MatchNum|AgencyName|AgencyGroup|OfficeName|TeamName|MatchType|MatchStatus|MatchName|MatchOpenDate|MatchCloseDate|SurveyType|YOSScheduledDate|YOSCompletionDate|YOSCompletionType|YOSStatus|Q1|Q2Neg|Q3Neg|Q4Neg|Q5|Q6|SocAccept|Q1b|Q2b|Q3b|Q4b|Q5b|Q6b|SocAcceptB|SocAcceptPrcnt|Q7Neg|Q8|Q9|Q10Neg|Q11Neg|Q12|SchComp|Q7b|Q8b|Q9b|Q10b|Q11b|Q12b|SchCompB|SchCompPrcnt|Q13|Q14|Q15|EdExpect|Q13b|Q14b|Q15b|EdExpectb|EdExpectPrcnt|Q16|Q17|Q18|Q19|Grades|Q16b|Q17b|Q18b|Q19b|Gradesb|GradesPrcnt|Q20Neg|Q21Neg|Q22Neg|Q23Neg|Q24Neg|Q25Neg|Q26Neg|RiskAtt|Q20b|Q21b|Q22b|Q23b|Q24b|Q25b|Q26b|RiskAttb|RiskAttPrcnt|Q27|Q28|Q29|PTrust|Q27b|Q28b|Q29b|PTrustb|PTrustPrcnt|Q30Neg|Q31Neg|Truancy|Q30b|Q31b|Truancyb|TruancyPrcnt|Q32|SpAdult|Q32b|SpAdultb|SpAdultPrcnt|Q33Neg|JJustice|Q33b|JJusticeB|JJusticePrcnt|MatchSupportLevel|MatchReportSources|MatchClosureReasons|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildGrade|ChildLivingSituation|ChildIncomeLevel|ChildFamilyAssistance|ChildFreeReducedLunch|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|ChildPartKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolPartKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|MatchKey|MatchTypeKey|SiteTypeKey|MatchActivityKey|SiteKey|StatusKey|MatchSupportLevelKey|MatchReportSourceKey|ChildReportSourceKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|YOSSurveyKey|PriorBaselineYOSSurveyKey|YOSStatusKey|YOSCompletionTypeKey|SurveyTypeKey|CustodialAdultEmployerHash
CM39|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM39|2015-04-14|2015-10-07|Baseline|2015-03-26|2015-04-14|Complete|Done|2|1|3|1|2|3|2|||||||||2|4|2|2|3|2|2.5|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Moved|5.8||1|2|1|1|F|Multi-race (Hispanic & White)||13|No|Mother|28205|7|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community||Pending Match|F|White||30|28205|Bachelors Degree|Separated|Business|28205|0|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504205508|504207619|35|0|2|504157187|1|0|2|500820606|2||-2||4|3|500014681||-2|500014681|-2|0|5|||17159|12|||1|863991|-1|4|3|44|610388910998118020
CM6|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM6|2015-04-30|2015-06-25|Baseline|2015-04-23|2015-04-30|Complete|Done|1|1|1|4|4|4|2.5|||||||||2|2|3|3|3|4|2.83|||||||||4|4|4|4||||||5|5|5|3|4.5|||||||4|4|4|4|4|4|4|4||||||||||1|4|1|2||||||4|1|2.5|||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|1.8||2|2|1|1|F|Black||11|No|Mother|28269|5|One Parent: Female|$50,000 to $59,999|Y|No||School|General Community||Match Support|F|White||27|28202|Some College|Single|Transport: Flight Attendant||2|1|Local TV|Media|Big|General Community||Enrollment|277|60|598|500000170|500017732|504243465|504245581|31|0|2|504173742|1|0|2|500824646|2||-2||4|1|||-2||-2|0|4|||7438|1|||1|873076|-1|4|3|44|2806833304218536184
CM78|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM78|2015-05-31|2016-03-14|Baseline|2015-05-14|2015-05-31|Complete|Done|4|2|4|1|3|4|3|||||||||2|4|4|3|1|4|3|||||||||3|2|4|3||||||2|3|1|5|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|PERL 2014-2016|Child/Family: Moved|9.5||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28134|4|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28273|Bachelors Degree|Single|Architect|28273|0|11|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|504202968|504205079|36|0|1|504285700|1|0|1|500827095|2||-2||4|2|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|881906|-1|4|3|44|7165641474360673060
CM87|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM87|2015-06-02|2016-04-27|Baseline|2015-05-05|2015-06-02|Complete|Done|3|2|4|1|4|4|3|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||3|4|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|10.8||1|1|1|1|M|Black||15|No|Mother|28273|8|One Parent: Female|$35,000 to $39,999||No|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||30|28208|Bachelors Degree|Single|Self-Employed, Entrepreneur|28078|2|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504159888|504161941|31|0|1|504240720|1|0|1|500825834|2||-2||4|3|500014681|500014681|-2|500014681|-2|34|2|||17159|12|||1|877407|-1|4|3|44|8491998754880714879
CM42|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM42|2015-06-18|2015-12-29|Baseline|2015-05-28|2015-06-18|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|4|3|2|4|3|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||4|3|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|6.4||1|1|1|1|M|Black||13|Yes|Mother|28214|5|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Asian|Indian|49|28203|Bachelors Degree|Married|Tech: Engineer|28204|10|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504217755|504219869|31|0|1|504131744|4|18|1|500828564|2||-2||4|1||500000294|-2||-2|34|2|||17159|12|||1|890821|-1|4|3|44|7000602719972091240
CM70|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM70|2015-06-23|2016-03-03|Baseline|2015-06-23|2015-06-23|Complete|Done|2|4|4|3|3|3|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016|Child/Family: Moved|8.3||1|1|1|1|F|Black||13|No|Mother|28134|6|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||30|28277|Bachelors Degree|Single|Business: Clerical|28277|1|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502205926|502206355|31|0|2|504225335|1|0|2|500831147|2||-2||4|1|500014681|500014681|-2||-2|0|5|||7464|9|||1|908891|-1|4|3|44|6178126991714892144
CM64|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM64|2015-06-28|2016-02-24|Baseline|2015-06-28|2015-06-28|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red|PERL 2014-2016|Child/Family: Time constraints|7.9||1|1|2|2|M|Black||11|No|Mother|28226|3|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|504198439|504200550|31|0|1|504230177|1|0|1|500831539|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||7462|13|||1|910542|-1|4|3|44|0
CM9|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM9|2015-06-29|2015-09-23|Baseline|2015-06-16|2015-06-29|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|3|1|2|4|3|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|2|3.71||||||||||3|4|4|3.67||||||3|1|2|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|2.8||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28031||Single|Service: Restaurant|28078|0|2|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504186384|1|0|1|500830331|2||-2||4|3|500014681|500014681|-2|500000294, 500014681|-2|0|4|||7464|9|||1|905704|-1|4|3|44|3402014428779854546
CM13|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM13|2015-08-11|2015-11-30|Baseline|2015-08-06|2015-08-11|Complete|Done|4|4|2|2|4|4|3.33|||||||||3|4|3|3|4|3|3.33|||||||||3|3|4|3.33||||||2|4|5|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Feels incompatible with child/family|3.6||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28212|6|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community|PERL 2014-2016|Enrollment|F|White||47|28270|Some College|Married|Homemaker|29020|18|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|504280484|504282684|36|0|2|504226821|1|0|2|500835375|2||-2||4|3|500014681|500014681|-2||-2|0|3|||7464|9|||1|924522|-1|4|3|44|4694273237201497095
CM10|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM10|2015-09-23|2015-12-29|Baseline|2015-09-11|2015-09-23|Complete|Done|4|2|4|2|4|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|Amachi|Child: Lost interest|3.2||1|1|1|1|F|Black||10|Yes|GrandMother|28217|4|Grandparents|Less than $10,000|Y|Yes||School|General Community|Amachi|Match Support|F|White||32|28277|Masters Degree|Divorced|Tech: Computer/Programmer|28277|0|3|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|504195472|504197572|31|0|2|504222207|1|0|2|500839514|2||-2||4|1|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|933343|-1|4|3|44|0
CM22|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM22|2015-10-21|2016-03-04|Baseline|2015-10-01|2015-10-21|Complete|Done|2|4|4|4|4|4|3.67|||||||||1|4|2|2|2|3|2.33|||||||||4|4|4|4||||||2|3|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||1|1||||4|4||||Green|PERL 2014-2016|Child/Family: Moved|4.4||1|1|2|2|M|Black||14|No|Mother|28212|5|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|Amachi, PERL 2014-2016|Enrollment|M|White||30|28209|Bachelors Degree|Married|Real Estate: Realtor|28217|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|503863366|503865360|31|0|1|504322037|1|0|1|500843765|2||-2||4|1|500014681|500000294, 500014681|-2||-2|0|5|||46|2|||1|939888|-1|4|3|44|0
CM34|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM34|2015-12-07|2016-05-24|Baseline|2015-11-06|2015-12-07|Complete|Done|3|4|2|2|3|4|3|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||2|3|4|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|5.6||1|1|1|1|M|Black||14|No|Mother|28027|7|One Parent: Female|$25,000 to $29,999||Yes||School|General Community||Match Support|M|White||24|28262||Single|Medical: Healthcare Worker|28025|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|502129820|502130249|31|0|1|504474407|1|0|1|500858150|2||-2||4|3|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|957862|-1|4|3|44|2881622112345502539
CM30|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM30|2015-12-14|2016-05-19|Baseline|2015-11-17|2015-12-14|Complete|Done|3|4|4|4|3|2|3.33|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|2|3|2.67||||||2|3|2.5||||||||||3|3||||Green|PERL 2014-2016|Volunteer: Moved|5.2||1|1|1|1|F|Black||16|No|Mother|28215|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||25|28205|Bachelors Degree|Single|Business|28031|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017777|503611723|503613600|31|0|2|504295160|1|0|2|500860670|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|10|||17159|12|||1|962728|-1|4|3|44|0
CM71|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM71|2015-12-17|2016-08-29|Baseline|2015-12-07|2015-12-17|Complete|Done|4|2|4|2|4|4|3.33|||||||||2|4|2|2|2|2|2.33|||||||||4|3|3|3.33||||||3|4|2|4|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment, PERL 2014-2016|Volunteer: Lost contact with child/agency|8.4||1|1|1|1|M|Black||14|No|Mother|28269|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||RTBM|M|Black||40|28269|Bachelors Degree|Married|Tech: Support, Writing|28269|4|0|Local Radio|Media|Big|General Community|Amachi, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|504245120|504247236|31|0|1|504396885|31|0|1|500865817|2||-2||4|1|500007920, 500011315, 500011316, 500014681||-2|500000294, 500007920, 500011315, 500011316, 500014681|-2|0|4|||7437|1|||1|970842|-1|4|3|44|1546374315672654438
CM2|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM2|2015-12-18|2016-01-08|Baseline|2015-12-08|2015-12-17|Complete|Done|3|3|3|3|4|4|3.33|||||||||2|4|3|3|4|4|3.33|||||||||4|4|4|4||||||2|4|3|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|0.7||1|1|1|1|F|Black||15|No|Mother|28269|8|One Parent: Female|$30,000 to $34,999||Yes||School|General Community|VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|F|White||26|28078|Masters Degree|Single|Business: Marketing|28269|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|277|60|598|500000170|500017777|504458036|504460294|31|0|2|504416792|1|0|2|500866388|2||-2||4|2||500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|971455|-1|4|3|44|3086452374500817499
CM56|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM56|2016-01-14|2016-08-29|Baseline|2015-11-09|2016-01-14|Complete|Done|3|3|3|1|2|3|2.5|||||||||2|3|3|4|3|4|3.17|||||||||4|4|4|4||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Lost contact with child/agency|7.5||1|1|1|1|F|Black||10|No|Mother|28056|4|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||RTBM|F|White||30|28209|Bachelors Degree|Single|Finance: Banking|28211|3|2|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|504407275|504409521|31|0|2|504393547|1|0|2|500857377|2||-2||4|1|500014681||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|958346|-1|4|3|44|0
CM51|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM51|2016-01-21|2016-08-29|Baseline|2016-01-11|2016-01-21|Complete|Done|3|4|4|1|4|4|3.33|||||||||2|2|3|2|1|2|2|||||||||4|3|3|3.33||||||2|5|3|4|3.5|||||||1|1|2|4|3|3|4|2.57||||||||||2|4|3|3||||||2|4|3|||||1|1||||3|3||||Green|PERL 2014-2016|Volunteer: Feels incompatible with child/family|7.3||1|1|1|1|M|Black||15|No|Mother|28269|7|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Multi-race (Black & White)||27|28115|Bachelors Degree|Single|Business|28115|4|4|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500017777|504268284|504270481|31|0|1|503172653|36|0|1|500871097|2||-2||4|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|981397|-1|4|3|44|2378213070582218846
CM14|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM14|2016-01-30|2016-05-20|Baseline|2016-01-14|2016-01-30|Complete|Done|4|2|4|4|4|4|3.67|||||||||2|3|3|3|1|3|2.5|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|Volunteer: Moved|3.6||2|2|1|1|F|Black||12|No|Mother|28214|5|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||32|28208|Bachelors Degree|Single|Journalist/Media||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503976557|503978568|31|0|2|504365048|1|0|2|500871811|2||-2||4|1|500007920, 500011315, 500011316||-2||-2|34|2|||7464|9|||1|982536|-1|4|3|44|3198188609986797983
CM74|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM74|2016-05-24|2017-02-23|Baseline|2016-05-10|2016-05-24|Complete|Done|2|1|1|2|1|1|1.33|||||||||3|2|3|3|3|2|2.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|2|1|2||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|9||1|1|1|1|M|Black||15|No|Mother|28208|9|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|PHD|Single|Self-Employed, Entrepreneur|30604|4|0|Local Print|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504347348|504349572|31|0|1|504566830|1|0|1|500892524|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|34|2|||7439|1|||1|1022954|-1|4|3|44|7044657180546140448
CM60|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM60|2016-05-27|2017-01-20|Baseline|2016-05-04|2016-05-27|Complete|Done|3|4|2|4|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|3|4|4|3.86||||||||||3|3|3|3||||||3|2|2.5|||||1|1||||4|4||||Red||Child: Severity of challenges|7.8||1|1|1|1|M|Black||14|No|Mother|28215|7|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|M|White||23|28205|Bachelors Degree|Single|Finance|28210|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500008321|504318423|504320644|31|0|1|504561410|1|0|1|500891770|2||-2||4|3|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1020756|-1|4|3|44|2141487034287122220
CM62|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM62|2016-05-31|2017-01-27|Baseline|2016-05-02|2016-05-31|Complete|Done|2|3|4|3|3|3|3|||||||||3|3|3|2|3|3|2.83|||||||||4|3|2|3||||||2|3|5|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|3|3|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|Volunteer: Lost contact with child/agency|7.9||1|1|2|2|M|White||14|No|Mother|28214|7|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community||Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|504231264|504233379|1|0|1|504230177|1|0|1|500891315|2||-2||4|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|0|3|||7462|13|||1|1019394|-1|4|3|44|0
CM25|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM25|2016-06-20|2016-11-03|Baseline|2016-05-11|2016-06-20|Complete|Done|2|2|3|2|3|2|2.33|||||||||3|3|3|2|3|4|3|||||||||4|4|4|4||||||5|3|1|3|3|||||||4|4|4|4|3|4|2|3.57||||||||||2|2|1|1.67||||||4|4|4|||||1|1||||3|3||||Green||Volunteer: Lost contact with child/agency|4.5||1|1|1|1|F|Black||14|No|GrandMother|28105|9|Grandparents|$45,000 to $49,999||Yes|BBBS National Site|Web Link|General Community||RTBM|F|Black||39|28105|Bachelors Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504631841|504634252|31|0|2|504167347|31|0|2|500892753|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|1023753|-1|4|3|44|5605796235524810842
CM8|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|CM8|2016-12-22|2017-02-28|Baseline|2016-12-01|2016-12-19|Complete|Done|4|1|4|4|4|4|3.5|||||||||4|4|4|1|4|1|3|||||||||4|4|4|4||||||1|1|5|5|3|||||||4|4|4|3|3|3|4|3.57||||||||||4|4|4|4||||||1|1|1|||||1|1||||4|4||||Red||Child/Family: Moved|2.2||1|1|1|1|M|Black||14|No|Mother|28215|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Black||32|28213|Masters Degree|Married|Finance: Auditor|28202|0|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500020753|504851045|504853547|31|0|1|504774982|31|0|1|500932246|2||-2||4|3||500014681|-2|500007920, 500011315, 500011316|-2|0|5|||46|2|||1|1112091|-1|4|3|44|2141487034287122220
