GroupB|ChildPartKey|VolPartKey
M2|501045214|500953330
M3|500261295|500188435
M4|500826592|501314246
M5|500186682|500887363
M6|500185601|501082220
M7|500546821|500790181
M8|500874765|502038804
M9|502142541|501905673
M10|500474486|500491064
M11|500186956|500189727
M12|500186106|500778380
M13|500186435|500189358
M14|502436202|502642999
M15|500395038|500392006
M16|501347056|501217000
M17|502045254|502171015
M18|502601023|502546883
M19|502824908|502891382
M20|500185907|500697782
M21|502893765|502874079
M22|502431164|502850528
M23|500408135|500189709
M24|500186260|500189139
M25|501516900|501438601
M26|502966254|502895517
M27|502714405|502764673
M28|501092911|501176101
M29|500799303|500798390
M30|500186905|500189677
M31|501300101|500346193
M32|500733695|500307108
M33|500185723|501310677
M34|501060196|501036081
M35|500968246|501179573
M36|500185571|500188438
M37|501641337|500835981
M38|501506214|501588885
M39|501645192|501519306
M40|502205848|502624702
M41|501868921|501382633
M42|502537477|500189507
M43|503236068|503976384
M44|501631547|502170945
M45|500871683|500933829
M46|501811385|502460013
M47|500186742|502397541
M48|501185594|501153366
M49|500186133|500188930
M50|501626226|502036832
M51|500997880|500990660
M52|502588461|502636478
M53|503469094|501717376
M54|501201377|501497622
M55|500185778|500188776
M56|502863781|503002010
M57|501402710|501728845
M58|503052841|503122069
M59|503268324|503253968
M60|502308593|502262702
M61|500185812|500188912
M62|500948129|501891556
M63|502185074|502490418
M64|503216769|503344849
M65|502570396|502545897
M66|502045258|502190790
M67|502510347|502677833
M68|500796255|501846438
M69|500252077|501365749
M70|502370669|503472866
M71|501237971|501598429
M72|503425736|503519747
M73|502421176|503497451
M74|500341548|504323327
M75|504043491|503984584
M76|501621811|501621016
M77|503026933|503758613
M78|500186645|500189545
M79|500887862|500923430
M80|502839827|503311280
M81|504031009|503971990
M82|501604443|501729878
M83|500826594|500920342
M84|501378357|501174997
M85|502578459|502869485
M86|502604900|502582742
M87|502974629|503188801
M88|501212047|501242250
M89|503110827|503278385
M90|502499851|502690262
M91|504447856|502087592
M92|504042248|502056302
M93|502982301|503442370
M94|502319972|502911091
M95|500814240|500981509
M96|500187081|500189197
M97|504070330|504032595
M98|501936316|501872326
M99|503026286|503259120
M100|504425940|502716664
M101|501000843|503106526
M102|502277840|503953636
M103|503671116|503672609
M104|503013779|501311929
M105|501919423|502034798
M106|504031043|503776239
M107|504031043|503956879
M108|500361200|500368628
M109|500378354|501181060
M110|501011735|502473442
M111|502725777|502710032
M112|502530688|502166996
M113|500931662|500894084
M114|503662199|503639494
M115|502255150|502392989
M116|501716763|502112513
M117|500186952|500189723
M118|502839019|502432390
M119|502702145|502204211
M120|503360420|503831013
M121|502570183|502570153
M122|500243491|502919490
M123|502172536|501279665
M124|502180719|502391505
M125|502551092|502366844
M126|502670076|501391123
M127|500938154|501446421
M128|504043289|502366876
M129|501300013|500346193
M130|500970495|500965698
M131|500970267|502084649
M132|502571727|502769619
M133|500958307|500876132
M134|503417576|503594017
M135|503255669|500188812
M136|502674024|502660051
M137|501157075|502978065
M138|503804225|503881040
M139|501309634|501046221
M140|503448711|503576769
M141|504493589|504314218
M142|502885468|502954219
M143|502371558|502528355
M144|502275241|502394690
M145|502129650|502598777
M146|501725162|501833178
M147|503124706|503609606
M148|502526965|502881104
M149|502431187|503015009
M150|503546374|503890372
M151|500271303|501291358
M152|504447951|504272897
M153|500724632|500803551
M154|502124485|501905673
M155|504042320|502779828
M156|502589869|502701252
M157|502912141|502932948
M158|502197477|502422929
M159|502206673|502668179
M160|504043455|503972115
M161|504454538|504311707
M162|504513842|504431507
M163|501361902|501307192
M164|503476243|503334174
M165|502700505|503029324
M166|500545328|501033808
M167|500545326|500697845
M168|502083429|502653045
M169|501726201|501734664
M170|503833956|503635291
M171|501786018|503914867
M172|501376745|500725077
M173|504043477|501245666
M174|503533026|502485670
M175|502067798|502062408
M176|501529921|502554719
M177|502702827|503969458
M178|504495905|504366540
M179|501083790|503984623
M180|501428903|501441245
M181|504445088|504368282
M182|502133283|504277979
M183|503014417|503518076
M184|504447755|504434419
M185|502307585|501519450
M186|504043271|503974114
M187|502920861|503097126
M188|502570188|502366830
M189|504447916|504130536
M190|503635703|503979778
M191|501340097|501934966
M192|502710796|502926804
M193|504426368|500863980
M194|500764138|503707921
M195|504043114|502261758
M196|504447778|504350981
M197|502097843|502643791
M198|504043467|503971844
M199|500340183|503868914
M200|503443162|500234684
M201|502828131|502881454
M202|500829028|501978180
M203|502868969|503574667
M204|502469903|502868874
M205|504043252|503974167
M206|504059403|503658554
M207|503813942|503873603
M208|504043100|503962672
M209|504043445|503922166
M210|502602958|502578040
M211|504169896|503987952
M212|501195410|501277677
M213|503873575|504004351
M214|503923102|503996589
M215|504426028|504357594
M216|503796616|503828896
M217|502761850|503632186
M218|503216855|503969586
M219|503587930|500942257
M220|501735420|500956022
M221|500713817|501834795
M222|501234606|501233675
M223|502221847|502654877
M224|502551045|503859553
M225|504454510|504357339
M226|502763473|502828246
M227|504050643|503969686
M228|504426151|504431643
M229|504043352|503969666
M230|501833031|502427342
M231|502580335|502677590
M232|503524036|503913408
M233|504454500|503529603
M234|503767186|503788125
M235|504085882|503977000
M236|503236129|503682677
M237|503236129|504434419
M238|503236165|503163281
M239|501096791|503803014
M240|504043184|504024311
M241|504043120|503974816
M242|502555551|503207140
M243|503578835|503605630
M244|500824037|500789337
M245|504842862|504300098
M246|504043105|503969642
M247|504180420|504001561
M248|502581328|503144090
M249|502063945|502295138
M250|502338225|502312449
M251|500186245|502989318
M252|501227649|503316978
M253|504050627|503976447
M254|504445059|501631588
M255|500783100|500777047
M256|503296945|503381327
M257|502760967|502666332
M258|500905037|501564519
M259|504050561|503971898
M260|501631140|501628976
M261|503149009|503199095
M262|500740296|502893901
M263|502234504|502129464
M264|504043501|504001561
M265|504454641|500800975
M266|504425996|504272278
M267|504494261|504423999
M268|503602174|503615576
M269|502171910|502141964
M270|502866475|502961396
M271|504447927|503868542
M272|504447891|503984584
M273|504447891|504739188
M274|503983132|503995895
M275|504440300|504313945
M276|503597088|503642924
M277|502478428|502555822
M278|503496889|503490051
M279|501597228|501397328
M280|502319984|502290677
M281|504426057|504363902
M282|502537469|502056302
M283|502537469|503323641
M284|504419900|504351222
M285|501143674|502958999
M286|500826100|503877762
M287|500910037|500856100
M288|500843863|501078655
M289|504445029|504272155
M290|501288021|501249338
M291|500936718|501027885
M292|504043155|503985283
M293|504099617|503984599
M294|501825910|501196986
M295|504447802|504350780
M296|502610186|502913393
M297|504426106|504355965
M298|503187841|503789478
M299|501604887|503999324
M300|500465506|500496966
M301|504104035|504214658
M302|501353940|502710990
M303|504043305|503776239
M304|501376223|503976447
M305|501376223|503969375
M306|502064627|500773055
M307|502482642|503118336
M308|502264006|502274748
M309|502766037|503605985
M310|501525308|501536144
M311|504063426|504152304
M312|501074345|501158523
M313|502753870|503869569
M314|502531929|504397371
M315|502549829|502594393
M316|500934908|502107314
M317|502552947|503881539
M318|502393980|502928199
M319|504043202|503971855
M320|503712470|503952262
M321|504050578|503969533
M322|504043211|503969563
M323|500395499|501027885
M324|500280148|502118494
M325|504089115|504081485
M326|504090244|504121323
M327|503611723|504295160
M328|504449675|504461244
M329|504426315|503796728
M330|502593613|502601730
M331|503225805|503317460
M332|504454746|504339857
M333|503212298|500189616
M334|502304267|503343217
M335|504269922|504285435
M336|500727291|500857838
M337|502179379|502161458
M338|504034181|504053608
M339|504454486|504300098
M340|503624220|503605851
M341|503379566|503407492
M342|504495937|504355841
M343|500382177|500188566
M344|503472839|503503841
M345|503395663|503735537
M346|502589865|502625828
M347|503681619|503680923
M348|504419831|503985283
M349|504426322|503972115
M350|504425700|504445539
M351|503955527|504285092
M352|504426175|504445758
M353|503934189|503918487
M354|503678291|503680714
M355|503556065|501284751
M356|503441463|504122275
M357|504460043|504314082
M358|504831646|503605851
M359|502193174|503100143
M360|502876870|503104166
M361|503690133|503605679
M362|503484186|503355490
M363|501434147|501926474
M364|501721760|501755476
M365|502591898|503002003
M366|502787401|503122442
M367|503326540|503852999
M368|504419824|504455318
M369|504425599|504349061
M370|504004117|503929259
M371|503681650|503661517
M372|502980965|503091130
M373|502980958|503008664
M374|504456568|504380428
M375|500847570|502542379
M376|504426348|504363925
M377|501842678|502335257
M378|502979759|503234517
M379|500826603|502672644
M380|503681628|504024551
M381|504888350|503599329
M382|504454736|503605671
M383|504451240|504432323
M384|502552438|502549491
M385|504447817|504422986
M386|504416080|504349689
M387|503746685|503961087
M388|500765381|501579025
M389|504129007|504137446
M390|502828137|502446364
M391|502402515|502537081
M392|502244776|502143351
M393|504440280|503028265
M394|504831472|504339626
M395|503606415|503665457
M396|504447831|504349089
M397|503635439|503605799
M398|503503500|503390470
M399|504445105|504447607
M400|504454672|503885836
M401|501725168|503828482
M402|504235352|504200139
M403|504449679|504447687
M404|503318447|503537303
M405|504425892|504352616
M406|504451307|504356262
M407|504393421|504395484
M408|504154291|503862054
M409|504031334|503882331
M410|503216820|504024735
M411|504419837|504368264
M412|503602228|503605726
M413|501833026|502451325
M414|504444913|504272227
M415|504447870|504320091
M416|500796261|503790153
M417|504440272|503281135
M418|501194563|503477116
M419|504444978|504357304
M420|503005868|502935610
M421|500496598|501383928
M422|504023342|504173078
M423|504207073|504201268
M424|504440264|504267500
M425|504454695|503605851
M426|504159888|504240720
M427|503821678|504468148
M428|504883840|504742660
M429|504287270|504024992
M430|503805173|503799347
M431|504425766|504287751
M432|504445152|504355816
M433|503532788|503939365
M434|504426069|504350928
M435|502990571|503400909
M436|504444999|504448559
M437|504445133|503969458
M438|504425789|504287751
M439|504425789|504353872
M440|504148143|504559007
M441|502317500|502658498
M442|501224282|503347558
M443|504089161|504078362
M444|504089161|504393611
M445|500545470|500815012
M446|503834613|503790527
M447|504081466|504098772
M448|501076082|502687269
M449|503533022|503534544
M450|504075196|504108003
M451|504428620|504035546
M452|502859187|503090888
M453|502030263|501923553
M454|503634083|503605644
M455|501247269|501914025
M456|504444952|504284272
M457|502809446|502909383
M458|500570756|502889143
M459|504440287|504382284
M460|504397554|504206321
M461|504454712|504214615
M462|502501997|504227306
M463|504440292|504364944
M464|502247579|502681447
M465|501401583|504338671
M466|502051702|503378835
M467|504425918|504383897
M468|504174131|503997551
M469|504416061|504465459
M470|501253195|500395148
M471|504289347|504428167
M472|504416147|504212639
M473|503569117|503583743
M474|504454572|504359810
M475|502549826|501223094
M476|502549826|503431300
M477|502549826|504037091
M478|503831166|503861120
M479|504220177|504309758
M480|502699353|503945609
M481|501989028|503039778
M482|504425672|504448500
M483|503023832|503139766
M484|503831971|504011759
M485|502255225|502312682
M486|504440275|504342087
M487|501904523|503979230
M488|502845758|502944923
M489|504454594|504249944
M490|501811395|500876892
M491|504440268|504315884
M492|504831598|504431507
M493|501332658|501814288
M494|502495501|502508181
M495|503803718|503930530
M496|502983808|503140432
M497|504416042|504072039
M498|504416042|504557665
M499|503041998|503110820
M500|502146600|503483337
M501|501604446|502664359
M502|504451288|503976447
M503|503635399|503605621
M504|501068963|503906067
M505|502612404|504226710
M506|502612404|503790988
M507|502663937|503296990
M508|504454656|504387544
M509|504347348|504566830
M510|504454566|504448602
M511|501641325|501715652
M512|501627668|503921388
M513|502270499|502510107
M514|501010684|503491643
M515|501123191|502153920
M516|504831621|504357339
M517|503611732|504421910
M518|503681630|503162750
M519|504831552|504359810
M520|502180724|502391505
M521|500784687|503531111
M522|502287066|504056150
M523|504976123|504685043
M524|500917189|504538036
M525|504473782|504550297
M526|504834787|504808345
M527|504662357|504791469
M528|503230648|503169561
M529|501611456|501876475
M530|503974135|503860995
M531|503974135|504341793
M532|504842890|504780315
M533|503246887|503253208
M534|504454583|504274695
M535|504842854|500953330
M536|504089143|504072039
M537|501372080|502500246
M538|504089098|504037139
M539|501809541|501620528
M540|504076406|503831499
M541|504416180|503630789
M542|504416180|504399592
M543|504834756|504767391
M544|502252828|502602451
M545|504423117|504359583
M546|501716720|501878786
M547|503728057|503788318
M548|504831502|504775164
M549|503899239|503871007
M550|503722616|503707316
M551|503722616|504343006
M552|503623969|503976684
M553|503635425|503606058
M554|504039275|504461897
M555|504526221|504349689
M556|504526221|504396970
M557|503633871|503855574
M558|504183446|503979203
M559|504183446|504267362
M560|501247286|501247141
M561|504312104|503754104
M562|504312104|504766848
M563|504471621|504580592
M564|503782093|504545677
M565|501390344|501380163
M566|501390345|502966998
M567|502979699|504127445
M568|503413167|504190868
M569|503044619|503021454
M570|502821865|504267500
M571|503678239|500189616
M572|503678239|503689039
M573|501831581|500715453
M574|503071479|503051382
M575|504410184|503979778
M576|501529924|502199360
M577|504458036|504416792
M578|502569117|502538689
M579|504859855|504784459
M580|504416166|503799347
M581|501536733|501418563
M582|504698283|504765309
M583|501185592|501255830
M584|501771263|501622704
M585|504831667|504780301
M586|504089123|504383897
M587|504089123|503680769
M588|503624276|504786758
M589|503770826|503820142
M590|503328958|503574852
M591|501253965|502985911
M592|503944459|504260502
M593|504089059|504024774
M594|504416202|504394234
M595|504268284|503172653
M596|504207081|504060437
M597|500961274|500403000
M598|503770380|503833456
M599|503758675|503792275
M600|504428649|504396801
M601|503704573|503883049
M602|502183217|501733851
M603|503707241|503767700
M604|503863366|504322037
M605|502896719|502959645
M606|503224764|504130394
M607|504831713|504380428
M608|503318449|503775488
M609|501599416|500188567
M610|502183053|503073638
M611|504631841|504167347
M612|504160892|504171934
M613|502566369|503065299
M614|504870363|504719047
M615|504506841|504024774
M616|503219503|503589945
M617|503816186|504090792
M618|502920377|502942994
M619|503566749|503605700
M620|503063769|504299841
M621|503511553|503504991
M622|500868942|500947018
M623|503110829|503130981
M624|503917561|504206321
M625|502229042|503849760
M626|504526211|504528256
M627|503634718|503595858
M628|503961917|504052039
M629|504831449|504719321
M630|504910946|504687842
M631|501938282|502356100
M632|501152789|503604690
M633|502245129|502670839
M634|504298668|504372921
M635|504831525|504765443
M636|503492214|504272278
M637|503021417|503115600
M638|501662021|503759352
M639|501091420|503946168
M640|504081573|503880925
M641|504081573|504317495
M642|502000252|502127058
M643|502902247|502801082
M644|503515724|503689721
M645|502008563|503400112
M646|504416129|504399706
M647|501147999|503112265
M648|504888396|504767070
M649|502700503|502931327
M650|504231264|504230177
M651|503813952|503829786
M652|504416115|504397175
M653|504842873|503969533
M654|501273088|503079327
M655|503952645|503942996
M656|503923436|501306527
M657|504333795|504348509
M658|503535105|504127300
M659|504859921|504353872
M660|504416012|504397015
M661|503838769|503948333
M662|504861242|504786813
M663|501069450|500887364
M664|504416100|504455617
M665|503874068|504196201
M666|503361148|502459922
M667|504045474|504228594
M668|504087114|503605618
M669|502863776|503029273
M670|501014187|501404007
M671|502303088|502445797
M672|502335675|502305990
M673|503849038|503930671
M674|502858216|503376842
M675|504831574|504756883
M676|504831771|504784525
M677|504245120|504396885
M678|501213488|501225276
M679|503587461|503541106
M680|502254067|503590595
M681|501092822|503854063
M682|501092822|503854063
M683|503441472|503551607
M684|504855873|504783357
M685|502178448|504024654
M686|504851045|504774982
M687|502619926|504288677
M688|502619926|502642260
M689|502273093|502252422
M690|504842845|504794021
M691|503711736|501121735
M692|504831791|503529603
M693|502183420|502264770
M694|503937201|503582646
M695|503913977|503898216
M696|503913977|503898216
M697|504867822|504743932
M698|504880135|504738710
M699|502829894|503443998
M700|504574961|504676344
M701|502549830|504035546
M702|502549830|502462453
M703|502107146|504090344
M704|504221476|504231286
M705|504831698|504751575
M706|503690173|503604304
M707|504318423|504561410
M708|502359051|502242295
M709|501788776|501698382
M710|502825916|502367677
M711|504154297|504201847
M712|503999208|503973970
M713|502753873|503146044
M714|502186245|504248899
M715|503016111|503135600
M716|502436198|503255826
M717|503643026|503377601
M718|503643026|504315865
M719|503791020|503783913
M720|501143676|503315012
M721|503803127|503866013
M722|504129013|504577506
M723|504150667|503845717
M724|504150667|504242094
M725|503217134|503605778
M726|503633782|502441938
M727|504089044|503255983
M728|503524258|500497043
M729|504333730|504349844
M730|503602213|503606038
M731|503544893|503844843
M732|504054633|504068503
M733|502776307|502483716
M734|502255156|502946412
M735|502529397|500188946
M736|503999199|503973076
M737|504348416|504242094
M738|503479095|503915425
M739|501863951|501601161
M740|504013295|504146637
M741|504545166|503788318
M742|503021552|502951522
M743|504396237|503604304
M744|503497835|503507978
M745|504855816|504839044
M746|504410234|504368847
M747|503429736|503850437
M748|502943644|503671882
M749|502943644|503899413
M750|503166335|503729353
M751|502875279|504151222
M752|503999194|503611445
M753|503017622|503095382
M754|504172774|504040677
M755|502945480|502919780
M756|501142903|501236825
M757|501721579|501687513
M758|503381531|500540549
M759|503690154|502542324
M760|504396225|503605618
M761|504410165|504445343
M762|504410165|504403681
M763|504416580|504504983
M764|501721762|503471102
M765|501721761|503023854
M766|502236953|502232559
M767|504013291|503979108
M768|503941174|503207130
M769|502308197|502325667
M770|502506397|503039829
M771|504057301|503796968
M772|504057301|503796968
M773|502821218|504244628
M774|501843066|504152982
M775|504076403|504415946
M776|502507408|502673562
M777|504170222|503853917
M778|501295538|502897530
M779|503756716|503596238
M780|504038196|504062905
M781|504235369|503937954
M782|502225378|502245842
M783|502129820|504474407
M784|503452963|503489818
M785|503717073|503853194
M786|503652810|500189256
M787|502336272|503743688
M788|501222138|500189173
M789|503972507|500189600
M790|502222545|502196116
M791|502255210|502255794
M792|501254255|501356688
M793|504007361|503605824
M794|504507791|504650231
M795|504655474|503853917
M796|502197486|502870668
M797|503953654|503976139
M798|502255223|501823103
M799|503217214|504373953
M800|503217214|503350133
M801|502583662|503943422
M802|502583662|504286292
M803|502583660|503944507
M804|503679979|504191848
M805|504410212|503973076
M806|504691840|504535890
M807|502278985|500220237
M808|503552606|501052547
M809|504732530|504893030
M810|503755565|503814505
M811|504013056|503976618
M812|504013056|504219921
M813|503632799|503567146
M814|501332660|503579743
M815|501332660|504556335
M816|502605331|503090281
M817|504348425|503911472
M818|501252806|501320197
M819|504416818|503988229
M820|503617980|503573243
M821|503421607|503520561
M822|504284556|504260574
M823|503654364|504076011
M824|501314104|501170940
M825|503917550|504577899
M826|504013304|503910182
M827|504564027|504766711
M828|501662033|503655814
M829|503977573|501601161
M830|503977573|504047655
M831|503662377|503573326
M832|504410257|503979108
M833|504401898|504875613
M834|503052850|503028888
M835|504331538|503843020
M836|504439764|504392917
M837|503959684|503985328
M838|503535102|503882165
M839|503989203|504066226
M840|503268271|502993922
M841|502868923|502832013
M842|504999127|504999362
M843|504230613|503995309
M844|504333777|504355120
M845|501837686|503754104
M846|504425160|504509415
M847|501755470|502038804
M848|503328946|503371779
M849|501319029|504558901
M850|501319029|503078205
M851|503452335|503845505
M852|504068125|504241807
M853|504152757|503979778
M854|502866083|503378884
M855|502866079|503378886
M856|504507408|504651211
M857|504401907|504355133
M858|501722052|502030533
M859|501597169|501563612
M860|504333786|504359851
M861|502763524|503839682
M862|502763524|504370632
M863|502763524|504370632
M864|503413169|504092153
M865|503292843|503233785
M866|504893713|504783221
M867|503628199|503966130
M868|504328960|504215323
M869|504855805|503605799
M870|504401919|504396776
M871|504416613|504368299
M872|504416613|504776839
M873|503462811|503365326
M874|504672339|504870474
M875|502728289|502339145
M876|502721278|502701096
M877|502700500|502824634
M878|502763379|503613615
M879|504410201|503605799
M880|502551048|501472128
M881|502912138|503857059
M882|502763968|502939016
M883|504205508|504157187
M884|503870487|503813685
M885|503915384|503995835
M886|504517520|501284751
M887|504517520|504355611
M888|503610365|503615532
M889|503879123|503889097
M890|503688885|503606993
M891|504396338|504353900
M892|503898651|503494199
M893|501712048|502405439
M894|502353937|501672025
M895|503723868|503940354
M896|504100809|503979771
M897|502249189|502485458
M898|503405468|502944301
M899|503405468|504322859
M900|504401940|504368976
M901|503743876|503908096
M902|504602680|504579649
M903|504868978|504855899
M904|504423105|503911379
M905|503851354|503962684
M906|504202968|504285700
M907|504748250|504885284
M908|503506115|503552068
M909|502987717|503559146
M910|504348606|504368342
M911|504038302|504099787
M912|504030009|503910147
M913|502939347|503598887
M914|504410173|504350008
M915|502997224|502939526
M916|502576641|502537061
M917|502471024|502685747
M918|502073665|503245956
M919|503924157|504277947
M920|504808434|504557160
M921|502205926|504225335
M922|504875016|503908898
M923|504250982|504349938
M924|504416684|504338378
M925|504237243|504456306
M926|503833936|502489398
M927|504139056|503991266
M928|503063881|503125383
M929|504247189|504228103
M930|503671715|503576626
M931|503671715|504324165
M932|504423077|504359606
M933|503594290|503508074
M934|502930499|502564910
M935|503770823|503850589
M936|503689574|503577882
M937|504165911|504030347
M938|504626085|504396349
M939|504333815|504348456
M940|504431587|504475369
M941|501859854|502044100
M942|503893808|504546078
M943|503893808|503976460
M944|503163476|503119713
M945|502335365|503603503
M946|504633835|504775410
M947|504161470|504396335
M948|503718061|503472779
M949|502375449|503493703
M950|502969236|503567563
M951|504242976|504198992
M952|502728419|504011804
M953|504007349|503981896
M954|503629812|503497377
M955|504450770|504359867
M956|504218954|504099424
M957|504217755|504131744
M958|502097794|502425119
M959|502184849|503145815
M960|503071350|503421602
M961|503071350|500831828
M962|503281941|503907559
M963|504517593|504526149
M964|503996783|503911472
M965|504554067|503373934
M966|504333747|504359691
M967|501951335|504368723
M968|502261100|502284382
M969|504416740|503355514
M970|502252822|504229640
M971|503692165|503216970
M972|502083438|502657267
M973|501853851|502922901
M974|503012569|502949193
M975|503756602|503825615
M976|504075185|504169746
M977|502335325|503500437
M978|504416703|504401855
M979|502392338|504744814
M980|504410188|504335835
M981|502385620|503633995
M982|502335383|503493859
M983|502262109|503605726
M984|504348774|503911351
M985|502882034|502983700
M986|503584428|503839843
M987|502786012|503553020
M988|502813481|503009633
M989|504025425|503948833
M990|502722096|504213418
M991|503575828|504188100
M992|503575828|504686759
M993|503241922|503507368
M994|504416720|504438102
M995|504030013|503910089
M996|502416642|503500482
M997|503663975|503854225
M998|503663975|504468271
M999|502634923|501197016
M1000|504280484|504226821
M1001|504910266|504829494
M1002|503666549|504106972
M1003|503666553|500991324
M1004|504869056|504788305
M1005|503034769|503650997
M1006|504100841|503964951
M1007|504016980|503931457
M1008|503469072|503478672
M1009|503469072|504202910
M1010|504155180|502462446
M1011|504431606|504355024
M1012|502637766|503016558
M1013|502375441|503507295
M1014|502582366|503858870
M1015|503710095|503872736
M1016|503496815|503673962
M1017|503250358|504861106
M1018|504338170|504465810
M1019|502747706|502618438
M1020|504399552|504544485
M1021|504853140|503605824
M1022|503610226|503935226
M1023|504013021|503910269
M1024|504792692|504760167
M1025|504416788|504353866
M1026|502873189|502882530
M1027|503720575|503714604
M1028|504976117|503605644
M1029|502207223|503251424
M1030|502355228|503507223
M1031|503869451|504135282
M1032|503552498|503538554
M1033|504855744|504783146
M1034|503774057|503665969
M1035|503532014|503694720
M1036|503532014|504408440
M1037|504626128|504632567
M1038|503207102|503688236
M1039|504417121|504579745
M1040|504143296|503540922
M1041|504358312|504048355
M1042|504937152|504797758
M1043|504474573|504349165
M1044|504474573|504685043
M1045|501806165|501706064
M1046|504416598|502432606
M1047|502183411|500189229
M1048|502787404|503485414
M1049|504416752|504396349
M1050|504025428|503911351
M1051|504333764|503908898
M1052|504517710|504475369
M1053|504626092|504349844
M1054|504410223|504445343
M1055|503637786|503577771
M1056|504054004|504265163
M1057|502097375|503901690
M1058|504410217|504359867
M1059|504592666|504625671
M1060|504176462|504109704
M1061|503418316|503493771
M1062|504736266|504634630
M1063|503704203|503493888
M1064|503704203|504297059
M1065|503995803|503963125
M1066|504013115|503675532
M1067|503547661|503731665
M1068|503884921|504160910
M1069|503952082|504546069
M1070|503629807|503603514
M1071|503533041|504183712
M1072|502552445|502545537
M1073|502395420|503497477
M1074|503946469|504188283
M1075|504410249|504369534
M1076|504869115|504349938
M1077|504436181|504741299
M1078|503821686|504460050
M1079|503229410|503493684
M1080|504396333|502542324
M1081|502278991|502263116
M1082|502335396|503507119
M1083|503704276|503507098
M1084|503704276|504306171
M1085|504628514|504599441
M1086|504333802|504354941
M1087|504463138|504819424
M1088|504176233|503500482
M1089|504471617|504458762
M1090|502458458|504387453
M1091|502979757|503161988
M1092|502234905|504334608
M1093|502234905|502799047
M1094|504227502|504460839
M1095|503270485|504039802
M1096|503270485|504574450
M1097|504231267|504379684
M1098|503978153|504039547
M1099|504489376|504604779
M1100|502933371|503080292
M1101|502933371|503911379
M1102|504886657|504807149
M1103|504200641|504222624
M1104|502173768|503831898
M1105|503807556|502105224
M1106|503636487|503899296
M1107|503590328|503874645
M1108|502223076|502694717
M1109|503895740|503765053
M1110|503895740|504364485
M1111|504171035|504150234
M1112|502761742|503041890
M1113|504013104|503933411
M1114|504333758|504484385
M1115|504437000|503979153
M1116|504427276|504354996
M1117|503512877|503893014
M1118|504039826|503980178
M1119|504275306|504359606
M1120|504038458|503971368
M1121|504200631|503404737
M1122|504416771|504349862
M1123|501314348|502205797
M1124|504396318|503605621
M1125|503976557|504365048
M1126|503976557|504538747
M1127|504038255|504034443
M1128|503254146|503509874
M1129|504049432|503908413
M1130|504410241|503605964
M1131|503701025|503576358
M1132|504040012|503935151
M1133|502789637|504034331
M1134|502789637|503542037
M1135|502789637|504703410
M1136|503355095|503373533
M1137|503401214|503758808
M1138|504133883|503868128
M1139|503756537|503403281
M1140|503281891|503507494
M1141|502234486|504359670
M1142|502813499|503633204
M1143|504133877|503908101
M1144|504310625|503442370
M1145|504439749|503605644
M1146|504886640|503754104
M1147|504205445|503796968
M1148|504030001|503935202
M1149|502245343|502526001
M1150|504133872|504225360
M1151|504041825|503907538
M1152|504041825|504303741
M1153|504416044|504623074
M1154|503472232|503444888
M1155|504861201|504804012
M1156|504051660|504277513
M1157|504049365|503908435
M1158|503629858|503507250
M1159|503629858|504303791
M1160|502347820|502419409
M1161|502347820|504547241
M1162|503689205|503689218
M1163|504530586|503694720
M1164|504861229|504798600
M1165|503770372|503594093
M1166|504675071|500353496
M1167|502391396|503228398
M1168|504065282|504168627
M1169|504886567|504799615
M1170|504861191|504783413
M1171|504103367|503907299
M1172|504908795|504024654
M1173|504890014|504807342
M1174|504016998|503931397
M1175|503718040|503449923
M1176|503492220|503521240
M1177|504260159|504639152
M1178|503530345|502460114
M1179|503312337|504201470
M1180|504112178|503916397
M1181|504085860|503605925
M1182|504870329|504814162
M1183|503703048|503354824
M1184|504150685|504378557
M1185|504150685|504186384
M1186|502875668|503114677
M1187|504268884|504240747
M1188|504565095|504860995
M1189|504878306|504775341
M1190|503777913|503572872
M1191|503777913|503907463
M1192|504290756|504315689
M1193|502559020|503590913
M1194|503602276|503381037
M1195|504899975|504359583
M1196|504861210|504890087
M1197|504998006|504303308
M1198|503885975|504620475
M1199|503885975|503885544
M1200|504019066|503931438
M1201|504152161|504180963
M1202|504886516|503255983
M1203|502969243|503837125
M1204|503739899|503802084
M1205|503652763|503985312
M1206|504280334|504556921
M1207|503637810|503603518
M1208|503637810|503901690
M1209|503565188|503814392
M1210|503565188|504265907
M1211|504861159|504801626
M1212|502629201|502893231
M1213|504870336|504348456
M1214|503424337|503446943
M1215|503195998|503507195
M1216|503195998|503905482
M1217|504869078|504359691
M1218|502290468|502873884
M1219|502383218|504867282
M1220|503629852|503613527
M1221|503629852|503907559
M1222|504861120|504242094
M1223|502222548|502214317
M1224|502367953|502658210
M1225|504932757|504311367
M1226|504908812|504024992
M1227|504536121|504562411
M1228|504539986|504793129
M1229|504908748|504821304
M1230|504103364|503907420
M1231|502776261|503995722
M1232|502776261|503540978
M1233|502068488|503953186
M1234|503486227|503555261
M1235|503810996|503799211
M1236|504861100|504798309
M1237|504166613|503823941
M1238|504106278|504043172
M1239|504890029|504060437
M1240|502763403|503603510
M1241|502763403|503905493
M1242|503866348|503862591
M1243|502162237|503151333
M1244|503707963|503507325
M1245|503707963|504302535
M1246|503770356|503479599
M1247|504070362|503507276
M1248|504234460|503812408
M1249|504875023|504475369
M1250|504540553|503680923
M1251|503670769|503493268
M1252|503670769|503905510
M1253|504312629|504262612
M1254|504312569|504208036
M1255|503941222|503889588
M1256|503929747|503910740
M1257|503644180|503493918
M1258|503644180|504327166
M1259|503638969|503503174
M1260|503391535|503497423
M1261|503391535|504306107
M1262|502431040|502609637
M1263|502766031|501946079
M1264|504343306|504109000
M1265|503565637|503604089
M1266|504049262|503907248
M1267|504890059|504394474
M1268|504878293|504632567
M1269|503196044|503509836
M1270|503196044|504324154
M1271|502746641|503540909
M1272|502746641|503907262
M1273|504671571|504308223
M1274|504890041|504817368
M1275|504861049|504354941
M1276|502527969|503169378
M1277|503996753|503911411
M1278|504049370|503517772
M1279|504049370|504301152
M1280|503259350|503370160
M1281|504908826|504829966
M1282|504240231|504523981
M1283|503204695|503506209
M1284|503204695|504301092
M1285|503779546|504625641
M1286|503669127|504220439
M1287|504870344|503911379
M1288|504870349|504359606
M1289|504870355|504798428
M1290|503779482|504510616
M1291|503779482|503108667
M1292|502763413|503577783
M1293|502763413|503907351
M1294|504960112|504789046
M1295|504013280|503908838
M1296|504629037|504619538
M1297|503686272|503817633
M1298|503691322|503763297
M1299|504184668|503338695
M1300|503143377|503109316
M1301|503196065|503497346
M1302|503196065|504308470
M1303|503745285|503655183
M1304|502934728|503516330
M1305|504886538|504829898
M1306|503609425|503837417
M1307|504230975|504284612
M1308|503723888|503858682
M1309|502602926|503808719
M1310|504861132|504771994
M1311|503217239|503666439
M1312|502299232|503510609
M1313|502653228|502192090
M1314|504861085|504391145
M1315|504870325|504349862
M1316|504041972|503897715
M1317|502324604|502657850
M1318|502211032|502276859
M1319|503492511|503852376
M1320|504635786|504662207
M1321|504026659|504744796
M1322|502274606|502441954
M1323|504100771|504000676
M1324|503650948|504063702
M1325|504357732|504576046
M1326|503644199|503540939
M1327|503644199|504296433
M1328|504153965|504372591
M1329|503470937|500188541
M1330|504886558|504822645
M1331|504944637|504324154
M1332|504908775|504806684
M1333|504041849|503995703
M1334|504110036|504043678
M1335|503629844|503608281
M1336|503629844|504307866
M1337|504030027|503908898
M1338|503408595|503490264
M1339|504870394|504557665
M1340|503996736|503880784
M1341|504083467|504003996
M1342|504861175|504952358
M1343|504861175|504349844
M1344|503503497|503775803
M1345|503637763|503507441
M1346|503637763|504307795
M1347|504878263|504797062
M1348|502749239|503507342
M1349|502749239|503905466
M1350|504526251|504475303
M1351|504134537|503852298
M1352|504005669|503908386
M1353|504942804|504807056
M1354|502464508|502901720
M1355|504628103|504469742
M1356|502426625|504274174
M1357|503569115|503619714
M1358|503623886|504803107
M1359|503745242|503480703
M1360|502859181|502638002
M1361|503795417|503762193
M1362|503741920|503696505
M1363|503741920|504976126
M1364|504870414|504787136
M1365|504662612|504595097
M1366|503718051|503489016
M1367|502298007|501202092
M1368|504059510|504000163
M1369|504059510|504359587
M1370|504221885|504188499
M1371|502842247|503305101
M1372|504049252|503901627
M1373|504049252|504297141
M1374|503198334|503907463
M1375|503904008|503820652
M1376|504714089|504679648
M1377|504388136|504360253
M1378|504388136|503869569
M1379|504526331|500994796
M1380|502619308|503710698
M1381|503545940|503804018
M1382|504577421|504771021
M1383|504049238|503907477
M1384|504049238|504297082
M1385|504198439|504230177
M1386|503704249|503497234
M1387|503704249|504303308
M1388|504619450|504619589
M1389|504619450|504884038
M1390|503794892|504175530
M1391|504041768|503907444
M1392|504041768|504296433
M1393|504937026|504303240
M1394|504468539|504306056
M1395|504526307|504441484
M1396|503418236|503671882
M1397|504531588|504127246
M1398|504093590|503907351
M1399|504042013|503999137
M1400|504970052|504743981
M1401|504952387|504306107
M1402|503214533|503540968
M1403|503214533|504307950
M1404|502982459|503565143
M1405|502982459|504669593
M1406|504184746|504183176
M1407|504059549|504109643
M1408|503515718|503443502
M1409|503515718|504368058
M1410|504628520|504409458
M1411|503418298|503497508
M1412|503418298|504303764
M1413|503634724|504107959
M1414|503543014|503546166
M1415|503254195|503608280
M1416|503254195|504386413
M1417|504295805|504337975
M1418|504617847|504580008
M1419|502425281|502529075
M1420|502458411|502479222
M1421|504637328|504995988
M1422|504637328|504583576
M1423|504003061|504169596
M1424|502948870|502984009
M1425|503644166|503497274
M1426|504711954|504718024
M1427|503637696|503540493
M1428|503381519|503803833
M1429|504944612|504297059
M1430|503217195|503695805
M1431|504184145|503907282
M1432|504184145|504308470
M1433|504456498|504766383
M1434|504243465|504365625
M1435|504243465|504173742
M1436|504049414|503898561
M1437|503067218|503526377
M1438|503329148|503225539
M1439|503737886|503844296
M1440|503764144|503784339
M1441|503694415|503723380
M1442|504700175|504649796
M1443|503956230|504026743
M1444|504049221|503897618
M1445|504049221|504306171
M1446|503853254|504163053
M1447|504526285|504530191
M1448|504194601|504032490
M1449|503505378|503796728
M1450|503446279|503842555
M1451|503585510|504817967
M1452|503585510|504179374
M1453|504078916|503497302
M1454|504078916|504311135
M1455|502656083|503108132
M1456|502920379|503497697
M1457|504875300|504877937
M1458|504531004|504455232
M1459|504039192|504344501
M1460|504231007|504163497
M1461|504581060|504503934
M1462|503867922|503834583
M1463|504004518|504055712
M1464|502782687|502760157
M1465|503296668|503922155
M1466|504524360|504302471
M1467|504126227|504846755
M1468|504126227|504042887
M1469|503388408|503761210
M1470|502882555|503438025
M1471|504441613|504310955
M1472|503229456|503603496
M1473|503411965|503792970
M1474|503383959|503572248
M1475|504049169|504002563
M1476|504049169|504307866
M1477|504274120|504255905
M1478|504658548|504789938
M1479|504658548|504629735
M1480|503206081|503497526
M1481|503206081|504296357
M1482|504432726|504430061
M1483|502869627|502932955
M1484|504240016|504155486
M1485|504240016|504911868
M1486|503297711|503353908
M1487|504179804|504337207
M1488|504058316|503984749
M1489|504388295|504404378
M1490|504122670|504179830
M1491|504030099|503994598
M1492|504005675|502635965
M1493|504647175|504759286
M1494|502776079|503573272
M1495|504073587|503904297
M1496|504666129|504583619
M1497|504907815|504878315
M1498|502643841|504076732
M1499|502643841|503991357
M1500|504078931|503905510
M1501|504835647|504545759
M1502|504819474|505001672
M1503|503718011|503281135
M1504|502610111|501041084
M1505|503076808|503688665
M1506|503389942|503191064
M1507|504442301|504296402
M1508|504530688|504528677
M1509|504207638|504357457
M1510|504041737|503901650
M1511|504888357|504850919
M1512|504345626|504373316
M1513|504975900|504998038
M1514|504932738|504307950
M1515|504115691|504068384
M1516|503355399|503428702
M1517|503585540|503798839
M1518|503585540|504301494
M1519|504050657|503929917
M1520|503931637|504068281
M1521|504848419|504941003
M1522|504517631|504284567
M1523|503246892|503350295
M1524|502688939|503023856
M1525|504234369|504116244
M1526|504022991|504545438
M1527|503801691|504142324
M1528|502543702|503346987
M1529|502543702|504874916
M1530|502544010|502641777
M1531|504553935|504682974
M1532|504041835|503895081
M1533|504041835|504303741
M1534|504556546|504283498
M1535|503921502|504063702
M1536|503889301|504021478
M1537|504495775|504376009
M1538|504495775|504376009
M1539|504640447|504266263
M1540|503720519|504207546
M1541|503281864|503897642
M1542|503569406|503534366
M1543|504918317|504932049
M1544|502931159|503802032
M1545|503402178|503468005
M1546|503586001|503568168
M1547|503586069|503541572
M1548|504134912|503909509
M1549|504970032|504037091
M1550|504095778|503916388
M1551|504095778|504307795
M1552|504176244|503901671
M1553|504176244|504324165
M1554|504937135|504694440
M1555|503779386|504333970
M1556|504254978|504379733
M1557|504875019|504396349
M1558|504605286|504579876
M1559|503214548|503500393
M1560|503214548|503901650
M1561|504896389|504301129
M1562|503630433|504025162
M1563|504205503|504191463
M1564|504278828|504354967
M1565|504976138|504709284
M1566|504838542|504930064
M1567|504951152|504775091
M1568|504862022|504930361
M1569|504592676|504742988
M1570|504137677|504026893
M1571|504137677|504032683
M1572|503315297|503507566
M1573|503315297|504308458
M1574|504049186|503898609
M1575|504049186|504302535
M1576|504063660|503507139
M1577|504063660|504307828
M1578|504063660|504306023
M1579|503229418|503907312
M1580|503229418|504310910
M1581|502934732|503537424
M1582|504106223|504043405
M1583|504106223|504579772
M1584|504106223|504579805
M1585|504195472|504222207
M1586|504652703|504629049
M1587|503204707|503497191
M1588|503204707|504302580
M1589|504951143|504301152
M1590|504167666|504035902
M1591|503471046|503489178
M1592|502778215|503291713
M1593|504478043|504306207
M1594|504050669|503925833
M1595|503259551|503371077
M1596|503259551|504219483
M1597|504532725|503951023
M1598|504379951|504736110
M1599|504443661|504311367
M1600|504186133|504122609
M1601|504449710|504708194
M1602|504449710|504311336
M1603|504005000|504241664
M1604|504407275|504393547
M1605|503834826|504139505
M1606|504759201|504322037
M1607|503720474|503638772
M1608|503720474|504685604
M1609|504478270|504307889
M1610|503873009|503953864
M1611|502946633|502893902
M1612|503582752|503771996
M1613|503634722|503597445
M1614|503671417|504022116
M1615|503230851|503317475
M1616|504468544|504297069
M1617|504498650|504131389
M1618|504165894|504138163
M1619|503401421|504818783
M1620|504442284|504302566
M1621|504563369|504600175
M1622|504231269|503927707
M1623|504412845|504727827
M1624|504059287|504210666
M1625|504530709|500189256
M1626|503144476|503453981
M1627|504417080|504872445
M1628|503433219|503890372
M1629|503836529|503876514
M1630|504390954|504231700
M1631|503662361|503740772
M1632|503835875|503926804
M1633|504933441|504712714
M1634|503471483|503641249
M1635|503471483|504631163
M1636|503804106|502255664
M1637|503804106|503988181
M1638|504486089|502643791
M1639|504051221|503972520
M1640|503224812|503385277
M1641|504495854|504303214
M1642|504401349|504856770
M1643|504476395|504302545
M1644|504260162|504639207
M1645|503589761|504552375
M1646|503589761|503582412
M1647|503669403|503553049
M1648|503669403|504549032
M1649|504896413|504296421
M1650|504168597|504161094
M1651|503001538|503380945
M1652|504468562|504556956
M1653|503321228|503412979
M1654|504660516|503922166
M1655|504211769|504100154
M1656|504495820|504297164
M1657|504495820|504297164
M1658|503650774|503526078
M1659|503995241|503924249
M1660|504449730|504307828
M1661|503314773|504176084
M1662|503022461|504323998
M1663|504918193|504884057
M1664|504391010|504614273
M1665|503873448|503889163
M1666|504495871|503901733
M1667|503468785|503856524
M1668|503391580|503509851
M1669|503391580|504303256
M1670|503565647|503577080
M1671|503565647|503865770
M1672|504297445|504306075
M1673|504495828|504296415
M1674|503637758|503498727
M1675|503637758|504297025
M1676|504101686|503907516
M1677|503461190|503672434
M1678|503812210|504084695
M1679|503418294|503507180
M1680|503418294|504311115
M1681|504932802|504718131
M1682|504046908|504349113
M1683|503681425|503786945
M1684|504811851|504883582
M1685|503241971|503901671
M1686|503602769|504787610
M1687|503602769|503919845
M1688|504724296|504746325
M1689|504122686|504171365
M1690|504462301|503680396
M1691|504478000|504306150
M1692|503911799|503956879
M1693|503661137|504531427
M1694|503661137|503507155
M1695|503644157|504605644
M1696|503644157|503500364
M1697|504441601|504306403
M1698|504449694|504311015
M1699|503226693|503035671
M1700|503883171|502138981
M1701|504601619|504611053
M1702|504042033|503916425
M1703|504042033|504303791
M1704|503587467|503886373
M1705|504918404|504629049
M1706|504600029|504579912
M1707|504600029|504884009
M1708|503778456|503787440
M1709|504619564|504579789
M1710|504345299|504397824
M1711|504403567|504689704
M1712|503589735|503488419
M1713|504909745|504634278
M1714|503062537|503455629
M1715|504976151|504722603
M1716|503774068|503866555
M1717|504604960|504374080
M1718|503866363|503946948
M1719|503862843|503926694
M1720|504468558|504296388
M1721|503476611|503495634
M1722|503856979|504170817
M1723|504449703|504302426
M1724|504106075|503995246
M1725|503967629|504276405
M1726|504445747|504321583
M1727|504399529|504803637
M1728|504392725|504697126
M1729|504579529|503853917
M1730|504443675|504310910
M1731|504605295|504875740
M1732|504605295|504629024
M1733|504507824|504575855
M1734|504081854|503905493
M1735|504478286|504297003
M1736|504601244|504577016
M1737|504112150|503907569
M1738|504112150|504296357
M1739|503471487|502163847
M1740|504943196|504712668
M1741|504931624|504731990
M1742|503454717|503323641
M1743|504049330|503905491
M1744|504203765|504766376
M1745|504886739|504000676
M1746|504577424|503698988
M1747|504842848|504676684
M1748|504922812|500189256
M1749|504936878|503216970
M1750|504220461|503633204
M1751|504220461|504029691
M1752|503225825|504862689
M1753|503225825|503551624
M1754|504262369|504538390
M1755|504934152|504707562
M1756|504919512|504892783
M1757|503585543|500189320
M1758|504930090|504741770
M1759|504932947|504722595
M1760|504902017|501028238
M1761|504932921|504725071
M1762|504932725|504719725
M1763|504886700|504777354
M1764|504673056|504845407
M1765|503953662|503952799
M1766|504934155|504708831
M1767|504574836|504303283
M1768|503798419|502994003
M1769|504970016|504708027
M1770|503996764|503889103
M1771|504933050|504707396
M1772|504153377|504487777
M1773|504932900|504718207
M1774|504933011|504718087
M1775|504931636|504722516
M1776|504219209|504301519
M1777|504030927|503905447
M1778|504530646|504637067
M1779|504220029|504198281
M1780|504965759|504718233
M1781|504404998|504481744
M1782|503286862|503386901
M1783|504039337|504011759
M1784|503663973|503865770
M1785|503663973|504568754
M1786|504943089|504725175
M1787|504425557|504124868
M1788|504298787|504325174
M1789|503739912|503929189
M1790|504965797|504719673
M1791|504970025|504718076
M1792|503637911|503507211
M1793|504599974|504579851
M1794|504599974|504905469
M1795|503978163|504510675
M1796|504933006|504708229
M1797|504185266|504213307
M1798|503663417|504057497
M1799|504033095|503900507
M1800|504033095|504708147
M1801|504254967|504209409
M1802|504473041|504582115
M1803|503530548|503635342
M1804|503833932|503698988
M1805|504468548|504297196
M1806|504241299|504194344
M1807|504727612|504822117
M1808|503834833|503968276
M1809|504929993|504716201
M1810|503290655|504326647
M1811|503955220|503874105
M1812|503366783|503493458
M1813|504967850|504718021
M1814|504965771|504718182
M1815|504929976|504712694
M1816|504441617|504296345
M1817|504443588|504308465
M1818|503496397|503797696
M1819|504029216|503916972
M1820|504029216|504307988
M1821|504030970|503995921
M1822|504929983|504741735
M1823|504449801|504296421
M1824|504443634|504297141
M1825|503644251|503288713
M1826|503644251|504375905
M1827|504956436|504725140
M1828|504576297|504308458
M1829|504942885|504732009
M1830|503629828|503497539
M1831|503629828|504306008
M1832|504971582|504708804
M1833|504932937|504719691
M1834|503965808|504180840
M1835|504517488|503853917
M1836|503558194|503527934
M1837|503661150|503603498
M1838|503661150|504297094
M1839|504960078|504707677
M1840|504106167|504026893
M1841|504442292|504375946
M1842|504533508|504443510
M1843|503575837|503825634
M1844|504487104|502924751
M1845|504998024|504718378
M1846|504998017|504714248
M1847|503579909|503552956
M1848|503798824|503895001
M1849|504930097|504707501
M1850|504103356|503896267
M1851|503554921|503556149
M1852|503654738|503853843
M1853|504931611|504709361
M1854|504442313|504297082
M1855|504037433|504722559
M1856|503856172|503961801
M1857|503644282|503521705
M1858|503644282|504301111
M1859|503617871|503786945
M1860|504971614|504708240
M1861|505001625|504716181
M1862|504819428|504805078
M1863|504579544|502143796
M1864|504101750|503898526
M1865|503805008|504322860
M1866|504934159|504709318
M1867|504029245|503907342
M1868|504029245|504719766
M1869|504956449|504712902
M1870|504960064|504719639
M1871|503644208|503540957
M1872|503644208|504301129
M1873|504033059|503898570
M1874|504933160|504709325
M1875|504966805|504843117
M1876|504933392|504707250
M1877|504073275|504032411
M1878|505011025|504707532
M1879|503717075|503842851
M1880|503717075|504270682
M1881|504652697|504579805
M1882|504599957|504579744
M1883|504599957|504871177
M1884|504612286|504634827
M1885|504106116|504043276
M1886|504106116|504579862
M1887|504035892|503905466
M1888|504095796|503905482
M1889|503902854|504273752
M1890|504033104|503907262
M1891|504231851|503291779
M1892|504930076|504709344
M1893|504388144|504365599
M1894|503572810|503785317
M1895|504532539|504467958
M1896|504468571|504301055
M1897|504468571|504707239
M1898|504886770|504771529
M1899|504883829|504629735
M1900|503804124|504284484
M1901|504915869|504933506
M1902|504348389|504667599
M1903|504538972|502171015
M1904|504400213|503961801
M1905|504081829|503916445
M1906|504155409|504606544
M1907|504041991|503898591
M1908|504933110|504719709
M1909|504033052|503896236
M1910|504033052|504732663
M1911|504956421|504727760
M1912|504272839|504114967
M1913|504629014|504619516
M1914|504629014|504619516
M1915|504967881|504707461
M1916|504952245|504757125
M1917|505022089|504741631
M1918|503661106|503608284
M1919|503661106|504303240
M1920|504937124|504828127
M1921|504275417|504249590
M1922|503781255|504179316
M1923|504917122|504453155
M1924|503993975|503947272
M1925|504095814|503901733
M1926|504456510|504829731
M1927|503862846|504765492
M1928|504357786|504163106
M1929|504041716|503916375
M1930|504579602|504634278
M1931|504069856|502591360
M1932|504026699|504659125
M1933|504449794|504303177
M1934|504447302|504307845
M1935|504096330|503992956
M1936|504096289|503776419
M1937|504044312|503862152
M1938|504029267|504375960
M1939|504433829|504470539
M1940|504443697|504307612
M1941|504180621|504624656
M1942|503774486|503792812
M1943|504049133|503907282
M1944|504095817|503995722
M1945|504834879|504666284
M1946|504303891|504553488
M1947|504524465|504438216
M1948|504524465|504438216
M1949|504041803|503897667
M1950|504699174|504744195
M1951|503960671|504107327
M1952|504447323|504303681
M1953|504405002|504241664
M1954|504182796|504378001
M1955|504112110|504409289
M1956|504682143|504313521
M1957|504690665|502240986
M1958|504982340|504755956
M1959|504532089|504631918
M1960|504919506|504871597
M1961|504447304|504306107
M1962|504101661|503925846
M1963|504101661|504302447
M1964|504049279|503898540
M1965|504049279|504741711
M1966|504478304|504443741
M1967|504478304|504721191
M1968|504495891|504306089
M1969|503978167|504529749
M1970|504168599|504166556
M1971|504505830|504419128
M1972|505026952|504725007
M1973|504495791|504452192
M1974|504075474|503792949
M1975|504636958|504549037
M1976|504592686|504594988
M1977|504951117|504671040
M1978|504188050|504845940
M1979|504998019|504739301
M1980|504915468|504349057
M1981|504461758|504468576
M1982|504496553|504419043
M1983|504496553|504723806
M1984|504345301|504373845
M1985|504622170|504802975
M1986|504495730|504428689
M1987|504495730|504428689
M1988|504478319|504419161
M1989|504478319|504723859
M1990|504997997|504729038
M1991|504617761|504911953
M1992|504478033|504442352
M1993|504956464|504901170
M1994|504571845|504442352
M1995|504571845|504731823
M1996|504970056|504764294
M1997|504505823|504416646
M1998|504505823|504741636
M1999|504525282|504452202
M2000|504525282|504732675
M2001|504502423|504452221
M2002|504461688|504442316
M2003|504461688|504723876
M2004|504998028|504731856
M2005|504276350|504273397
M2006|504960292|504714143
M2007|504211341|504224356
M2008|504960210|504666420
M2009|504453477|503803589
M2010|504478083|504438031
M2011|504505846|504438050
M2012|504505846|504723759
M2013|504918273|504871256
M2014|504260164|504523141
M2015|504963048|504724989
M2016|504241295|503542037
M2017|504965733|504739346
M2018|504496656|504419085
M2019|504496656|504723816
M2020|504502456|504428583
M2021|504502456|504739362
M2022|504478022|504428560
M2023|504478022|504452221
M2024|504530664|504363589
M2025|504461329|504442387
M2026|504366634|504346767
M2027|505004269|504729049
M2028|504461792|504418898
M2029|504997973|504729023
M2030|504439153|500189709
M2031|504960282|504833597
M2032|504360025|503844843
M2033|504524429|504442387
M2034|504524429|504729038
M2035|504441583|504441249
M2036|504441583|504739276
M2037|504461293|504452241
M2038|504461293|504721236
M2039|504502404|504418950
M2040|504502404|504732709
M2041|504530464|504428766
M2042|504530464|504739376
M2043|504524449|504442325
M2044|504524449|504934167
M2045|504533461|504565015
M2046|504965745|504721170
M2047|504997959|504741689
M2048|504415884|504930194
M2049|504524390|504438266
M2050|504442355|500790181
M2051|504502465|504438196
M2052|504819441|504805076
M2053|504502442|504428719
M2054|504918305|504875774
M2055|504620049|504659863
M2056|504899050|504850064
M2057|504951130|504806060
M2058|504918090|504883844
M2059|504461307|504452261
M2060|504461307|504725042
M2061|502527168|501646021
M2062|502374716|503560077
M2063|503490571|503645850
M2064|502874566|502894480
M2065|503895506|504026849
M2066|503706992|503709061
M2067|503673635|502143796
M2068|503779460|503659745
M2069|504050606|503972019
M2070|501872144|502063676
M2071|502455004|502680045
M2072|504059280|503998203
M2073|503355390|503843020
M2074|503467766|503543048
M2075|500896588|500924445
M2076|501023408|501356600
M2077|503860710|504115693
M2078|502215233|504119825
M2079|502485856|503544124
M2080|500186798|500189825
M2081|500771746|500996153
M2082|501513669|500824400
M2083|501609876|501425392
M2084|500881634|500816190
M2085|504043329|503918707
M2086|500835156|500466903
M2087|501132052|501356464
M2088|501129781|500189245
M2089|501488919|501392684
M2090|504042339|503984783
M2091|504043224|503985439
M2092|501160242|502325100
M2093|504043260|503969480
M2094|502445356|501026290
M2095|504043128|503985272
M2096|504043397|503922094
M2097|503239475|503162880
M2098|500337327|500189300
M2099|500399844|500188569
M2100|504419889|503976384
M2101|502785308|502736971
M2102|504043170|503974104
M2103|504445232|504431681
M2104|502034298|500188638
M2105|502137546|501641708
M2106|502763586|500189754
M2107|501101149|500834694
M2108|501618024|501500078
M2109|503633704|503604638
M2110|504416193|504394474
M2111|502300563|502101059
M2112|502445373|502453180
M2113|502505660|504331356
M2114|500577150|501734288
M2115|504416147|504212639
M2116|503635533|503604414
M2117|504308876|504215512
M2118|504579590|504397175
M2119|501129794|500922570
M2120|502813454|502855397
M2121|503624326|503605964
M2122|504012972|503975669
M2123|503292494|503216525
M2124|502813470|502889718
M2125|502813513|502915648
M2126|504401898|504350243
M2127|502776341|502631040
M2128|503610353|503973144
M2129|503996726|503355514
M2130|503012569|502966672
M2131|504396299|503973970
M2132|503292427|503282196
M2133|503250358|501721806
M2134|503779471|503040015
M2135|503610226|504260675
M2136|502813527|502691411
M2137|503807530|503381588
M2138|503292675|503282391
M2139|504396213|503615576
M2140|503249895|503372833
M2141|502290745|501944716
M2142|504183436|504053150
M2143|504198005|504222771
M2144|502369374|501876592
M2145|504257276|504250952
M2146|504184625|504016261
M2147|503694497|503550540
M2148|504936816|504528677
M2149|504220499|504045698
M2150|503457000|503552518
M2151|504449667|504633714
M2152|502813442|502656402
