AgencyName|AgencyGroup|OfficeName|TeamName|MatchType|MatchStatus|MatchOpenDate|MatchCloseDate|SurveyType|YOSScheduledDate|YOSCompletionDate|YOSCompletionType|YOSStatus|Q1|Q2Neg|Q3Neg|Q4Neg|Q5|Q6|SocAccept|Q1b|Q2b|Q3b|Q4b|Q5b|Q6b|SocAcceptB|SocAcceptPrcnt|Q7Neg|Q8|Q9|Q10Neg|Q11Neg|Q12|SchComp|Q7b|Q8b|Q9b|Q10b|Q11b|Q12b|SchCompB|SchCompPrcnt|Q13|Q14|Q15|EdExpect|Q13b|Q14b|Q15b|EdExpectb|EdExpectPrcnt|Q16|Q17|Q18|Q19|Grades|Q16b|Q17b|Q18b|Q19b|Gradesb|GradesPrcnt|Q20Neg|Q21Neg|Q22Neg|Q23Neg|Q24Neg|Q25Neg|Q26Neg|RiskAtt|Q20b|Q21b|Q22b|Q23b|Q24b|Q25b|Q26b|RiskAttb|RiskAttPrcnt|Q27|Q28|Q29|PTrust|Q27b|Q28b|Q29b|PTrustb|PTrustPrcnt|Q30Neg|Q31Neg|Truancy|Q30b|Q31b|Truancyb|TruancyPrcnt|Q32|SpAdult|Q32b|SpAdultb|SpAdultPrcnt|Q33Neg|JJustice|Q33b|JJusticeB|JJusticePrcnt|MatchSupportLevel|MatchReportSources|MatchClosureReasons|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildGrade|ChildLivingSituation|ChildIncomeLevel|ChildFamilyAssistance|ChildFreeReducedLunch|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|ChildPartKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolPartKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|MatchKey|MatchTypeKey|SiteTypeKey|MatchActivityKey|SiteKey|StatusKey|MatchSupportLevelKey|MatchReportSourceKey|ChildReportSourceKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|YOSSurveyKey|PriorBaselineYOSSurveyKey|YOSStatusKey|YOSCompletionTypeKey|SurveyTypeKey|CustodialAdultEmployerHash
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-08|NaT|Baseline|2014-11-25|2015-01-08|Complete|Done|4|3|4|2|4|4|3.5|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||25.9||1|1|1|1|M|Multi-race (Black & White)||13|Yes|Aunt|28031|6|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||51|28031|Masters Degree|Married|Real Estate: Realtor|28031|2|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020753|503654364|503656324|36|0|1|504076011|1|0|1|500799134|2||-2||2|1||500000294|-2||-2|0|4|||7438|1|||1|825549|-1|4|3|44|6178126991714892144
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-08|NaT|Followup|2016-01-08|2016-02-26|Declined|Late||||||||4|3|4|2|4|4|3.5|||||||||3|4|4|4|4|4|3.83||||||4|4|4|4|||||||5|5|5|4|4.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Green|||25.9||1|1|1|1|M|Multi-race (Black & White)||13|Yes|Aunt|28031|6|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||51|28031|Masters Degree|Married|Real Estate: Realtor|28031|2|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020753|503654364|503656324|36|0|1|504076011|1|0|1|500799134|2||-2||2|1||500000294|-2||-2|0|4|||7438|1|||1|839581|825549|4|1|45|6178126991714892144
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-08|NaT|Followup|2017-01-08|2017-02-20|Complete|Done|3|3|3|2|3|3|2.83|4|3|4|2|4|4|3.5|-19.14|3|4|3|3|3|3|3.17|3|4|4|4|4|4|3.83|-17.23|4|4|4|4|4|4|4|4|0|4|5|4|4|4.25|5|5|5|4|4.75|-10.53|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|3|3|3|4|4|4|4|-25|2|2|2|4|4|4|-50|2|2|2|2|0|4|4|4|4|0|Green|||25.9||1|1|1|1|M|Multi-race (Black & White)||13|Yes|Aunt|28031|6|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||51|28031|Masters Degree|Married|Real Estate: Realtor|28031|2|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020753|503654364|503656324|36|0|1|504076011|1|0|1|500799134|2||-2||2|1||500000294|-2||-2|0|4|||7438|1|||1|998525|825549|4|3|45|6178126991714892144
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-09|2017-01-27|Followup|2016-01-09|2016-02-29|Declined|Late||||||||4|1|4|1|4|4|3|||||||||2|4|4|2|3|4|3.17||||||4|4|4|4|||||||4|2|2|4|3||||||||||3|4|4|4|4|4|3|3.71||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Red||Child/Family: Lost contact with volunteer/agency|24.6||1|2|1|2|M|Black||15|No|Mother|28206|7|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|M|White||31|28205|Masters Degree|Single|Business|28262|8|0|Duke Energy|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500013781|503635533|503580712|31|0|1|503604414|1|0|1|500807416|2||-2||4|3|||-2||-2|0|4|||16705|3|||1|840080|667227|4|1|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-09|2017-01-27|Followup|2017-01-09|2017-01-13|Declined|Done||||||||4|1|4|1|4|4|3|||||||||2|4|4|2|3|4|3.17||||||4|4|4|4|||||||4|2|2|4|3||||||||||3|4|4|4|4|4|3|3.71||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Red||Child/Family: Lost contact with volunteer/agency|24.6||1|2|1|2|M|Black||15|No|Mother|28206|7|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|M|White||31|28205|Masters Degree|Single|Business|28262|8|0|Duke Energy|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500013781|503635533|503580712|31|0|1|503604414|1|0|1|500807416|2||-2||4|3|||-2||-2|0|4|||16705|3|||1|999472|667227|4|1|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-12|2015-08-31|Baseline|2014-09-02|2015-01-12|Complete|Done|4|2|3|2|1|2|2.33|||||||||1|4|4|2|1|4|2.67|||||||||3|4|4|3.67||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red||Child/Family: Moved|7.6||1|1|1|1|F|Multi-race (Black & White)||14|No|Mother|28217|7|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||49|28210|Masters Degree|Divorced|Education|28211|6|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503535105|503536977|36|0|2|504127300|1|0|2|500805104|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|789387|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-12|2016-04-18|Baseline|2014-12-18|2015-01-12|Complete|Done|1|3|3|4|3|2|2.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|3|4.25|||||||4|4|4|4|4|4|4|4||||||||||1|1|1|1||||||4|3|3.5|||||2|2||||4|4||||Green||Child: Family structure changed|15.2||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$40,000 to $44,999||No||Self|General Community||Match Support|M|White||30|28205|Bachelors Degree|Living w/ Significant Other|Finance: Banking|28217|3|4|Igniting Breakfast|Special Event|Big|General Community||Match Support|277|60|598|500000170|500021785|502107146|502107573|31|0|1|504090344|1|0|1|500804987|2||-2||4|1|||-2||-2|0|10|||17266|8|||1|834811|-1|4|3|44|7151546326379863072
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-12|2016-04-18|Followup|2016-01-12|2016-03-01|Declined|Late||||||||1|3|3|4|3|2|2.67|||||||||4|4|4|4|4|4|4||||||4|4|4|4|||||||5|4|5|3|4.25||||||||||4|4|4|4|4|4|4|4||||||1|1|1|1|||||4|3|3.5||||2|2||||4|4||Green||Child: Family structure changed|15.2||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$40,000 to $44,999||No||Self|General Community||Match Support|M|White||30|28205|Bachelors Degree|Living w/ Significant Other|Finance: Banking|28217|3|4|Igniting Breakfast|Special Event|Big|General Community||Match Support|277|60|598|500000170|500021785|502107146|502107573|31|0|1|504090344|1|0|1|500804987|2||-2||4|1|||-2||-2|0|10|||17266|8|||1|840420|834811|4|1|45|7151546326379863072
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-13|NaT|Baseline|2014-12-17|2015-01-13|Complete|Done|3|3|2|3|3|3|2.83|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|3|3|3|3.57||||||||||3|4|2|3||||||4|3|3.5|||||1|1||||4|4||||Yellow|PERL 2014-2016||25.8||1|1|1|1|F|Black||15|Yes|Mother|28212|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||25|28213|Bachelors Degree|Single|Retail: Mgt||0|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504076406|504078432|31|0|2|503831499|31|0|2|500807374|2||-2||2|2|500014681|500014681|-2|500014681|-2|0|5|||17159|12|||1|834438|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-13|NaT|Baseline|2015-01-07|2015-01-13|Complete|Done|3|2|4|2|3|3|2.83|||||||||2|3|3|3|3|4|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|||25.8||1|1|1|1|F|Black||16|No|Mother|28105|10|One Parent: Female|$35,000 to $39,999|Y|Yes|Other|Faith Organization|General Community||Match Support|F|Black||27|28227|Bachelors Degree|Single|Finance: Banking|29715|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|504090244|504092274|31|0|2|504121323|31|0|2|500806857|2||-2||2|1|||-2||-2|5635|9|||46|2|||1|839314|-1|4|3|44|2359037990929827326
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-13|NaT|Baseline|2015-01-07|2015-01-13|Complete|Done|4|3|3|3|4|4|3.5|||||||||2|4|4|3|3|4|3.33|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|2|2.5|||||1|1||||4|4||||Green|||25.8||1|1|1|1|M|Black||16|No|Mother|28227|8|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community||Match Support|M|White||30|28202|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|504034181|504036199|31|0|1|504053608|1|0|1|500806936|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|839397|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-13|NaT|Followup|2016-01-13|2016-01-31|Complete|Done|3|3|4|4|3|3|3.33|3|2|4|2|3|3|2.83|17.67|2|4|4|4|2|4|3.33|2|3|3|3|3|4|3|11|4|4|4|4|4|4|4|4|0|3|3|5|4|3.75|4|4|4|4|4|-6.25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|3|2.5|3|4|3.5|-28.57|2|2|2|2|0|4|4|4|4|0|Green|||25.8||1|1|1|1|F|Black||16|No|Mother|28105|10|One Parent: Female|$35,000 to $39,999|Y|Yes|Other|Faith Organization|General Community||Match Support|F|Black||27|28227|Bachelors Degree|Single|Finance: Banking|29715|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|504090244|504092274|31|0|2|504121323|31|0|2|500806857|2||-2||2|1|||-2||-2|5635|9|||46|2|||1|841070|839314|4|3|45|2359037990929827326
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-13|NaT|Followup|2016-01-13|2016-01-19|Complete|Done|4|3|3|3|3|3|3.17|4|3|3|3|4|4|3.5|-9.43|3|3|3|3|3|3|3|2|4|4|3|3|4|3.33|-9.91|4|4|4|4|4|4|4|4|0|5|4|4|4|4.25|4|4|5|4|4.25|0|4|4|4|4|4|3|3|3.71|4|4|4|4|4|4|3|3.86|-3.89|3|4|3|3.33|3|4|4|3.67|-9.26|4|2|3|3|2|2.5|20|2|2|1|1|100|4|4|4|4|0|Green|||25.8||1|1|1|1|M|Black||16|No|Mother|28227|8|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community||Match Support|M|White||30|28202|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|504034181|504036199|31|0|1|504053608|1|0|1|500806936|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|841097|839397|4|3|45|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-13|NaT|Followup|2016-01-13|2016-01-31|Complete|Done|3|3|3|3|3|3|3|3|3|2|3|3|3|2.83|6.01|3|4|3|3|3|3|3.17|3|4|3|3|3|3|3.17|0|4|4|3|3.67|4|4|4|4|-8.25|3|3|5|4|3.75|4|5|4|5|4.5|-16.67|4|4|4|4|4|4|3|3.86|4|4|4|4|3|3|3|3.57|8.12|3|4|3|3.33|3|4|2|3|11|3|3|3|4|3|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Yellow|PERL 2014-2016||25.8||1|1|1|1|F|Black||15|Yes|Mother|28212|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||25|28213|Bachelors Degree|Single|Retail: Mgt||0|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504076406|504078432|31|0|2|503831499|31|0|2|500807374|2||-2||2|2|500014681|500014681|-2|500014681|-2|0|5|||17159|12|||1|841104|834438|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-13|NaT|Followup|2017-01-13|2017-01-12|Complete|Done|3|4|4|4|3|3|3.5|3|2|4|2|3|3|2.83|23.67|3|4|4|4|4|4|3.83|2|3|3|3|3|4|3|27.67|4|4|4|4|4|4|4|4|0|3|5|5|5|4.5|4|4|4|4|4|12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|2|3|3|4|3.5|-14.29|2|2|2|2|0|4|4|4|4|0|Green|||25.8||1|1|1|1|F|Black||16|No|Mother|28105|10|One Parent: Female|$35,000 to $39,999|Y|Yes|Other|Faith Organization|General Community||Match Support|F|Black||27|28227|Bachelors Degree|Single|Finance: Banking|29715|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|504090244|504092274|31|0|2|504121323|31|0|2|500806857|2||-2||2|1|||-2||-2|5635|9|||46|2|||1|989317|839314|4|3|45|2359037990929827326
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-18|NaT|Followup|2016-01-18|2016-01-27|Complete|Done|1|1|1|1|4|4|2|||||||||2|4|4|1|1|4|2.67|||||||||4|4|4|4||||||4|4|5|2|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||25.6||1|1|1|1|F|Black||10|Yes|Mother|28208|5|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||27|29730|Bachelors Degree|Married|Finance|28277|3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504115691|504117725|31|0|2|504068384|1|0|2|500807126|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||17159|12|||1|902579||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-18|NaT|Followup|2017-01-18|2017-01-18|Complete|Done|4|1|1|1|2|2|1.83|||||||||2|4|3|1|1|3|2.33|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||25.6||1|1|1|1|F|Black||10|Yes|Mother|28208|5|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||27|29730|Bachelors Degree|Married|Finance|28277|3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504115691|504117725|31|0|2|504068384|1|0|2|500807126|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||17159|12|||1|987781||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-23|NaT|Baseline|2015-01-13|2015-01-23|Complete|Done|4|1|4|4|4|4|3.5|||||||||4|4|4|4|3|4|3.83|||||||||1|3|1|1.67||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|3|2|||||1|1||||4|4||||Green|PERL 2014-2016||25.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||37|28215|Masters Degree|Married|Finance: Banking|28262|15|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503224764|503226552|31|0|1|504130394|31|0|1|500807724|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|840786|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-23|NaT|Followup|2016-01-23|2016-02-28|Declined|Done||||||||4|1|4|4|4|4|3.5|||||||||4|4|4|4|3|4|3.83||||||1|3|1|1.67|||||||4|4|4|4|4||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||1|3|2||||1|1||||4|4||Green|PERL 2014-2016||25.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||37|28215|Masters Degree|Married|Finance: Banking|28262|15|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503224764|503226552|31|0|1|504130394|31|0|1|500807724|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|844078|840786|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-23|NaT|Followup|2017-01-23|2017-02-28|Declined|Done||||||||4|1|4|4|4|4|3.5|||||||||4|4|4|4|3|4|3.83||||||1|3|1|1.67|||||||4|4|4|4|4||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||1|3|2||||1|1||||4|4||Green|PERL 2014-2016||25.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||37|28215|Masters Degree|Married|Finance: Banking|28262|15|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503224764|503226552|31|0|1|504130394|31|0|1|500807724|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|999038|840786|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-26|2016-05-10|Baseline|2015-01-23|2015-01-26|Complete|Done|3|4|4|3|4|4|3.67|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green||Child/Family: Moved|15.4||1|1|1|1|M|Multi-race (Black & White)||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||30|28203|Masters Degree|Single|Finance: Banking|28262|4|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504054633|504056657|36|0|1|504068503|1|0|1|500809809|2||-2||4|1|||-2||-2|0|4|||17159|12|||1|844194|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-26|2016-05-10|Followup|2016-01-26|2016-01-26|Complete|Done|3|3|4|3|3|3|3.17|3|4|4|3|4|4|3.67|-13.62|4|4|3|4|3|4|3.67|4|4|4|4|2|4|3.67|0|4|4|4|4|4|4|4|4|0|4|4|5|3|4|5|5|5|5|5|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|2|2|2|4|2|3|-33.33|1|1|2|2|-50|4|4|4|4|0|Green||Child/Family: Moved|15.4||1|1|1|1|M|Multi-race (Black & White)||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||30|28203|Masters Degree|Single|Finance: Banking|28262|4|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504054633|504056657|36|0|1|504068503|1|0|1|500809809|2||-2||4|1|||-2||-2|0|4|||17159|12|||1|844821|844194|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-26|2016-05-04|Followup|2016-01-26|2016-04-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Feels incompatible with volunteer|15.2||2|2|1|1|F|Black||11|No|Mother|28217|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||24|28213||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500021785|504126227|504128262|31|0|2|504042887|31|0|2|500807321|2||-2||4|1||500007920, 500011315, 500011316|-2||-2|0|4|||46|2|||1|856465||4|0|45|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-26|NaT|Followup|2016-01-26|2016-01-23|Complete|Done|1|4|4|2|3|3|2.83|3|4|2|2|3|4|3|-5.67|4|4|4|4|4|4|4|2|3|3|4|3|4|3.17|26.18|4|1|4|3|3|3|3|3|0|4|4|3|4|3.75|3|4|3|3|3.25|15.38|4|4|4|4|4|4|4|4|4|4|4|4|3|4|4|3.86|3.63|4|4|4|4|3|4|3|3.33|20.12|2|4|3|1|4|2.5|20|2|2|2|2|0|4|4|4|4|0|Green|||25.3||2|2|1|1|F|Black||14|No|Mother|28206|8|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||30|28205|Bachelors Degree|Single|Human Services|28203|1|2|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|503816186|501097065|31|0|2|504090792|1|0|2|500807024|2||-2||2|1|||-2||-2|0|10|||130|1|||1|844734|745502|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-26|NaT|Followup|2016-01-26|2016-04-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||25.3||3|3|2|2|F|Black||11|No|Mother|28216|2|One Parent: Female|Unknown||Yes|TV|Media|General Community||Match Support|F|Black||48|28203|Bachelors Degree|Married|Business: Mgt, Admin|28202|1|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502324604|502325039|31|0|2|502657850|31|0|2|500808029|2||-2||2|1|||-2||-2|56|1|||7464|9|||1|844951||4|0|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-27|2016-11-09|Baseline|2014-09-19|2015-01-27|Complete|Done|3|3|4|3|2|3|3|||||||||3|3|2|2|3|3|2.67|||||||||4|3|3|3.33||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|3|3||||||4|4|4|||||1|1||||4|4||||Red|PERL 2014-2016|Child: Lost interest|21.4||1|1|4|5|F|White||14|No|Mother|28025|8|One Parent: Female|$35,000 to $39,999||No||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|277|60|598|500000170|500020753|503923436|503925443|1|0|2|501306527|1|0|2|500806777|2||-2||4|3|500014681|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||7464|9|||1|793984|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-27|2016-11-09|Followup|2016-01-27|2016-01-22|Complete|Done|3|2|3|4|3|3|3|3|3|4|3|2|3|3|0|2|4|3|4|2|3|3|3|3|2|2|3|3|2.67|12.36|4|4|4|4|4|3|3|3.33|20.12|3|3|5|5|4|4|4|4|5|4.25|-5.88|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|3|2|2.67|2|4|3|3|-11|4|2|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Red|PERL 2014-2016|Child: Lost interest|21.4||1|1|4|5|F|White||14|No|Mother|28025|8|One Parent: Female|$35,000 to $39,999||No||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|277|60|598|500000170|500020753|503923436|503925443|1|0|2|501306527|1|0|2|500806777|2||-2||4|3|500014681|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||7464|9|||1|845299|793984|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-27|NaT|Followup|2016-01-27|2016-02-04|Complete|Done|3|3|3|2|3|3|2.83|3|3|2|2|4|3|2.83|0|2|2|3|2|2|3|2.33|2|3|3|3|4|3|3|-22.33|4|4|4|4|4|4|4|4|0|1|3|1|1|1.5|3|4|3|2|3|-50|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|2|2.67|4|4|4|4|-33.25|2|2|2|3|3|3|-33.33|2|2|2|2|0|4|4|4|4|0|Yellow|PERL 2014-2016||25.3||2|2|1|1|F|Hispanic|Other South American|14|No|Mother|28212|8|Two Parent|Unknown||Yes|Big|Neighbor/Friend|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|Hispanic||26|28215|Bachelors Degree|Single|Student: College||0|0|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|277|60|598|500000170|500020753|502215233|502215660|3|15|2|504119825|3|0|2|500808734|2||-2||2|2|500014681|500011312, 500014681|-2|500000294, 500014681|-2|6854|8|||7464|9|||1|845417|645412|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-27|NaT|Followup|2016-01-27|2016-03-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||25.3||1|1|1|1|M|Black||10|No|Mother|28262|4|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Tech: Engineer|28027|3|11|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|503801691|503803668|31|0|1|504142324|1|0|1|500808169|2||-2||2|1|||-2|500000294|-2|0|10|||17159|12|||1|910628||4|1|45|386356889061704511
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-28|2015-03-05|Baseline|2015-01-26|2015-01-28|Complete|Done|4|3|2|3|3|4|3.17|||||||||3|4|3|2|2|4|3|||||||||4|4|4|4||||||3|5|4|4|4|||||||3|4|4|4|4|3|3|3.57||||||||||3|3|4|3.33||||||2|3|2.5|||||1|1||||4|4||||Green||Child: Lost interest|1.2||1|1|1|1|F|Black||15|No|Mother|28273|8|One Parent: Male|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|Black||37|28273|Masters Degree|Single|Business|29715|3|0|Current/Previous Big|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500013781|504174131|504143662|31|0|2|503997551|31|0|2|500810212|2||-2||4|1|||-2||-2|0|4|||17159|12|||1|845041|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-28|2017-02-28|Baseline|2015-01-28|2015-01-28|Complete|Done|4|2|4|1|4|4|3.17|||||||||2|4|4|1|2|4|2.83|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|25||1|1|1|1|M|Black||11|No|GrandMother|28215|1|One Parent: Female|$35,000 to $39,999|Y|Yes||School|General Community||Enrollment|M|White||26|28205|Bachelors Degree|Single|Business: Mgt, Admin|28205|1|7|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020753|503853254|503855248|31|0|1|504163053|1|0|1|500809956|2||-2||4|3|||-2|500000294|-2|0|4|||17159|12|||1|845753|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-28|2017-02-28|Followup|2016-01-28|2016-03-28|Declined|Late||||||||4|2|4|1|4|4|3.17|||||||||2|4|4|1|2|4|2.83||||||4|4|4|4|||||||3|4|3|4|3.5||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|2|2||||2|2||||4|4||Red||Volunteer: Lost contact with child/agency|25||1|1|1|1|M|Black||11|No|GrandMother|28215|1|One Parent: Female|$35,000 to $39,999|Y|Yes||School|General Community||Enrollment|M|White||26|28205|Bachelors Degree|Single|Business: Mgt, Admin|28205|1|7|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020753|503853254|503855248|31|0|1|504163053|1|0|1|500809956|2||-2||4|3|||-2|500000294|-2|0|4|||17159|12|||1|845756|845753|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-28|2017-02-28|Followup|2017-01-28|2017-02-02|Complete|Done|2|4|4|4|4|4|3.67|4|2|4|1|4|4|3.17|15.77|2|3|4|4|2|4|3.17|2|4|4|1|2|4|2.83|12.01|4|4|4|4|4|4|4|4|0|4|5|5|3|4.25|3|4|3|4|3.5|21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|2|2|2|100|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|25||1|1|1|1|M|Black||11|No|GrandMother|28215|1|One Parent: Female|$35,000 to $39,999|Y|Yes||School|General Community||Enrollment|M|White||26|28205|Bachelors Degree|Single|Business: Mgt, Admin|28205|1|7|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020753|503853254|503855248|31|0|1|504163053|1|0|1|500809956|2||-2||4|3|||-2|500000294|-2|0|4|||17159|12|||1|1007671|845753|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-29|2016-05-03|Baseline|2013-12-05|2015-01-28|Complete|Done|3|4|4|3|4|3|3.5|||||||||3|3|3|3|3|4|3.17|||||||||4|4|4|4||||||3|3|3|3|3|||||||3|4|4|4|2|3|2|3.14||||||||||3|4|3|3.33||||||3|3|3|||||1|1||||4|4||||Green||Child: Lost interest|15.1||1|1|1|1|F|Black||16|No|Mother|28212|8|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|F|Black||26|28213|Bachelors Degree|Single|Finance|28269|2|1|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500021785|503441463|501290021|31|0|2|504122275|31|0|2|500810468|2||-2||4|1|||-2||-2|0|4|||130|1|||1|685875|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-01-29|2016-05-03|Followup|2016-01-29|2016-03-28|Declined|Late||||||||3|4|4|3|4|3|3.5|||||||||3|3|3|3|3|4|3.17||||||4|4|4|4|||||||3|3|3|3|3||||||||||3|4|4|4|2|3|2|3.14||||||3|4|3|3.33|||||3|3|3||||1|1||||4|4||Green||Child: Lost interest|15.1||1|1|1|1|F|Black||16|No|Mother|28212|8|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|F|Black||26|28213|Bachelors Degree|Single|Finance|28269|2|1|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500021785|503441463|501290021|31|0|2|504122275|31|0|2|500810468|2||-2||4|1|||-2||-2|0|4|||130|1|||1|846129|685875|4|1|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-30|NaT|Baseline|2015-01-22|2015-01-30|Complete|Done|4|1|3|2|3|4|2.83|||||||||2|2|2|3|2|2|2.17|||||||||3|3|3|3||||||2|3|4|5|3.5|||||||4|4|4|4|3|4|3|3.71||||||||||3|3|2|2.67||||||3|1|2|||||2|2||||4|4||||Green|||25.2||1|1|1|1|F|Hispanic|Other South American|16|No|Mother|28215|7|Two Parent|$10,000 to $14,999|Y|Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||30|28211|Masters Degree|Married|Tech: Support, Writing|28202|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020753|503860710|503862704|3|15|2|504115693|1|0|2|500809450|2||-2||2|1||500011312|-2||-2|0|10|||17159|12|||1|843664|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-30|NaT|Followup|2016-01-30|2016-03-14|Declined|Done||||||||4|1|3|2|3|4|2.83|||||||||2|2|2|3|2|2|2.17||||||3|3|3|3|||||||2|3|4|5|3.5||||||||||4|4|4|4|3|4|3|3.71||||||3|3|2|2.67|||||3|1|2||||2|2||||4|4||Green|||25.2||1|1|1|1|F|Hispanic|Other South American|16|No|Mother|28215|7|Two Parent|$10,000 to $14,999|Y|Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||30|28211|Masters Degree|Married|Tech: Support, Writing|28202|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020753|503860710|503862704|3|15|2|504115693|1|0|2|500809450|2||-2||2|1||500011312|-2||-2|0|10|||17159|12|||1|847095|843664|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-31|NaT|Baseline|2015-01-21|2015-01-31|Complete|Done|4|2|4|3|3|4|3.33|||||||||1|3|3|1|2|2|2|||||||||4|4|4|4||||||3|4|2|2|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||4|2|3|||||2|2||||4|4||||Green|PERL 2014-2016||25.2||1|1|1|1|M|Black||13|No|Mother|28105|6|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||28|28105|Bachelors Degree|Single|Business: Human Resources|28204|1|2|Other|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503413169|503415024|31|0|1|504092153|1|0|1|500809276|2||-2||2|1|500014681|500014681|-2|500014681|-2|34|2|||7671|13|||1|843357|-1|4|3|44|3714886275549507192
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-31|NaT|Followup|2016-01-31|2016-01-30|Complete|Done|3|1|2|4|1|3|2.33|||||||||2|3|3|2|1|3|2.33|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||25.2||2|2|1|1|F|White||11|No|Father|28081|4|One Parent: Male|Unknown||Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||32|28226|Bachelors Degree|Married|Business: Mgt, Admin|10006|1|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503634724|503636659|1|0|2|504107959|1|0|2|500809650|2||-2||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||17159|12|||1|847217||4|3|45|1786514887916898235
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-31|NaT|Followup|2016-01-31|2016-04-16|Expired|Late||||||||4|2|4|3|3|4|3.33|||||||||1|3|3|1|2|2|2||||||4|4|4|4|||||||3|4|2|2|2.75||||||||||4|4|4|4|4|4|3|3.86||||||3|4|2|3|||||4|2|3||||2|2||||4|4||Green|PERL 2014-2016||25.2||1|1|1|1|M|Black||13|No|Mother|28105|6|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||28|28105|Bachelors Degree|Single|Business: Human Resources|28204|1|2|Other|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503413169|503415024|31|0|1|504092153|1|0|1|500809276|2||-2||2|1|500014681|500014681|-2|500014681|-2|34|2|||7671|13|||1|847222|843357|4|0|45|3714886275549507192
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-01-31|NaT|Followup|2017-01-31|2017-02-07|Complete|Done|4|1|2|1|1|3|2|||||||||1|4|3|2|1|3|2.33|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|3|4|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||25.2||2|2|1|1|F|White||11|No|Father|28081|4|One Parent: Male|Unknown||Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||32|28226|Bachelors Degree|Married|Business: Mgt, Admin|10006|1|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503634724|503636659|1|0|2|504107959|1|0|2|500809650|2||-2||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||17159|12|||1|989003||4|3|45|1786514887916898235
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-06|2016-08-08|Baseline|2015-01-23|2015-02-06|Complete|Done|2|1|1|1|4|1|1.67|||||||||1|3|4|4|4|4|3.33|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|PERL 2014-2016|Child: Severity of challenges|18||1|1|1|1|M|White||11|No|Mother|28081|3|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Hispanic||31|28083|Some College|Married|Business: Mgt, Admin||14|3|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504059549|504061573|1|0|1|504109643|3|0|2|500809931|2||-2||4|3|500014681|500014681, 500016374|-2|500014681, 500016374|-2|0|5|||46|2|||1|844355|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-06|2016-08-08|Followup|2016-02-06|2016-02-29|Complete|Done|4|2|2|1|1|1|1.83|2|1|1|1|4|1|1.67|9.58|1|3|3|1|1|2|1.83|1|3|4|4|4|4|3.33|-45.05|4|4|4|4|4|4|4|4|0|2|4|1|5|3|5|5|5|5|5|-40|4|4|4|4|4|4|2|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|4|4|4|4|4|4|0|2|3|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Red|PERL 2014-2016|Child: Severity of challenges|18||1|1|1|1|M|White||11|No|Mother|28081|3|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Hispanic||31|28083|Some College|Married|Business: Mgt, Admin||14|3|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504059549|504061573|1|0|1|504109643|3|0|2|500809931|2||-2||4|3|500014681|500014681, 500016374|-2|500014681, 500016374|-2|0|5|||46|2|||1|849404|844355|4|3|45|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-06|NaT|Baseline|2015-01-29|2015-02-06|Complete|Done|3|4|3|2|4|3|3.17|||||||||2|2|3|2|3|2|2.33|||||||||4|4|4|4||||||5|2||1||||||||4|4|4|4|4|4|4|4||||||||||2|3|1|2||||||4|2|3|||||2|2||||4|4||||Green|PERL 2014-2016||25||1|1|1|1|M|Black||16|No|Mother|28205|9|One Parent: Female|$10,000 to $14,999|Y|Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|White||36|28269|Bachelors Degree|Married|Self-Employed, Entrepreneur|28269|7|5|Other|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504063426|504065453|31|0|1|504152304|1|0|1|500810827|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|56|1|||7671|13|||1|846141|-1|4|3|44|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-06|NaT|Followup|2016-02-06|2016-04-22|Expired|Late||||||||3|4|3|2|4|3|3.17|||||||||2|2|3|2|3|2|2.33||||||4|4|4|4|||||||5|2||1|||||||||||4|4|4|4|4|4|4|4||||||2|3|1|2|||||4|2|3||||2|2||||4|4||Green|PERL 2014-2016||25||1|1|1|1|M|Black||16|No|Mother|28205|9|One Parent: Female|$10,000 to $14,999|Y|Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|White||36|28269|Bachelors Degree|Married|Self-Employed, Entrepreneur|28269|7|5|Other|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504063426|504065453|31|0|1|504152304|1|0|1|500810827|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|56|1|||7671|13|||1|849206|846141|4|0|45|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-09|NaT|Baseline|2015-01-22|2015-02-09|Complete|Done|2|4|4|2|1|3|2.67|||||||||2|4|4|2|2|3|2.83|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green|||24.9||1|1|1|1|F|Black||17|No|Mother|28217|8|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Black||24|28273|Some College|Single|Finance: Accountant|28226|6|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|504169896|504172004|31|0|2|503987952|31|0|2|500809606|2||-2||2|1||500014681|-2||-2|0|4|||46|2|||1|843833|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-09|NaT|Followup|2016-02-09|2016-03-28|Declined|Late||||||||2|4|4|2|1|3|2.67|||||||||2|4|4|2|2|3|2.83||||||4|4|4|4|||||||3|4|3|4|3.5||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||3|3|3||||2|2||||4|4||Green|||24.9||1|1|1|1|F|Black||17|No|Mother|28217|8|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Black||24|28273|Some College|Single|Finance: Accountant|28226|6|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|504169896|504172004|31|0|2|503987952|31|0|2|500809606|2||-2||2|1||500014681|-2||-2|0|4|||46|2|||1|849673|843833|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-13|2015-11-30|Baseline|2015-01-20|2015-02-13|Complete|Done|4|2|4|3|3|4|3.33|||||||||2|3|3|2|3|3|2.67|||||||||3|3|3|3||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||1|3|1|1.67||||||4|3|3.5|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|9.5||1|1|1|1|M|Black||16|No|Mother|28212|8|One Parent: Female|$35,000 to $39,999||Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|White||57|28226|Some College|Single|Business: Sales|28134|10|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|504129007|504131049|31|0|1|504137446|1|0|1|500809001|2||-2||4|3|500014681|500014681|-2|500014681|-2|56|1|||17159|12|||1|842899|-1|4|3|44|2197933814735019388
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-17|2015-09-04|Baseline|2015-02-05|2015-02-17|Complete|Done|4|1|4|2|4|4|3.17|||||||||3|4|3|4|3|4|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|1|3.57||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Lost contact with child/agency|6.5||1|1|1|1|M|Black||12|No|Mother|28216|4|One Parent: Female|$45,000 to $49,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||28|28214|Some College|Single|Transport: Driver||0|1|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|504065282|504067309|31|0|1|504168627|31|0|1|500812249|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|4|||46|2|||1|848860|-1|4|3|44|139697663694671798
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-17|2016-04-18|Followup|2016-02-17|2016-04-01|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||3|3||||Red|PERL 2014-2016|Volunteer: Moved|14||1|1|1|1|F|White||10|No|Mother|28078|3|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|PERL 2014-2016|Enrollment|F|White||38|28031|Some College|Single|Real Estate: Realtor|28031|8|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|504134912|504136949|1|0|2|503909509|1|0|2|500813035|2||-2||4|3|500014681|500014681|-2|500014681|-2|0|4|||46|2|||1|916459||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-17|NaT|Baseline|2014-12-18|2015-02-17|Complete|Done|4|4|4|4|4|4|4|||||||||2|2|4|4|2|4|3|||||||||4|3|4|3.67||||||3|3|3|2|2.75|||||||2|4|4|4|3|1|3|3||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||24.6||1|1|1|1|M|Black||16|No|Mother|28208|9|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||45|28273|Masters Degree|Married|Finance: Banking|28269|0|1|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|502552947|502553400|31|0|1|503881539|31|0|1|500804943|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|834754|-1|4|3|44|427143067147514567
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-17|NaT|Followup|2016-02-17|2016-05-03|Expired|Late||||||||4|4|4|4|4|4|4|||||||||2|2|4|4|2|4|3||||||4|3|4|3.67|||||||3|3|3|2|2.75||||||||||2|4|4|4|3|1|3|3||||||4|4|4|4|||||1|4|2.5||||2|2||||4|4||Green|PERL 2014-2016||24.6||1|1|1|1|M|Black||16|No|Mother|28208|9|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||45|28273|Masters Degree|Married|Finance: Banking|28269|0|1|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|502552947|502553400|31|0|1|503881539|31|0|1|500804943|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|851957|834754|4|0|45|427143067147514567
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-23|2017-02-28|Followup|2016-02-23|2016-03-31|Complete|Done|2|2|2|2|3|3|2.33|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||2|2|2|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|24.2||1|1|1|1|M|Multi-race (Black & White)||10|Yes|Mother|28204|1|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||26|28216|Bachelors Degree|Single|Tech: Engineer|28078|0|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503812210|503814187|36|0|1|504084695|1|0|1|500810906|2||-2||4|2|||-2||-2|0|10|||46|2|||1|991756||4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-24|NaT|Baseline|2014-09-26|2015-02-24|Complete|Done|3|4|4|4|4|3|3.67|||||||||2|4|2|4|4|4|3.33|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||1|1||||4|4||||Green|PERL 2014-2016||24.4||1|1|1|1|M|Black||12|No|Mother|28216|5|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||50|28211|Juris Doctorate (JD)|Married|Law: Lawyer|28211|17|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|503533041|503534897|31|0|1|504183712|1|0|1|500813495|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||7496|10|||1|796339|-1|4|3|44|1786514887916898235
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-24|NaT|Baseline|2015-02-18|2015-02-24|Complete|Done|3|2|1|1|3|2|2|||||||||1|4|1|1|2|1|1.67|||||||||4|2|2|2.67||||||2|3|3|5|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016||24.4||1|1|1|1|F|Black||12|Yes|Mother|28217|6|One Parent: Female|$20,000 to $24,999||No|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||28|28205|Bachelors Degree|Single|Journalist/Media|28202|4|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504171035|504173143|31|0|2|504150234|1|0|2|500814425|2||-2||2|1|500014681|500014681|-2|500014681|-2|34|2|||46|2|||1|852645|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-24|NaT|Followup|2016-02-24|2016-02-23|Complete|Done|4|4|1|4|4|1|3|3|2|1|1|3|2|2|50|1|4|4|1|1|3|2.33|1|4|1|1|2|1|1.67|39.52|4|4|4|4|4|2|2|2.67|49.81|3|3|3|4|3.25|2|3|3|5|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|1|3|2|3|3|3|-33.33|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||24.4||1|1|1|1|F|Black||12|Yes|Mother|28217|6|One Parent: Female|$20,000 to $24,999||No|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||28|28205|Bachelors Degree|Single|Journalist/Media|28202|4|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504171035|504173143|31|0|2|504150234|1|0|2|500814425|2||-2||2|1|500014681|500014681|-2|500014681|-2|34|2|||46|2|||1|854312|852645|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-24|NaT|Followup|2016-02-24|2016-04-19|Declined|Late||||||||3|4|4|4|4|3|3.67|||||||||2|4|2|4|4|4|3.33||||||4|4|4|4|||||||4|3|3|3|3.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||3|3|3||||1|1||||4|4||Green|PERL 2014-2016||24.4||1|1|1|1|M|Black||12|No|Mother|28216|5|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||50|28211|Juris Doctorate (JD)|Married|Law: Lawyer|28211|17|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|503533041|503534897|31|0|1|504183712|1|0|1|500813495|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||7496|10|||1|854688|796339|4|1|45|1786514887916898235
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-24|NaT|Followup|2017-02-24|2017-02-22|Complete|Done|4|4|4|4|3|3|3.67|3|2|1|1|3|2|2|83.5|2|4|3|2|4|4|3.17|1|4|1|1|2|1|1.67|89.82|4|4|4|4|4|2|2|2.67|49.81|3|2|2|2|2.25|2|3|3|5|3.25|-30.77|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|3|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||24.4||1|1|1|1|F|Black||12|Yes|Mother|28217|6|One Parent: Female|$20,000 to $24,999||No|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||28|28205|Bachelors Degree|Single|Journalist/Media|28202|4|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504171035|504173143|31|0|2|504150234|1|0|2|500814425|2||-2||2|1|500014681|500014681|-2|500014681|-2|34|2|||46|2|||1|997409|852645|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-26|2016-10-31|Baseline|2014-08-26|2015-02-26|Complete|Done|3|2|3|2|2|4|2.67|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red||Child/Family: Moved|20.1||1|1|1|1|M|Black||12|No|Mother|28269|5|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|M|White||34|28078|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28078|1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503884921|503876064|31|0|1|504160910|1|0|1|500814243|2||-2||4|3|||-2||-2|0|10|||46|2|||1|787794|-1|4|3|44|3501831218874457455
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-26|2017-01-12|Baseline|2015-02-22|2015-02-26|Complete|Done|4|4|3|2|4|4|3.5|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||1|5|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Time constraint|22.5||1|1|1|1|F|Black||12|No|Mother|28213|5|One Parent: Female|$45,000 to $49,999||Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Enrollment|F|Black||21|28269|Some College|Single|Business: Sales|28269|0|5|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|504038255|504040273|31|0|2|504034443|31|0|2|500814943|2||-2||4|1|500014681|500014681|-2|500014681|-2|34|2|||46|2|||1|853694|-1|4|3|44|8408514790530965815
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-26|2017-02-27|Followup|2016-02-26|2016-03-28|Complete|Done|4|4|4|4|4|4|4|3|2|2|2|3|3|2.5|60|2|4|3|2|4|3|3|3|4|3|4|1|2|2.83|6.01|4|4|4|4|4|4|4|4|0|3|3|2|3|2.75|3|3|4|5|3.75|-26.67|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|3|3.86|-3.89|4|4|4|4|4|4||||3|1|2|3|2|2.5|-20|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Time constraint|24||2|2|1|1|F|Black||14|No|Mother|28215|3|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||42|28216|Associate Degree|Married|Business: Clerical|28202|8|0|Duke Energy|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500013781|502875279|502876679|31|0|2|504151222|31|0|2|500815521|2||-2||4|3|||-2||-2|0|10|||16705|3|||1|855238|406736|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-26|2016-10-31|Followup|2016-02-26|2016-04-08|Complete|Done|3|2|3|3|3|3|2.83|3|2|3|2|2|4|2.67|5.99|2|3|3|3|3|4|3|2|4|3|3|2|3|2.83|6.01|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|3|3|3|3|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|4|4|4|4|-25|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Red||Child/Family: Moved|20.1||1|1|1|1|M|Black||12|No|Mother|28269|5|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|M|White||34|28078|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28078|1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503884921|503876064|31|0|1|504160910|1|0|1|500814243|2||-2||4|3|||-2||-2|0|10|||46|2|||1|855256|787794|4|3|45|3501831218874457455
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-26|2017-01-12|Followup|2016-02-26|2016-02-25|Complete|Done|3|3|3|3|3|2|2.83|4|4|3|2|4|4|3.5|-19.14|2|4|2|3|3|2|2.67|2|4|4|2|2|4|3|-11|4|4|4|4|4|4|4|4|0|1|5|3|2|2.75|1|5|4|5|3.75|-26.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|2|4|3|4|3|3.5|-14.29|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016|Volunteer: Time constraint|22.5||1|1|1|1|F|Black||12|No|Mother|28213|5|One Parent: Female|$45,000 to $49,999||Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Enrollment|F|Black||21|28269|Some College|Single|Business: Sales|28269|0|5|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|504038255|504040273|31|0|2|504034443|31|0|2|500814943|2||-2||4|1|500014681|500014681|-2|500014681|-2|34|2|||46|2|||1|855432|853694|4|3|45|8408514790530965815
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-26|NaT|Baseline|2015-02-24|2015-02-26|Complete|Done|3|3|4|3|3|3|3.17|||||||||4|4|3|4|4|3|3.67|||||||||4|4|3|3.67||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|||24.3||1|1|1|1|M|Black||14|No|Mother|28278|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|Black||29|28209|Bachelors Degree|Single|Finance|20877|0|8|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|504160892|504162947|31|0|1|504171934|31|0|1|500815454|2||-2||2|1|||-2||-2|0|4|||130|1|||1|854521|-1|4|3|44|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-26|NaT|Followup|2016-02-26|2016-05-12|Expired|Late||||||||3|3|4|3|3|3|3.17|||||||||4|4|3|4|4|3|3.67||||||4|4|3|3.67|||||||4|4|5|5|4.5||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|2|2.5||||1|1||||4|4||Green|||24.3||1|1|1|1|M|Black||14|No|Mother|28278|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|Black||29|28209|Bachelors Degree|Single|Finance|20877|0|8|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|504160892|504162947|31|0|1|504171934|31|0|1|500815454|2||-2||2|1|||-2||-2|0|4|||130|1|||1|855224|854521|4|0|45|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-02-27|2015-04-30|Baseline|2015-02-12|2015-02-27|Comprehension|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|PERL 2014-2016|Child: Severity of challenges|2||1|1|1|1|M|Black||11|No|Mother|28202|2|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||26|28205|Bachelors Degree|Single|Business: Sales|28205|1|1|BBBS National Site|Web Link|Big|General Community||RTBM|277|60|598|500000170|500008321|504003061|504005076|31|0|1|504169596|1|0|1|500813623|2||-2||4|3|500014681|500014681|-2||-2|34|2|||46|2|||1|851135|-1|4|2|44|8861782924354204409
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-28|NaT|Followup|2016-02-28|2016-04-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||24.2||3|3|1|1|F|Black||10|Yes|Aunt|28227|3|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|White||69|28104||Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|502643841|502255582|31|0|2|504076732|1|0|2|500812797|2||-2||2|1||500000294|-2||-2|0|10|||46|2|||1|877278||4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-02|NaT|Baseline|2015-02-22|2015-03-02|Complete|Done|1|4|4|4|1|1|2.5|||||||||2|4|2|4|3|3|3|||||||||1|4|3|2.67||||||5|4|2|5|4|||||||4|4|4|4|3|4|4|3.86||||||||||4|3|2|3||||||3|2|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||24.2||1|1|1|1|F|Black||13|No|Mother|28216|6|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||33|28205|Bachelors Degree|Single|Tech: Sales, Mktg|28217|7|11|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|504038302|504040320|31|0|2|504099787|1|0|2|500815247|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|5|||7464|9|||1|853687|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-02|NaT|Baseline|2015-02-23|2015-03-02|Complete|Done|4|1|2|1|1|3|2|||||||||3|3|3|2|1|4|2.67|||||||||3|4|2|3||||||4|5|2|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Green|||24.2||1|1|1|1|M|Black||15|No|Mother|28105|7|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||45|28226|Bachelors Degree|Single|Insurance|28226|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|503413167|503415024|31|0|1|504190868|1|0|1|500815087|2||-2||2|1|||-2||-2|34|2|||17159|12|||1|853968|-1|4|3|44|3714886275549507192
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-02|NaT|Followup|2016-03-02|2016-05-17|Expired|Late||||||||1|4|4|4|1|1|2.5|||||||||2|4|2|4|3|3|3||||||1|4|3|2.67|||||||5|4|2|5|4||||||||||4|4|4|4|3|4|4|3.86||||||4|3|2|3|||||3|2|2.5||||2|2||||4|4||Green|PERL 2014-2016||24.2||1|1|1|1|F|Black||13|No|Mother|28216|6|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||33|28205|Bachelors Degree|Single|Tech: Sales, Mktg|28217|7|11|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|504038302|504040320|31|0|2|504099787|1|0|2|500815247|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|5|||7464|9|||1|856652|853687|4|0|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-02|NaT|Followup|2016-03-02|2016-05-17|Expired|Late||||||||4|1|2|1|1|3|2|||||||||3|3|3|2|1|4|2.67||||||3|4|2|3|||||||4|5|2|3|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|4|4||||1|1||||4|4||Green|||24.2||1|1|1|1|M|Black||15|No|Mother|28105|7|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||45|28226|Bachelors Degree|Single|Insurance|28226|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|503413167|503415024|31|0|1|504190868|1|0|1|500815087|2||-2||2|1|||-2||-2|34|2|||17159|12|||1|856713|853968|4|0|45|3714886275549507192
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-09|2016-01-27|Baseline|2015-02-13|2015-03-09|Complete|Done|4|2|1|1|1|3|2|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|1|3||||||4|4|4|||||2|2||||4|4||||Red|PERL 2014-2016|Child/Family: Moved|10.6||1|1|1|1|M|Black||12|No|Mother|29301|5|Two Parent|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28203|Bachelors Degree|Single|Business|28208|0|1|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504152161|504154211|31|0|1|504180963|1|0|1|500813750|2||-2||4|3|500014681|500014681|-2|500014681|-2|0|4|||46|2|||1|851374|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-09|2016-03-23|Baseline|2015-03-05|2015-03-09|Complete|Done|3|4|4|4|2|3|3.33|||||||||2|3|4|4|4|4|3.5|||||||||4|4|3|3.67||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Time constraint|12.5||1|1|1|1|F|Black||15|No|Mother|28208|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||28|28204|Bachelors Degree|Single|Finance: Accountant|28277|0|3|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500018851|504075196|504048929|31|0|2|504108003|1|0|2|500817229|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|4|||46|2|||1|857926|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-12|NaT|Baseline|2015-03-03|2015-03-12|Complete|Done|4|3|1|3|4|4|3.17|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||23.9||1|1|1|1|M|Black||11|No|Mother|28215|3|One Parent: Female|$30,000 to $34,999||Yes||School|General Community||Match Support|M|Black||44|28173|Masters Degree|Married|Tech: Computer/Programmer|28202|7|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020910|503794892|503796869|31|0|1|504175530|31|0|1|500816649|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|857020|-1|4|3|44|3643651798871536206
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-12|NaT|Followup|2016-03-12|2016-05-27|Expired|Late||||||||4|3|1|3|4|4|3.17|||||||||2|4|4|2|3|4|3.17||||||4|4|4|4|||||||3|5|5|5|4.5||||||||||4|4|4|4|4|4|2|3.71||||||4|4|4|4|||||2|4|3||||2|2||||4|4||Green|||23.9||1|1|1|1|M|Black||11|No|Mother|28215|3|One Parent: Female|$30,000 to $34,999||Yes||School|General Community||Match Support|M|Black||44|28173|Masters Degree|Married|Tech: Computer/Programmer|28202|7|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020910|503794892|503796869|31|0|1|504175530|31|0|1|500816649|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|859786|857020|4|0|45|3643651798871536206
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-16|2016-08-02|Baseline|2015-02-24|2015-03-16|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|3|3|4|3.71||||||||||3|4|4|3.67||||||1|3|2|||||2|2||||4|4||||Green||Volunteer: Moved|16.6||1|1|1|1|F|Black||14|No|Mother|28213|6|One Parent: Female|$40,000 to $44,999||Yes|BBBS National Site|Web Link|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|F|Black||23|28262|Some College|Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504038196|504040273|31|0|2|504062905|31|0|2|500815275|2||-2||4|1||500007920, 500011315, 500011316|-2||-2|34|2|||17159|12|||1|854296|-1|4|3|44|8408514790530965815
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-16|2016-03-23|Baseline|2015-03-05|2015-03-16|Complete|Done|2|1|4|1|1|4|2.17|||||||||4|1|4|4|1|3|2.83|||||||||3|4|4|3.67||||||4|4|5|5|4.5|||||||4|4|4|4|3|4|2|3.57||||||||||4|3|4|3.67||||||2|2|2|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|12.3||1|1|1|1|M|Black||12|No|Mother|28211|4|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|Black||27|28215|High School Graduate|Single|Transport: Driver|28202|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503312337|503314167|31|0|1|504201470|31|0|1|500817147|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|857825|-1|4|3|44|4253272603994307857
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-16|2016-08-02|Followup|2016-03-16|2016-05-09|Complete|Late|3|4|4|4|4|4|3.83|4|4|4|3|4|4|3.83|0|3|4|4|4|2|4|3.5|4|4|4|4|4|4|4|-12.5|4|4|4|4|4|4|4|4|0|5|5|5|4|4.75|5|5|5|5|5|-5|4|4|4|4|4|4|3|3.86|4|4|4|4|3|3|4|3.71|4.04|3|3|4|3.33|3|4|4|3.67|-9.26|3|3|3|1|3|2|50|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|16.6||1|1|1|1|F|Black||14|No|Mother|28213|6|One Parent: Female|$40,000 to $44,999||Yes|BBBS National Site|Web Link|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|F|Black||23|28262|Some College|Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504038196|504040273|31|0|2|504062905|31|0|2|500815275|2||-2||4|1||500007920, 500011315, 500011316|-2||-2|34|2|||17159|12|||1|860623|854296|4|3|45|8408514790530965815
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-16|NaT|Followup|2016-03-16|2016-05-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||23.7||1|1|1|1|M|Black||10|No|Mother|28211|2|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||31|28209|Bachelors Degree|Married|Medical|70112|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|503314773|503314167|31|0|1|504176084|1|0|1|500817494|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|979708||4|1|45|4253272603994307857
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-17|2016-08-30|Followup|2016-03-17|2016-03-17|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|4|3|2|4|4|3.17|||||||||4|3|4|3.67||||||3|5|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Moved|17.5||2|2|1|1|M|Black||15||GrandMother|28227|3|One Parent: Female|Unknown|Y|Yes|AARTF|BBBS Board/Staff|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||25|28202|Bachelors Degree|Single|Finance: Banking|28202|0|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500018851|502287066|502287498|31|0|1|504056150|1|0|1|500814738|2||-2||4|1|500014681|500005291|-2|500014681|-2|7294|13|||17159|12|||1|861093||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-17|NaT|Baseline|2015-03-16|2015-03-17|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|3|4|1|2|4|2.67|||||||||4|4|4|4||||||5|1|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||1|1||||4|4||||Green|PERL 2014-2016||23.7||1|1|1|1|M|Black||12|No|Aunt|28216|7|One Parent: Female|$40,000 to $44,999||Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||33|28208|Masters Degree|Married|Finance|28202|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503946469|503948477|31|0|1|504188283|31|0|1|500818848|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|860764|-1|4|3|44|529594392811859839
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-17|NaT|Followup|2016-03-17|2016-03-15|Complete|Done|1|4|4|4|4|4|3.5|4|4|4|1|4|4|3.5|0|2|4|4|1|4|4|3.17|2|3|4|1|2|4|2.67|18.73|4|4|4|4|4|4|4|4|0|3|5|4|3|3.75|5|1|3|4|3.25|15.38|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|2|3|2.5|2|4|3|-16.67|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||23.7||1|1|1|1|M|Black||12|No|Aunt|28216|7|One Parent: Female|$40,000 to $44,999||Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||33|28208|Masters Degree|Married|Finance|28202|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503946469|503948477|31|0|1|504188283|31|0|1|500818848|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|861046|860764|4|3|45|529594392811859839
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-25|2016-09-29|Baseline|2015-03-23|2015-03-25|Complete|Done|3|4|4|4|3|3|3.5|||||||||4|2|4|4|4|4|3.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|2|3||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|18.2||1|1|1|1|M|White||16|No|Mother|28078|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance|28412|1|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500021785|504104035|504106070|1|0|1|504214658|1|0|1|500820084|2||-2||4|1|||-2||-2|0|5|||17159|12|||1|862933|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-25|2016-09-29|Followup|2016-03-25|2016-06-09|Expired|Late||||||||3|4|4|4|3|3|3.5|||||||||4|2|4|4|4|4|3.67||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|4|4|4|4|4||||||3|4|2|3|||||3|3|3||||2|2||||4|4||Green||Volunteer: Lost contact with child/agency|18.2||1|1|1|1|M|White||16|No|Mother|28078|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance|28412|1|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500021785|504104035|504106070|1|0|1|504214658|1|0|1|500820084|2||-2||4|1|||-2||-2|0|5|||17159|12|||1|863773|862933|4|0|45|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-26|2016-02-22|Baseline|2015-03-26|2015-03-26|Complete|Done|3|4|2|2|3|3|2.83|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||2|3|3|4|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Lost contact with child/agency|10.9||1|1|1|1|M|Black||13|No|Mother|28215|5|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||26|28204|Bachelors Degree|Single|Consultant|28244|1|6|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500018851|502722096|502722991|31|0|1|504213418|1|0|1|500820735|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|10|||17159|12|||1|864221|-1|4|3|44|8136849793711030748
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-26|2017-02-28|Baseline|2015-03-26|2015-03-26|Complete|Done|3|2|4|1|3|3|2.67|||||||||2|3|2|3|2|2|2.33|||||||||3|4|4|3.67||||||1|3|5|5|3.5|||||||4|4|4|4|4|3|3|3.71||||||||||2|4|3|3||||||1|3|2|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Moved|23.2||1|1|1|1|M|Black||14|No|Mother|28262|7|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||32|28262|Bachelors Degree|Single|Customer Service|28262|2|6|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|504045474|504047495|31|0|1|504228594|31|0|1|500820783|2||-2||4|3|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|864349|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-26|2017-02-28|Followup|2016-03-26|2016-04-22|Complete|Done|3|2|2|2|2|3|2.33|3|2|4|1|3|3|2.67|-12.73|2|3|3|2|3|3|2.67|2|3|2|3|2|2|2.33|14.59|3|2|2|2.33|3|4|4|3.67|-36.51|2|2|2|3|2.25|1|3|5|5|3.5|-35.71|4|4|4|4|4|4|3|3.86|4|4|4|4|4|3|3|3.71|4.04|3|3|3|3|2|4|3|3|0|2|3|2.5|1|3|2|25|2|2|2|2|0|4|4|4|4|0|Red|PERL 2014-2016|Volunteer: Moved|23.2||1|1|1|1|M|Black||14|No|Mother|28262|7|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||32|28262|Bachelors Degree|Single|Customer Service|28262|2|6|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|504045474|504047495|31|0|1|504228594|31|0|1|500820783|2||-2||4|3|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|864351|864349|4|3|45|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-26|NaT|Baseline|2015-03-10|2015-03-26|Complete|Done|2|1|2|1|3|4|2.17|||||||||1|4|2|2|3|4|2.67|||||||||2|3|3|2.67||||||4|5|4|5|4.5|||||||3|2|4|4|4|2|2|3||||||||||4|4|3|3.67||||||1|2|1.5|||||1|1||||4|4||||Yellow|||23.4||1|1|1|1|F|Black||11|No|Mother|28227|3|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||29|28226|Bachelors Degree|Single|Finance: Accountant|28202|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|504194601|504184323|31|0|2|504032490|1|0|2|500817776|2||-2||2|2|||-2||-2|0|4|||7464|9|||1|859018|-1|4|3|44|5822555200185981373
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-26|NaT|Followup|2016-03-26|2016-04-22|Complete|Done|4|2|3|2|3|4|3|2|1|2|1|3|4|2.17|38.25|3|3|3|3|4|3|3.17|1|4|2|2|3|4|2.67|18.73|4|4|4|4|2|3|3|2.67|49.81|3|3|3|3|3|4|5|4|5|4.5|-33.33|4|4|4|4|4|4|4|4|3|2|4|4|4|2|2|3|33.33|4|4|4|4|4|4|3|3.67|8.99|3|3|3|1|2|1.5|100|2|2|1|1|100|4|4|4|4|0|Yellow|||23.4||1|1|1|1|F|Black||11|No|Mother|28227|3|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||29|28226|Bachelors Degree|Single|Finance: Accountant|28202|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|504194601|504184323|31|0|2|504032490|1|0|2|500817776|2||-2||2|2|||-2||-2|0|4|||7464|9|||1|864248|859018|4|3|45|5822555200185981373
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-30|2017-02-27|Followup|2016-03-30|2016-05-16|Complete|Late|3|3|3|3|3|4|3.17|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|23||1|1|1|1|F|Black||10|Yes|Mother|28273|2|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Black||29|28269||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|504165894|504167953|31|0|2|504138163|31|0|2|500821104|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|952690||4|3|45|5161383151676749743
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-30|NaT|Followup|2016-03-30|2016-03-24|Complete|Done|4|3|3|1|4|4|3.17|||||||||1|4|2|1|1|2|1.83|||||||||4|4|4|4||||||2|2|2|2|2|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|||23.3||2|2|2|2|M|Black||10|Yes|Mother|28216|1|One Parent: Female|Less than $10,000||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||42|28205|Bachelors Degree|Married|Arts, Entertainment, Sports|28205|14|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020910|503565647|503567522|31|0|1|503865770|1|0|1|500819520|2||-2||2|1||500000294|-2|500000294|-2|34|2|||17159|12|||1|988940||4|3|45|1786514887916898235
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-31|2017-02-27|Baseline|2015-03-31|2015-03-31|Complete|Done|3|1|3|1|3|4|2.5|||||||||2|1|4|2|2|4|2.5|||||||||4|4|4|4||||||2|4|5|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|23||1|1|1|1|F|Black||13|No|Mother|28273|5|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Black||28|28105|Masters Degree|Single|Business: Human Resources|28078|0|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|504165911|504167953|31|0|2|504030347|31|0|2|500821362|2||-2||4|1|||-2||-2|0|4|||46|2|||1|865805|-1|4|3|44|5161383151676749743
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-31|2017-02-27|Followup|2016-03-31|2016-05-16|Complete|Late|3|3|3|3|3|3|3|3|1|3|1|3|4|2.5|20|3|4|4|3|3|4|3.5|2|1|4|2|2|4|2.5|40|4|4|4|4|4|4|4|4|0|4|4|4|4|4|2|4|5|4|3.75|6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Time constraint|23||1|1|1|1|F|Black||13|No|Mother|28273|5|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Black||28|28105|Masters Degree|Single|Business: Human Resources|28078|0|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|504165911|504167953|31|0|2|504030347|31|0|2|500821362|2||-2||4|1|||-2||-2|0|4|||46|2|||1|865829|865805|4|3|45|5161383151676749743
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-03-31|2016-08-29|Followup|2016-03-31|2016-06-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|VOL - Mentoring Hispanic Youth|Child: Family structure changed|17||1|1|1|1|M|Hispanic||10|No|Mother|28214|2|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|VOL - Mentoring Hispanic Youth|Match Support|M|Hispanic||40|28277|Bachelors Degree|Married|Insurance|28277|8|0|Current/Previous Big|Other Big|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|277|60|598|500000170|500017777|504059287|504061304|3|0|1|504210666|3|0|1|500819684|2||-2||4|3|500011312|500011312|-2|500011312|-2|0|5|||17159|12|||1|955440||4|0|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-31|NaT|Baseline|2015-03-14|2015-03-31|Complete|Done|1|4|4|3|4|4|3.33|||||||||2|4|3|3|2|2|2.67|||||||||4|4|4|4||||||2|4|3|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||3|3|2|2.67||||||3|2|2.5|||||2|2||||4|4||||Green|||23.2||1|1|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Business: Sales|28277|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|501843066|501843435|31|0|2|504152982|1|0|2|500818696|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|860440|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-31|NaT|Followup|2016-03-31|2016-04-22|Complete|Done|2|3|4|3|4|4|3.33|1|4|4|3|4|4|3.33|0|3|4|3|3|3|3|3.17|2|4|3|3|2|2|2.67|18.73|4|4|4|4|4|4|4|4|0|3|3|3|3|3|2|4|3|3|3|0|4|4|4|4|3|4|4|3.86|4|4|4|4|3|4|3|3.71|4.04|2|3|3|2.67|3|3|2|2.67|0|3|2|2.5|3|2|2.5|0|2|2|2|2|0|4|4|4|4|0|Green|||23.2||1|1|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Business: Sales|28277|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|501843066|501843435|31|0|2|504152982|1|0|2|500818696|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|866058|860440|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-13|2016-10-31|Baseline|2015-04-13|2015-04-13|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|18.6||1|1|1|1|M|Black||10|No|Mother|28212|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Business|33701|2|11|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504122670|504124721|31|0|1|504179830|1|0|1|500817495|2||-2||4|3|||-2||-2|0|4|||46|2|||1|869333|-1|4|1|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-13|2016-10-31|Followup|2016-04-13|2016-05-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|18.6||1|1|1|1|M|Black||10|No|Mother|28212|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Business|33701|2|11|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504122670|504124721|31|0|1|504179830|1|0|1|500817495|2||-2||4|3|||-2||-2|0|4|||46|2|||1|869334|869333|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-04-13|NaT|Baseline|2015-04-13|2015-04-13|Complete|Done|4|2|4|2|3|4|3.17|||||||||2|4|3|4|2|4|3.17|||||||||4|4|4|4||||||4|3|2|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||22.8||1|1|1|1|M|Black||13|No|Mother|28208|6|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||25|28203|Masters Degree|Single|Finance: Accountant|28202|0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504068125|504070152|31|0|1|504241807|1|0|1|500822990|2||-2||2|1|||-2||-2|0|10|||46|2|||1|869371|-1|4|3|44|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-04-13|NaT|Followup|2016-04-13|2016-04-22|Complete|Done|4|4|4|2|4|4|3.67|4|2|4|2|3|4|3.17|15.77|3|3|4|3|3|3|3.17|2|4|3|4|2|4|3.17|0|4|4|4|4|4|4|4|4|0|4|2|3|5|3.5|4|3|2|4|3.25|7.69|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|4|4|4|4|-8.25|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green|||22.8||1|1|1|1|M|Black||13|No|Mother|28208|6|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||25|28203|Masters Degree|Single|Finance: Accountant|28202|0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504068125|504070152|31|0|1|504241807|1|0|1|500822990|2||-2||2|1|||-2||-2|0|10|||46|2|||1|869384|869371|4|3|45|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-14|2015-10-07|Baseline|2015-03-26|2015-04-14|Complete|Done|2|1|3|1|2|3|2|||||||||2|4|2|2|3|2|2.5|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Moved|5.8||1|2|1|1|F|Multi-race (Hispanic & White)||13|No|Mother|28205|7|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community||Pending Match|F|White||30|28205|Bachelors Degree|Separated|Business|28205|0|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504205508|504207619|35|0|2|504157187|1|0|2|500820606|2||-2||4|3|500014681||-2|500014681|-2|0|5|||17159|12|||1|863991|-1|4|3|44|610388910998118020
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-04-14|NaT|Baseline|2015-04-13|2015-04-14|Complete|Done|3|1|1|3|2|1|1.83|||||||||2|3|2|1|2|2|2|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||3|2|2|2.33||||||4|4|4|||||2|2||||4|4||||Green|||22.8||1|1|1|1|F|Black||13|No|Mother|28205|5|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|Black||27|28262|Some College|Single|Medical: Healthcare Worker|28210|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504242976|504245092|31|0|2|504198992|31|0|2|500823043|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|869474|-1|4|3|44|3988279022378749151
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-04-14|NaT|Followup|2016-04-14|2016-04-22|Complete|Done|1|4|3|2|2|2|2.33|3|1|1|3|2|1|1.83|27.32|2|3|2|2|2|3|2.33|2|3|2|1|2|2|2|16.5|4|4|4|4|4|4|4|4|0|3|3|3|3|3|4|5|3|4|4|-25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|3|3|3.71|4.04|2|3|2|2.33|3|2|2|2.33|0|2|3|2.5|4|4|4|-37.5|2|2|2|2|0|4|4|4|4|0|Green|||22.8||1|1|1|1|F|Black||13|No|Mother|28205|5|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|Black||27|28262|Some College|Single|Medical: Healthcare Worker|28210|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504242976|504245092|31|0|2|504198992|31|0|2|500823043|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|869872|869474|4|3|45|3988279022378749151
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-16|2016-09-16|Baseline|2015-03-18|2015-04-16|Complete|Done|3|1|4|3|2|3|2.67|||||||||2|4|4|1|3|3|2.83|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|3|2|3.57||||||||||3|4|2|3||||||2|3|2.5|||||1|1||||4|4||||Green||Child: Lost interest|17.1||1|1|1|1|F|Black||11|No|Father|28205|4|One Parent: Male|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Black||56|28216|High School Graduate|Married|Unemployed||0|0|United Way|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500018851|504221885|504223999|31|0|2|504188499|31|0|2|500819243|2||-2||4|1|||-2||-2|0|4|||16263|6|||1|861392|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-16|2016-09-16|Followup|2016-04-16|2016-07-01|Expired|Late||||||||3|1|4|3|2|3|2.67|||||||||2|4|4|1|3|3|2.83||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|4|4|3|2|3.57||||||3|4|2|3|||||2|3|2.5||||1|1||||4|4||Green||Child: Lost interest|17.1||1|1|1|1|F|Black||11|No|Father|28205|4|One Parent: Male|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Black||56|28216|High School Graduate|Married|Unemployed||0|0|United Way|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500018851|504221885|504223999|31|0|2|504188499|31|0|2|500819243|2||-2||4|1|||-2||-2|0|4|||16263|6|||1|870525|861392|4|0|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-20|2016-08-01|Baseline|2015-04-07|2015-04-20|Complete|Done|3|4|4|4|4|3|3.67|||||||||1|4|4|1|1|1|2|||||||||4|3|2|3||||||5|4|3|4|4|||||||4|4|4|4|3|3|3|3.57||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Lost contact with child/agency|15.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$15,000 to $19,999||Yes||Relative|General Community|PERL 2014-2016|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Engineer||0|2|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503679979|503226552|31|0|1|504191848|1|0|1|500822162|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|3|||7464|9|||1|867614|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-20|2016-08-01|Followup|2016-04-20|2016-06-15|Declined|Late||||||||3|4|4|4|4|3|3.67|||||||||1|4|4|1|1|1|2||||||4|3|2|3|||||||5|4|3|4|4||||||||||4|4|4|4|3|3|3|3.57||||||4|4|3|3.67|||||4|3|3.5||||2|2||||4|4||Green|PERL 2014-2016|Volunteer: Lost contact with child/agency|15.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$15,000 to $19,999||Yes||Relative|General Community|PERL 2014-2016|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Engineer||0|2|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503679979|503226552|31|0|1|504191848|1|0|1|500822162|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|3|||7464|9|||1|871528|867614|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-21|2015-12-02|Baseline|2015-04-11|2015-04-21|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|3|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Feels incompatible with child/family|7.4||1|1|2|2|M|Black||14|No|Mother|28213|7|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community|PERL 2014-2016|RTBM|M|White||32|28202|Masters Degree|Single|Finance: Accountant|28202|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|503917561|503962680|31|0|1|504206321|1|0|1|500822824|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|868959|-1|4|3|44|6084148439133243542
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-27|2016-09-16|Baseline|2015-03-24|2015-04-27|Complete|Done|2|4|4|3|3|3|3.17|||||||||3|2|3|3|4|3|3|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|4|3|||||1|1||||4|4||||Green||Volunteer: Time constraint|16.7||1|1|1|1|F|Black||13|Yes|Mother|28208|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|F|White||33|28202|Bachelors Degree|Divorced|Business|28117|4|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018851|504075185|504048929|31|0|2|504169746|1|0|2|500822245|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|863157|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-27|2015-10-09|Baseline|2015-04-16|2015-04-27|Complete|Done|3|3|4|3|3|2|3|||||||||2|1|2|3|3|3|2.33|||||||||2|2|2|2||||||2|2|4|5|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|2|2.5|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Feels incompatible with child/family|5.4||2|2|2|2|F|Black||15|No|Mother|28262|8|One Parent: Female|$45,000 to $49,999||No||School|General Community|PERL 2014-2016|Match Support|F|Black||38|28269|Masters Degree|Single|Business|28262|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|277|60|598|500000170|500017777|503974135|503598965|31|0|2|503860995|31|0|2|500823546|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|870595|-1|4|3|44|1198499568025045356
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-27|2016-09-16|Followup|2016-04-27|2016-07-12|Expired|Late||||||||2|4|4|3|3|3|3.17|||||||||3|2|3|3|4|3|3||||||4|4|4|4|||||||3|4|4|5|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||2|4|3||||1|1||||4|4||Green||Volunteer: Time constraint|16.7||1|1|1|1|F|Black||13|Yes|Mother|28208|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|F|White||33|28202|Bachelors Degree|Divorced|Business|28117|4|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018851|504075185|504048929|31|0|2|504169746|1|0|2|500822245|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|874050|863157|4|0|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-28|2016-08-29|Baseline|2015-04-11|2015-04-28|Complete|Done|3|2|3|3|3|4|3|||||||||2|2|3|3|1|3|2.33|||||||||4|4|4|4||||||5|3|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|4|3|||||1|1||||4|4||||Red|VOL - Mentoring Hispanic Youth, PERL 2014-2016|Volunteer: Moved|16.1||1|1|1|1|M|Hispanic||14|No|Mother|28215|8|One Parent: Female|Unknown|Y|Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Enrollment|M|Hispanic||27|28262|Some College|Single|Finance: Banking|28228|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|277|60|598|500000170|500017777|504154297|504156341|3|0|1|504201847|3|0|1|500822827|2||-2||4|3|500011312, 500014681|500011312, 500014681|-2|500011312, 500014681|-2|0|10|||17159|12|||1|868966|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-28|2016-08-29|Followup|2016-04-28|2016-07-13|Expired|Late||||||||3|2|3|3|3|4|3|||||||||2|2|3|3|1|3|2.33||||||4|4|4|4|||||||5|3|4|4|4||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||2|4|3||||1|1||||4|4||Red|VOL - Mentoring Hispanic Youth, PERL 2014-2016|Volunteer: Moved|16.1||1|1|1|1|M|Hispanic||14|No|Mother|28215|8|One Parent: Female|Unknown|Y|Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Enrollment|M|Hispanic||27|28262|Some College|Single|Finance: Banking|28228|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|277|60|598|500000170|500017777|504154297|504156341|3|0|1|504201847|3|0|1|500822827|2||-2||4|3|500011312, 500014681|500011312, 500014681|-2|500011312, 500014681|-2|0|10|||17159|12|||1|874742|868966|4|0|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-29|2016-03-21|Baseline|2015-04-29|2015-04-29|Complete|Done|2|3|3|2|4|3|2.83|||||||||2|2|3|2|2|3|2.33|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|2|2|||||1|1||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|10.7||1|1|1|1|F|Black||11|No|Mother|28212|3|One Parent: Female|$25,000 to $29,999||Yes||School|General Community||Match Support|F|White||26|28205||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500017732|504231007|504233122|31|0|2|504163497|1|0|2|500825416|2||-2||4|1|||-2||-2|0|4|||17159|12|||1|875638|-1|4|3|44|8136849793711030748
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-04-30|2015-06-25|Baseline|2015-04-23|2015-04-30|Complete|Done|1|1|1|4|4|4|2.5|||||||||2|2|3|3|3|4|2.83|||||||||4|4|4|4||||||5|5|5|3|4.5|||||||4|4|4|4|4|4|4|4||||||||||1|4|1|2||||||4|1|2.5|||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|1.8||2|2|1|1|F|Black||11|No|Mother|28269|5|One Parent: Female|$50,000 to $59,999|Y|No||School|General Community||Match Support|F|White||27|28202|Some College|Single|Transport: Flight Attendant||2|1|Local TV|Media|Big|General Community||Enrollment|277|60|598|500000170|500017732|504243465|504245581|31|0|2|504173742|1|0|2|500824646|2||-2||4|1|||-2||-2|0|4|||7438|1|||1|873076|-1|4|3|44|2806833304218536184
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-04-30|NaT|Followup|2016-04-30|2016-06-15|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|PERL 2014-2016||22.2||1|1|2|2|M|Multi-race (Black & Hispanic)||10|Yes|GrandMother|28208|1|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community|Amachi, PERL 2014-2016|Match Support|M|Asian||33|28204|Bachelors Degree|Married|Business: Engineer|28007|3|9|Man Up Campaign|Media|Big|General Community|Amachi, PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503433219|503227914|38|0|1|503890372|4|0|1|500822826|2||-2||2|1|500014681|500000294, 500014681|-2|500000294, 500014681|-2|0|10|||17101|1|||1|958046||4|1|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-04|2016-05-19|Baseline|2015-05-03|2015-05-04|Complete|Done|3|4|1|2|4|3|2.83|||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||1|1||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|12.5||2|2|1|1|M|Black||10|Yes|Mother|28213|3|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community|Amachi|Match Support|M|White||31|28105|Bachelors Degree|Married|Consultant|43215|1|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504240016|504242131|31|0|1|504155486|1|0|1|500825676|2||-2||4|1||500000294|-2||-2|0|10|||17159|12|||1|876717|-1|4|3|44|3326174373441625173
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-04|2015-10-07|Baseline|2015-05-04|2015-05-04|Complete|Done|3|1|3|2|3|3|2.5|||||||||2|4|4|2|2|3|2.83|||||||||4|4|3|3.67||||||5|3|2|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Red||Child/Family: Moved|5.1||1|1|1|1|M|Black||14|Yes|Mother|28216|5|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Enrollment|M|Black||37|28213|Some College|Living w/ Significant Other|Self-Employed, Entrepreneur|28206|2|0|Current/Previous Big|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500013781|502821218|502822501|31|0|1|504244628|31|0|1|500825744|2||-2||4|3|||-2||-2|0|10|||17159|12|||1|877039|-1|4|3|44|6971797047831566199
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Baseline|2015-04-22|2015-05-04|Complete|Done|2|1|1|1|1|1|1.17|||||||||2|2|2|1|3|2|2|||||||||4|4|4|4||||||2|2|5|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||22.1||1|1|1|1|M|White||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999||Yes||School|General Community||Match Support|M|White||51|28173|Masters Degree|Married|Self-Employed, Entrepreneur|28173|19|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504235369|504237484|1|0|1|503937954|1|0|1|500824366|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|872406|-1|4|3|44|8961132295198487522
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Baseline|2015-04-24|2015-05-04|Complete|Done|4|2|3|3|3|4|3.17|||||||||2|3|3|3|2|3|2.67|||||||||4|3|3|3.33||||||4|3|2|2|2.75|||||||2|4|4|4|4|4|4|3.71||||||||||4|4|3|3.67||||||2|4|3|||||1|1||||4|4||||Green|||22.1||1|1|1|1|F|White||15|No|Mother|28227|8|One Parent: Female|$35,000 to $39,999||Yes||School|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Law: Paralegal|28211|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504235352|504237484|1|0|2|504200139|1|0|2|500825073|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|873520|-1|4|3|44|8961132295198487522
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Followup|2016-05-05|2016-05-09|Complete|Done|3|2|1|1|2|3|2|2|1|1|1|1|1|1.17|70.94|2|3|4|2|1|3|2.5|2|2|2|1|3|2|2|25|4|4|4|4|4|4|4|4|0|3|3|3|3|3|2|2|5|5|3.5|-14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|4|3.67|4|4|4|4|-8.25|3|4|3.5|4|4|4|-12.5|2|2|2|2|0|4|4|4|4|0|Green|||22.1||1|1|1|1|M|White||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999||Yes||School|General Community||Match Support|M|White||51|28173|Masters Degree|Married|Self-Employed, Entrepreneur|28173|19|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504235369|504237484|1|0|1|503937954|1|0|1|500824366|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|877351|872406|4|3|45|8961132295198487522
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Followup|2016-05-05|2016-05-09|Complete|Done|3|3|3|3|4|4|3.33|4|2|3|3|3|4|3.17|5.05|2|2|3|2|1|4|2.33|2|3|3|3|2|3|2.67|-12.73|3|3|2|2.67|4|3|3|3.33|-19.82|2|4|4|4|3.5|4|3|2|2|2.75|27.27|3|4|3|1|4|3|3|3|2|4|4|4|4|4|4|3.71|-19.14|3|3|2|2.67|4|4|3|3.67|-27.25|4|4|4|2|4|3|33.33|1|1|1|1|0|4|4|4|4|0|Green|||22.1||1|1|1|1|F|White||15|No|Mother|28227|8|One Parent: Female|$35,000 to $39,999||Yes||School|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Law: Paralegal|28211|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504235352|504237484|1|0|2|504200139|1|0|2|500825073|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|877359|873520|4|3|45|8961132295198487522
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-12|NaT|Followup|2016-05-12|2016-05-19|Complete|Done|3|1|2|2|1|4|2.17|||||||||2|1|4|4|4|4|3.17|||||||||2|4|4|3.33||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||21.8||1|1|1|1|F|White||10|No|Mother|28277|4|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community||Match Support|F|White||29|29708|Bachelors Degree|Married|Medical|28105|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|503889301|503891297|1|0|2|504021478|1|0|2|500823483|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|912396||4|3|45|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-13|NaT|Followup|2016-05-13|2016-05-25|Complete|Done|4|3|4|4|3|4|3.67|||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||21.8||1|1|1|1|F|White||10|No|Mother|28214|4|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community||Match Support|F|White||28|28206|Bachelors Degree|Single|Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|504231269|504233379|1|0|2|503927707|1|0|2|500826291|2||-2||2|1|||-2||-2|0|3|||46|2|||1|954853||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-19|2016-05-12|Baseline|2015-01-09|2015-05-19|Complete|Done|3|2|4|1|4|4|3|||||||||2|2|2|2|2|1|1.83|||||||||4|4|4|4||||||2|2|2|2|2|||||||4|4|4|4|4|4|4|4||||||||||3|4|2|3||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016|Child/Family: Lost contact with volunteer/agency|11.8||1|1|1|1|M|Black||14|No|Mother|28227|6|One Parent: Female|$10,000 to $14,999||Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Black||33|28215|Associate Degree|Single|Business|28202|0|3|Self|Self|Big|General Community|PERL 2014-2016|Enrollment|277|60|598|500000170|500020990|503941174|503943182|31|0|1|503207130|31|0|1|500825477|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|5|||7464|9|||1|839933|-1|4|3|44|7312235294346727700
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-19|NaT|Baseline|2015-01-27|2015-05-19|Complete|Done|3|4|4|4|3|3|3.5|||||||||3|2|3|3|2|3|2.67|||||||||4|3|3|3.33||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Green|||21.6||1|1|1|1|F|Black||15|No|Mother|28214|9|Two Parent|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|Black||22|28223||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504023342|504060686|31|0|2|504173078|31|0|2|500826184|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|845197|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-19|NaT|Followup|2016-05-19|2016-06-30|Complete|Done|2|4|4|4|4|4|3.67|3|4|4|4|3|3|3.5|4.86|2|3|3|4|3|3|3|3|2|3|3|2|3|2.67|12.36|3|3|3|3|4|3|3|3.33|-9.91|3|5|3|3|3.5|3|4|4|4|3.75|-6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|3|4|4|3.67|0|2|2|2|4|4|4|-50|2|2|2|2|0|4|4|4|4|0|Green|||21.6||1|1|1|1|F|Black||15|No|Mother|28214|9|Two Parent|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|Black||22|28223||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504023342|504060686|31|0|2|504173078|31|0|2|500826184|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|884131|845197|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-19|NaT|Followup|2016-05-19|2016-05-18|Complete|Done|4|4|4|1|4|4|3.5|4|4|4|1|2|2|2.83|23.67|2|4|3|1|1|3|2.33|4|2|1|1|2|4|2.33|0|4|4|4|4|1|4|4|3|33.33|4|4|4|4|4|4|3|3|5|3.75|6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|3|3.67|8.99|2|3|2.5|3|4|3.5|-28.57|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||21.6||2|2|1|1|M|White||13||GrandMother|28210|4|One Parent: Female|Unknown|Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||29|28217|Some College|Single|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503469072|503470938|1|0|1|504202910|1|0|1|500826264|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|884655|615797|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-19|NaT|Followup|2016-05-19|2016-05-18|Complete|Done|4|4|2|4|4|4|3.67|||||||||1|1|4|2|2|4|2.33|||||||||4|3|3|3.33||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|3|2.5|||||1|1||||4|4||||Green|PERL 2014-2016||21.6||1|1|1|1|F|White||10|No|GrandMother|28210|3|Other Relative|Unknown||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||28|28205|Some College|Single|Transport: Driver|28277|8|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504234369|503470938|1|0|2|504116244|35|0|2|500825294|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|910429||4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-20|2016-09-26|Baseline|2015-05-20|2015-05-20|Complete|Done|2|1|2|1|2|2|1.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child/Family: Moved|16.3||1|1|1|1|M|Black||14|No|Mother|28269|6|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|White||53|28203|Masters Degree|Married|Business: Sales|17601|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503874068|503876064|31|0|1|504196201|1|0|1|500827631|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|885162|-1|4|3|44|3501831218874457455
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-20|2016-09-26|Followup|2016-05-20|2016-06-28|Complete|Done|2|2|3|2|3|2|2.33|2|1|2|1|2|2|1.67|39.52|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|5|5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Red||Child/Family: Moved|16.3||1|1|1|1|M|Black||14|No|Mother|28269|6|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|White||53|28203|Masters Degree|Married|Business: Sales|17601|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503874068|503876064|31|0|1|504196201|1|0|1|500827631|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|885179|885162|4|3|45|3501831218874457455
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-22|NaT|Baseline|2015-05-22|2015-05-22|Complete|Done|3|1|4|2|3|4|2.83|||||||||3|4|3|3|2|4|3.17|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||21.5||1|1|2|2|F|Black||13|No|Mother|28212|7|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500018851|502930499|502931919|31|0|2|502564910|31|0|2|500828045|2||-2||2|1|||-2||-2|0|10|||17161|11|||1|887615|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-22|NaT|Followup|2016-05-22|2016-08-06|Expired|Late||||||||3|1|4|2|3|4|2.83|||||||||3|4|3|3|2|4|3.17||||||4|4|4|4|||||||4|5|5|4|4.5||||||||||4|4|4|4|4|4|2|3.71||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Green|||21.5||1|1|2|2|F|Black||13|No|Mother|28212|7|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500018851|502930499|502931919|31|0|2|502564910|31|0|2|500828045|2||-2||2|1|||-2||-2|0|10|||17161|11|||1|887617|887615|4|0|45|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-27|2015-07-14|Baseline|2015-05-21|2015-05-26|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|1|1.5|||||1|1||||4|4||||Yellow|PERL 2014-2016|Volunteer: Time constraint|1.6||2|2|1|1|M|American Indian or Alaska Native||14|No|Mother|28269|7|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||53|28027||Married|Tech: Management|28117|7|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500012459|504150667|504152735|6|0|1|503845717|1|0|1|500827880|2||-2||4|2|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|886556|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-27|NaT|Baseline|2011-04-29|2015-05-27|Complete|Done|4|4|4|4|3|4|3.83|||||||||3|4|3|4|3|4|3.5|||||||||4|4|4|4||||||3|5|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow|Cabarrus County||21.4||1|1|1|1|F|Black||15|No|Mother|28027|9|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community|2010-2012 OJJDP JJI, Cabarrus County|Match Support|F|White||27|28262|Associate Degree|Single|Self-Employed, Entrepreneur|28217|3|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502501997|502502446|31|0|2|504227306|1|0|2|500825847|2||500016307||2|2|500016374|500005291, 500016374|-2|500016374|-2|0|10|||17159|12|||1|273262|-1|4|3|44|2581014289501540602
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-27|NaT|Followup|2016-05-27|2016-06-14|Complete|Done|2|2|4|2|3|4|2.83|4|4|4|4|3|4|3.83|-26.11|2|4|4|4|2|4|3.33|3|4|3|4|3|4|3.5|-4.86|4|4|4|4|4|4|4|4|0|3|5|4|5|4.25|3|5|4|3|3.75|13.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|4|4|4|4|-8.25|3|2|2.5|4|4|4|-37.5|2|2|1|1|100|4|4|4|4|0|Yellow|Cabarrus County||21.4||1|1|1|1|F|Black||15|No|Mother|28027|9|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community|2010-2012 OJJDP JJI, Cabarrus County|Match Support|F|White||27|28262|Associate Degree|Single|Self-Employed, Entrepreneur|28217|3|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502501997|502502446|31|0|2|504227306|1|0|2|500825847|2||500016307||2|2|500016374|500005291, 500016374|-2|500016374|-2|0|10|||17159|12|||1|890411|273262|4|3|45|2581014289501540602
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-28|NaT|Baseline|2015-04-11|2015-05-28|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|4|3.5|||||1|1||||4|4||||Green|PERL 2014-2016||21.3||1|1|1|1|M|Multi-race (Black & Hispanic)||13|No|Mother|28208|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||29|28208|Masters Degree|Single|Finance: Accountant|28210|3|6|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|503924157|503926164|38|0|1|504277947|1|0|1|500827570|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|868958|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-28|NaT|Baseline|2015-05-11|2015-05-27|Complete|Done|2|2|2|1|1|3|1.83|||||||||2|3|3|4|3|3|3|||||||||4|4|4|4||||||2|3|4|2|2.75|||||||4|4|4|3|4|4|3|3.71||||||||||4|4|3|3.67||||||3|1|2|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||21.3||1|1|1|1|M|Black||11|No|Mother|28027|4|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||31|28027|Juris Doctorate (JD)|Married|Law: Lawyer|28036|2|10|Igniting Breakfast|Special Event|Big|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|502426625|502502446|31|0|1|504274174|1|0|1|500826502|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500000294, 500014681, 500016374|-2|0|10|||17266|8|||1|880022|-1|4|3|44|2581014289501540602
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-28|NaT|Followup|2016-05-28|2016-06-20|Complete|Done|3|4|4|2|3|3|3.17|2|2|2|1|1|3|1.83|73.22|2|4|3|2|2|3|2.67|2|3|3|4|3|3|3|-11|4|4|4|4|4|4|4|4|0|3|4|4|4|3.75|2|3|4|2|2.75|36.36|4|4|4|4|4|4|3|3.86|4|4|4|3|4|4|3|3.71|4.04|4|4|4|4|4|4|3|3.67|8.99|3|3|3|3|1|2|50|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016, Cabarrus County||21.3||1|1|1|1|M|Black||11|No|Mother|28027|4|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||31|28027|Juris Doctorate (JD)|Married|Law: Lawyer|28036|2|10|Igniting Breakfast|Special Event|Big|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|502426625|502502446|31|0|1|504274174|1|0|1|500826502|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500000294, 500014681, 500016374|-2|0|10|||17266|8|||1|890472|880022|4|3|45|2581014289501540602
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-28|NaT|Followup|2016-05-28|2016-06-29|Complete|Done|4|3|4|2|4|4|3.5|4|4|4|1|4|4|3.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|4|4|4|4.25|5|4|5|5|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3.67|8.99|3|3|3|3|4|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||21.3||1|1|1|1|M|Multi-race (Black & Hispanic)||13|No|Mother|28208|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||29|28208|Masters Degree|Single|Finance: Accountant|28210|3|6|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|503924157|503926164|38|0|1|504277947|1|0|1|500827570|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|891538|868958|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-29|2016-06-23|Baseline|2015-05-29|2015-05-29|Complete|Done|1|1|2|1|1|2|1.33|||||||||2|3|3|2|2|4|2.67|||||||||4|3|3|3.33||||||2|5|4|4|3.75|||||||4|4|4|4|4|4||||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016|Child/Family: Lost contact with volunteer/agency|12.8||1|1|1|1|F|Black||15|No|Mother|28227|8|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||22|28262||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504081466|504083495|31|0|2|504098772|1|0|2|500828761|2||-2||4|1|500014681|500014681|-2||-2|34|2|||17159|12|||1|892473|-1|4|3|44|4786128411006480901
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-05-31|2016-03-14|Baseline|2015-05-14|2015-05-31|Complete|Done|4|2|4|1|3|4|3|||||||||2|4|4|3|1|4|3|||||||||3|2|4|3||||||2|3|1|5|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|PERL 2014-2016|Child/Family: Moved|9.5||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28134|4|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28273|Bachelors Degree|Single|Architect|28273|0|11|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|504202968|504205079|36|0|1|504285700|1|0|1|500827095|2||-2||4|2|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|881906|-1|4|3|44|7165641474360673060
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-02|2016-04-27|Baseline|2015-05-05|2015-06-02|Complete|Done|3|2|4|1|4|4|3|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||3|4|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|10.8||1|1|1|1|M|Black||15|No|Mother|28273|8|One Parent: Female|$35,000 to $39,999||No|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||30|28208|Bachelors Degree|Single|Self-Employed, Entrepreneur|28078|2|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504159888|504161941|31|0|1|504240720|1|0|1|500825834|2||-2||4|3|500014681|500014681|-2|500014681|-2|34|2|||17159|12|||1|877407|-1|4|3|44|8491998754880714879
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-02|NaT|Followup|2016-06-02|2016-06-14|Complete|Done|2|3|4|3|2|2|2.67|3|3|2|3|2|3|2.67|0|3|3|3|3|3|3|3|3|2|3|2|2|3|2.5|20|4|4|4|4|4|3|4|3.67|8.99|4|4|4|4|4|3|3|3|1|2.5|60|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|3|4|2|3|22.33|2|2|2|4|4|4|-50|2|2|2|2|0|4|4|4|4|0|Green|mentor2.0, mentor2.0 2014||21.2||1|2|1|2|F|Hispanic||18|No|Mother|28217|9|One Parent: Female|Unknown|Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|F|Some Other Race||34|28216|Masters Degree|Living w/ Significant Other|Finance|28202|0|0|Local Print|Media|Big|General Community|mentor2.0 2014|Match Support|277|60|598|500000170|500022907|504043329|504045347|3|0|2|503918707|41|0|2|500828965|2||500015511||2|1|500014505, 500014506|500014505, 500014506|-2|500014506|-2|0|4|||7439|1|||1|897421|800009|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-03|NaT|Followup|2016-06-03|2016-06-14|Complete|Done|3|1|3|3|3|3|2.67|3|1|2|1|2|2|1.83|45.9|2|4|3|2|2|3|2.67|2|4|3|2|3|3|2.83|-5.65|4|3|3|3.33|4|4|3|3.67|-9.26|3|3|4|5|3.75|5|2|5|4|4|-6.25|4|4|4|4|3|3|3|3.57|4|4|4|3|1|4|3|3.29|8.51|3|3|2|2.67|2|3|4|3|-11|4|3|3.5|3|4|3.5|0|2|2|2|2|0|4|4|4|4|0|Green|mentor2.0, mentor2.0 2014||21.1||1|2|1|2|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown|Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|M|White||60|28211|Masters Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|277|60|598|500000170|500022907|504043397|504045415|31|0|1|503922094|1|0|1|500828963|2||500015511||2|1|500014505, 500014506|500014505, 500014506|-2|500014506|-2|0|4|||7671|13|||1|898565|800115|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-04|2017-02-06|Followup|2016-06-04|2016-07-30|Complete|Late|3|2|3|4|2|3|2.83|||||||||4|3|3|3|4|3|3.33|||||||||2|2|2|2||||||2|3|3|5|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||1|4|3|2.67||||||3|3|3|||||2|2||||4|4||||Red|Cabarrus County|Volunteer: Time constraint|20.1||1|3|1|2|F|White||9|No|Mother|28025|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|Cabarrus County|Pending Match|F|White||68|28025||Married|Retired||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|503694497|503696462|1|0|2|503550540|1|0|2|500828979|2||500016307||4|3|500016374|500016374|-2|500016374|-2|0|4|||7464|9|||1|1005416||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-09|2016-10-28|Followup|2016-06-09|2016-06-20|Complete|Done|4|1|2|2|2|3|2.33|||||||||4|4|4|3|4|3|3.67|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Green|mentor2.0, mentor2.0 2014|Child/Family: Moved|16.7||1|2|1|2|F|White||17|No|Mother|28217|9|One Parent: Female|Unknown|Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|F|White||44|28226|Masters Degree|Single|Human Services: Social Worker|28226|0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017786|504043224|504045242|1|0|2|503985439|1|0|2|500828962|2||500015511||4|1|500014505, 500014506|500014505, 500014506|-2||-2|0|4|||7462|13|||1|902193|799667|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-09|NaT|Followup|2016-06-09|2016-06-30|Complete|Done|2|4|2|4|4|2|3|3|4|4|4|4|4|3.83|-21.67|4|4|4|2|4|4|3.67|4|4|4|4|4|4|4|-8.25|4|4|4|4|4|4|4|4|0|4|3|5|5|4.25|3|5|5|5|4.5|-5.56|4|4|4|4|4|4|3|3.86|4|4|4|4|2|4|3|3.57|8.12|3|4|4|3.67|3|4|2|3|22.33|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green|||20.9||1|2|2|3|F|Black||13|No|Mother|28206|5|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|F|Black||27|28213|Bachelors Degree|Single|Finance|28202|0|5|Ally Financial|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500017732|503996726|503998741|31|0|2|503355514|31|0|2|500829491|2||-2||2|1|||-2||-1|0|4|||12831|3|||1|901778|792064|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-10|2016-10-28|Followup|2016-06-10|2016-06-30|Declined|Done||||||||3|3|3|2|2|3|2.67|||||||||3|4|4|3|3|4|3.5||||||4|4|4|4|||||||4|5|5|5|4.75||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|4|3||||1|1||||4|4||Yellow|mentor2.0, mentor2.0 2014|Child/Family: Lost contact with volunteer/agency|16.6||1|2|1|2|F|Black||17|No|Mother|28217|9|One Parent: Female|Unknown||Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|F|White||31|28278|Bachelors Degree|Married|Business: Mgt, Admin|28202|4|0|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|277|60|598|500000170|500017786|504043260|504045278|31|0|2|503969480|1|0|2|500829872|2||500015511||4|2|500014505, 500014506|500014505, 500014506|-2|500014506|-2|0|4|||7462|13|||1|903076|799585|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-16|2016-06-30|Baseline|2015-05-26|2015-06-16|Complete|Done|4|3|4|2|4|4|3.5|||||||||2|3|3|3|4|4|3.17|||||||||4|4|4|4||||||2|4|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||2|2|2|2||||||4|4|4|||||1|1||||4|4||||Yellow|PERL 2014-2016|Child: Lost interest|12.5||1|1|1|1|F|White||14|No|GrandMother|28277|7|Grandparents|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||30|28273|Bachelors Degree|Single|Business: Engineer|28273|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Enrollment|277|60|598|500000170|500013781|504221476|504223590|1|0|2|504231286|1|0|2|500828128|2||-2||4|2|500014681|500014681|-2|500014681|-2|0|5|||17159|12|||1|888610|-1|4|3|44|5605796235524810842
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Baseline|2015-05-29|2015-06-16|Complete|Done|3|3|4|3|3|4|3.33|||||||||2|4|3|3|2|4|3|||||||||4|3|4|3.67||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||20.7||1|1|1|1|M|Black||13|No|Mother|28216|6|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Business|28217|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504247189|504249305|31|0|1|504228103|1|0|1|500828700|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|892042|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Baseline|2015-06-09|2015-06-16|Complete|Done|4|2|4|4|3|3|3.33|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||1|2|1.5|||||2|2||||4|4||||Green|PERL 2014-2016||20.7||1|1|1|1|M|Black||15|No|GrandMother|28208|7|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|3|10|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503944459|503946467|31|0|1|504260502|1|0|1|500829606|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7462|13|||1|901862|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Followup|2016-06-16|2016-08-18|Declined|Late||||||||4|2|4|4|3|3|3.33|||||||||4|4|4|3|2|4|3.5||||||4|4|4|4|||||||4|3|5|5|4.25||||||||||4|4|4|4|3|4|3|3.71||||||4|4|3|3.67|||||1|2|1.5||||2|2||||4|4||Green|PERL 2014-2016||20.7||1|1|1|1|M|Black||15|No|GrandMother|28208|7|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|3|10|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503944459|503946467|31|0|1|504260502|1|0|1|500829606|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7462|13|||1|905636|901862|4|1|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Followup|2016-06-16|2016-08-31|Expired|Late||||||||3|3|4|3|3|4|3.33|||||||||2|4|3|3|2|4|3||||||4|3|4|3.67|||||||4|4|3|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|3|3||||1|1||||4|4||Green|||20.7||1|1|1|1|M|Black||13|No|Mother|28216|6|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Business|28217|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504247189|504249305|31|0|1|504228103|1|0|1|500828700|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|905690|892042|4|0|45|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-18|2015-12-29|Baseline|2015-05-28|2015-06-18|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|4|3|2|4|3|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||4|3|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|6.4||1|1|1|1|M|Black||13|Yes|Mother|28214|5|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Asian|Indian|49|28203|Bachelors Degree|Married|Tech: Engineer|28204|10|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504217755|504219869|31|0|1|504131744|4|18|1|500828564|2||-2||4|1||500000294|-2||-2|34|2|||17159|12|||1|890821|-1|4|3|44|7000602719972091240
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-18|NaT|Baseline|2015-06-10|2015-06-18|Complete|Done|2|4|4|3|4|3|3.33|||||||||2|4|4|1|1|3|2.5|||||||||4|4|4|4||||||3|2|2|4|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||1|1||||4|4||||Green|PERL 2014-2016||20.6||1|1|1|1|F|Black||15|No|Mother|28212|7|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||31|28204|Masters Degree|Single|Student: College||0|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|502979699|502981150|31|0|2|504127445|1|0|2|500829841|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7464|9|||1|902964|-1|4|3|44|415738029281868742
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-18|NaT|Followup|2016-06-18|2016-08-03|Declined|Late||||||||2|4|4|3|4|3|3.33|||||||||2|4|4|1|1|3|2.5||||||4|4|4|4|||||||3|2|2|4|2.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||2|4|3||||1|1||||4|4||Green|PERL 2014-2016||20.6||1|1|1|1|F|Black||15|No|Mother|28212|7|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||31|28204|Masters Degree|Single|Student: College||0|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|502979699|502981150|31|0|2|504127445|1|0|2|500829841|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7464|9|||1|906912|902964|4|1|45|415738029281868742
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-23|2016-03-03|Baseline|2015-06-23|2015-06-23|Complete|Done|2|4|4|3|3|3|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016|Child/Family: Moved|8.3||1|1|1|1|F|Black||13|No|Mother|28134|6|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||30|28277|Bachelors Degree|Single|Business: Clerical|28277|1|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502205926|502206355|31|0|2|504225335|1|0|2|500831147|2||-2||4|1|500014681|500014681|-2||-2|0|5|||7464|9|||1|908891|-1|4|3|44|6178126991714892144
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-24|2017-02-28|Baseline|2015-06-15|2015-06-24|Complete|Done|4|3|4|2|4|4|3.5|||||||||4|4|4|1|2|4|3.17|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4||||||||3|2|2.5|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|20.2||1|1|1|1|M|Black||12|Yes|Mother|28208|4|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community|Amachi, PERL 2014-2016|Match Support|M|White||30|28202|Masters Degree|Single|Finance: Accountant|28202|0|6|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504054004|504056028|31|0|1|504265163|1|0|1|500830573|2||-2||4|3|500014681|500000294, 500014681|-2||-2|34|2|||17159|12|||1|905463|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-24|2017-02-28|Followup|2016-06-24|2016-06-29|Complete|Done|4|3|4|3|4|4|3.67|4|3|4|2|4|4|3.5|4.86|4|4|4|2|4|4|3.67|4|4|4|1|2|4|3.17|15.77|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3|3|3.25|23.08|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4||||2|3|2.5|3|2|2.5|0|2|2|1|1|100|4|4|4|4|0|Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|20.2||1|1|1|1|M|Black||12|Yes|Mother|28208|4|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community|Amachi, PERL 2014-2016|Match Support|M|White||30|28202|Masters Degree|Single|Finance: Accountant|28202|0|6|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504054004|504056028|31|0|1|504265163|1|0|1|500830573|2||-2||4|3|500014681|500000294, 500014681|-2||-2|34|2|||17159|12|||1|909265|905463|4|3|45|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-25|NaT|Baseline|2015-06-12|2015-06-25|Complete|Done|3|2|1|1|3|4|2.33|||||||||2|2|3|2|3|1|2.17|||||||||1|3|2|2||||||5|3|4|5|4.25||||||||1|4|4|3|4|4|||||||||||4|4|4|4||||||1|2|1.5|||||1|1||||4|4||||Green|PERL 2014-2016||20.4||1|1|1|1|M|Black||16|No|Mother|28208|7|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Hispanic||26|28203|Bachelors Degree|Single|Business: Sales|53073|0|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|503955527|503957535|31|0|1|504285092|3|0|1|500830048|2||-2||2|1|500014681|500014681|-2||-2|0|5|||17159|12|||1|904321|-1|4|3|44|3380017483853696343
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-25|NaT|Followup|2016-06-25|2016-08-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||20.4||3|3|1|1|F|Black||13|No|GrandMother|28227|5|Grandparents|Unknown||No||Self|General Community||Match Support|F|Black||31|28210|Associate Degree|Single|Finance|28255|0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020753|502252822|502253254|31|0|2|504229640|31|0|2|500829933|2||-2||2|1|||-2||-2|0|10|||7671|13|||1|909577||4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-25|NaT|Followup|2016-06-25|2016-06-29|Complete|Done|2|2|2|2|3|3|2.33|3|2|1|1|3|4|2.33|0|2|3|2|2|3|2|2.33|2|2|3|2|3|1|2.17|7.37|2|2|2|2|1|3|2|2|0|3|2|2|3|2.5|5|3|4|5|4.25|-41.18|3|2|4|4|3|4|3|3.29||1|4|4|3|4|4|||4|4|4|4|4|4|4|4|0|2|2|2|1|2|1.5|33.33|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||20.4||1|1|1|1|M|Black||16|No|Mother|28208|7|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Hispanic||26|28203|Bachelors Degree|Single|Business: Sales|53073|0|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|503955527|503957535|31|0|1|504285092|3|0|1|500830048|2||-2||2|1|500014681|500014681|-2||-2|0|5|||17159|12|||1|909731|904321|4|3|45|3380017483853696343
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-26|2017-02-28|Followup|2016-06-26|2016-08-03|Complete|Done|3|4|4|4|2|3|3.33|2|1|2|1|1|1|1.33|150.38|2|4|3|1|1|4|2.5|3|1|3|1|1|3|2|25|4|2|2|2.67|4|4|4|4|-33.25|1|1|1|3|1.5|3|5|3|4|3.75|-60|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|3|3|2|2.67|1|3|1|1.67|59.88|4|2|3|1|2|1.5|100|2|2|1|1|100|4|4|4|4|0|Green||Child/Family: Lost contact with volunteer/agency|20.1||1|2|2|3|F|Black||14|No|Father|28205|6|One Parent: Male|Unknown||Yes||School|General Community||Match Support|F|White||49|28278|Masters Degree|Single|Business|28202|12|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500017732|503624326|503626215|31|0|2|503605964|1|0|2|500831308|2||-2||4|1|||-2||-1|0|4|||16705|3|||1|910195|661637|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-27|NaT|Baseline|2015-06-15|2015-06-27|Complete|Done|4|4|3|4|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|1|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Green|Cabarrus County||20.3||1|1|1|1|M|Multi-race (Black & Asian)||12|No|Mother|28025|7|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Asian||32|28025|Bachelors Degree|Married|Tech: Sales, Mktg|28202|8|9|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi, Cabarrus County, mentor2.0|Match Support|277|60|598|500000170|500022817|504051660|504053684|39|0|1|504277513|4|0|1|500830267|2||500016307||2|1|500016374|500016374|-2|500000294, 500014505, 500016374|-2|0|10|||7462|13|||1|905458|-1|4|3|44|887254134148570071
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-27|NaT|Followup|2016-06-27|2016-07-25|Complete|Done|2|1|1|1|1|2|1.33|4|4|3|4|4|4|3.83|-65.27|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|3|5|4.5|5|5|1|5|4|12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|3|3|3|1|1|1|200|2|2|2|2|0|4|4|4|4|0|Green|Cabarrus County||20.3||1|1|1|1|M|Multi-race (Black & Asian)||12|No|Mother|28025|7|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Asian||32|28025|Bachelors Degree|Married|Tech: Sales, Mktg|28202|8|9|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi, Cabarrus County, mentor2.0|Match Support|277|60|598|500000170|500022817|504051660|504053684|39|0|1|504277513|4|0|1|500830267|2||500016307||2|1|500016374|500016374|-2|500000294, 500014505, 500016374|-2|0|10|||7462|13|||1|910458|905458|4|3|45|887254134148570071
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-28|2016-02-24|Baseline|2015-06-28|2015-06-28|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red|PERL 2014-2016|Child/Family: Time constraints|7.9||1|1|2|2|M|Black||11|No|Mother|28226|3|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|504198439|504200550|31|0|1|504230177|1|0|1|500831539|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||7462|13|||1|910542|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-29|2015-09-23|Baseline|2015-06-16|2015-06-29|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|3|1|2|4|3|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|2|3.71||||||||||3|4|4|3.67||||||3|1|2|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|2.8||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28031||Single|Service: Restaurant|28078|0|2|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504186384|1|0|1|500830331|2||-2||4|3|500014681|500014681|-2|500000294, 500014681|-2|0|4|||7464|9|||1|905704|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-29|2016-09-27|Followup|2016-06-29|2016-08-19|Declined|Late||||||||3|1|4|4|3|4|3.17|||||||||4|3|4|2|1|4|3||||||4|3|3|3.33|||||||5|4|4|4|4.25||||||||||4|4|4|4|3|4|2|3.57||||||3|4|1|2.67|||||1|1|1||||2|2||||4|4||Red||Child/Family: Time constraints|15||2|2|1|1|F|Some Other Race||15|No|Aunt|28217|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||36|28210|Masters Degree|Single|Finance: Accountant|28202|6|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|502612404|500188044|41|0|2|504226710|1|0|2|500830721|2||-2||4|3|||-2||-2|0|10|||17159|12|||1|911353|788378|4|1|45|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-29|NaT|Baseline|2015-05-14|2015-06-29|Complete|Done|2|3|2|3|2|2|2.33|||||||||1|2|2|3|2|3|2.17|||||||||4|4|4|4||||||2|4|4|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|2|3||||||4|4|4|||||1|1||||4|4||||Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016||20.3||1|1|1|1|F|Hispanic||15|No|Mother|28215|9|One Parent: Female|Unknown||Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|White||45|28205|Associate Degree|Married|Tech: Computer/Programmer|28202|10|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504154291|504156341|3|0|2|503862054|1|0|2|500827743|2||-2||2|1|500011312, 500014681|500011312, 500014681|-2|500014681|-2|0|10|||17159|12|||1|881920|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-29|NaT|Followup|2016-06-29|2016-08-25|Declined|Late||||||||2|3|2|3|2|2|2.33|||||||||1|2|2|3|2|3|2.17||||||4|4|4|4|||||||2|4|4|5|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|3|2|3|||||4|4|4||||1|1||||4|4||Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016||20.3||1|1|1|1|F|Hispanic||15|No|Mother|28215|9|One Parent: Female|Unknown||Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|White||45|28205|Associate Degree|Married|Tech: Computer/Programmer|28202|10|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504154291|504156341|3|0|2|503862054|1|0|2|500827743|2||-2||2|1|500011312, 500014681|500011312, 500014681|-2|500014681|-2|0|10|||17159|12|||1|911350|881920|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-06-30|2016-08-22|Followup|2016-06-30|2016-06-28|Complete|Done|2|3|4|4|3|3|3.17|||||||||3|2|4|2|3|4|3|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Infraction of match rules/agency policies|13.8||1|1|2|2|M|White||10|No|Mother|28277|3|One Parent: Female|$40,000 to $44,999|Y|Yes||Self|General Community||Match Support|M|White||57|28105|Bachelors Degree|Married|Business: Sales|28203|11|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503921502|503891297|1|0|1|504063702|1|0|1|500831159|2||-2||4|1|||-2|500000294|-2|0|10|||17159|12|||1|912398||4|3|45|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-16|NaT|Followup|2016-07-16|2016-07-25|Complete|Done|2|3|4|4|3|2|3|3|4|4|4|3|3|3.5|-14.29|3|4|4|4|3|4|3.67|3|4|4|3|1|4|3.17|15.77|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|4|3|3|4|3.5|-7.14|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|||19.7||1|2|1|2|F|Black||17|No|Mother|28208|9|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|F|Black||27|28202|Masters Degree|Single|Business|28202|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|277|60|598|500000170|500017732|504042339|504044357|31|0|2|503984783|31|0|2|500833563|2||-2||2|1|||-2|500014506|-2|0|4|||7462|13|||1|916498|800017|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-17|2016-10-21|Baseline|2015-06-11|2015-07-17|Complete|Done|3|1|3|1|3|4|2.5|||||||||1|4|3|3|3|3|2.83|||||||||4|4|4|4||||||4|2|4|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Time constraint|15.2||1|1|1|1|F|Black||13|No|Mother|28213|5|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||28|28078|Bachelors Degree|Single|Business|28078|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504218954|504221068|31|0|2|504099424|1|0|2|500830251|2||-2||4|3|500014681|500014681|-2||-2|0|4|||46|2|||1|903482|-1|4|3|44|6178126991714892144
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-17|2016-10-21|Followup|2016-07-17|2016-08-30|Complete|Done|3|3|3|3|4|4|3.33|3|1|3|1|3|4|2.5|33.2|4|4|4|3|4|4|3.83|1|4|3|3|3|3|2.83|35.34|4|4|4|4|4|4|4|4|0|4|4|3|4|3.75|4|2|4|4|3.5|7.14|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|3|3.67|0|3|3|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Red|PERL 2014-2016|Volunteer: Time constraint|15.2||1|1|1|1|F|Black||13|No|Mother|28213|5|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||28|28078|Bachelors Degree|Single|Business|28078|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504218954|504221068|31|0|2|504099424|1|0|2|500830251|2||-2||4|3|500014681|500014681|-2||-2|0|4|||46|2|||1|916932|903482|4|3|45|6178126991714892144
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-23|2017-02-28|Followup|2016-07-23|2016-09-01|Declined|Done||||||||4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4||||||4|4|4|4|||||||4|4|3|4|3.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Yellow|PERL 2014-2016|Volunteer: Time constraint|19.3||1|2|1|2|F|Black||14|No|Mother|28205|6|One Parent: Female|Unknown||Yes||School|General Community|PERL 2014-2016|Match Support|F|White||31|28211|Masters Degree|Single|Finance: Accountant|28202|1|0|Duke Energy|Workplace Partner|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|504012972|504014987|31|0|2|503975669|1|0|2|500834251|2||-2||4|2|500014681|500014681|-2|500014681|-2|0|4|||16705|3|||1|918234|793644|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-23|NaT|Baseline|2015-07-23|2015-07-23|Complete|Done|4|3|4|1|4|4|3.33|||||||||2|3|3|2|1|4|2.5|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|||19.5||1|1|1|1|M|Black||15|No|Mother|28215|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||31|28202|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|504220177|504222291|31|0|1|504309758|1|0|1|500834242|2||-2||2|1|||-2||-2|0|4|||46|2|||1|918218|-1|4|3|44|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-23|NaT|Followup|2016-07-23|2016-10-07|Expired|Late||||||||4|3|4|1|4|4|3.33|||||||||2|3|3|2|1|4|2.5||||||4|4|4|4|||||||3|4|4|5|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|4|3.5||||2|2||||4|4||Green|||19.5||1|1|1|1|M|Black||15|No|Mother|28215|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||31|28202|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|504220177|504222291|31|0|1|504309758|1|0|1|500834242|2||-2||2|1|||-2||-2|0|4|||46|2|||1|918387|918218|4|0|45|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-23|NaT|Followup|2016-07-23|2016-07-22|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||19.5||2|2|1|1|F|Black||10||Mother|28216|4|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Business: Human Resources|28202|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|503259551|503261359|31|0|2|504219483|1|0|2|500831431|2||-2||2|1|||-2||-2|34|2|||7496|10|||1|933116||4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-27|2017-01-18|Baseline|2015-07-11|2015-07-27|Complete|Done|1|1|1|1|3|2|1.5|||||||||4|1|4|4|2|3|3|||||||||4|4|4|4||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|17.8||1|1|1|1|F|Black||10|No|Mother|28208|3|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Enrollment|F|Black||24|28262||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504274120|504276320|31|0|2|504255905|31|0|2|500832878|2||-2||4|3|||-2||-2|0|4|||17159|12|||1|914893|-1|4|3|44|2053394993324953440
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-27|2017-01-18|Followup|2016-07-27|2016-09-01|Complete|Done|3||3|2|4|3||1|1|1|1|3|2|1.5||4|4|4|4|4|4|4|4|1|4|4|2|3|3|33.33|4|4|4|4|4|4|4|4|0|4|4|4|4|4|5|4|3|3|3.75|6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|3|3.67|8.99|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|17.8||1|1|1|1|F|Black||10|No|Mother|28208|3|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Enrollment|F|Black||24|28262||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504274120|504276320|31|0|2|504255905|31|0|2|500832878|2||-2||4|3|||-2||-2|0|4|||17159|12|||1|919087|914893|4|3|45|2053394993324953440
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Baseline|2015-07-16|2015-07-27|Complete|Done|3|3|4|4|3|4|3.5|||||||||4|4|4|4|2|4|3.67|||||||||3|3|3|3||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green|||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||Relative|General Community||Match Support|F|White||29|28209|Bachelors Degree|Single|Retail: Mgt|28217|3|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504312629|504314787|31|0|2|504262612|1|0|2|500833665|2||-2||2|1|||-2||-2|0|3|||17159|12|||1|916650|-1|4|3|44|237874676114443178
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Baseline|2015-07-20|2015-07-27|Complete|Done|4|4|4|4|1|4|3.5|||||||||2|2|2|2|3|2|2.17|||||||||3|3|3|3||||||3|3|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Asian||28|28203|Bachelors Degree|Single|Consultant|28202|1|1|Current/Previous Big|Other Big|Big|General Community|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500008321|504312569|504314787|31|0|2|504208036|4|0|2|500833808|2||-2||2|1|500014681|500014681|-2|500014505, 500015184|-2|0|4|||17159|12|||1|917230|-1|4|3|44|237874676114443178
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Followup|2016-07-27|2016-09-01|Complete|Done|3|4|4|4|3|4|3.67|3|3|4|4|3|4|3.5|4.86|4|3|4|4|4|4|3.83|4|4|4|4|2|4|3.67|4.36|4|4|4|4|3|3|3|3|33.33|3|4|3|4|3.5|4|5|5|4|4.5|-22.22|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|4|3|3.33|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green|||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||Relative|General Community||Match Support|F|White||29|28209|Bachelors Degree|Single|Retail: Mgt|28217|3|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504312629|504314787|31|0|2|504262612|1|0|2|500833665|2||-2||2|1|||-2||-2|0|3|||17159|12|||1|918944|916650|4|3|45|237874676114443178
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Followup|2016-07-27|2016-09-01|Complete|Done|4|4|4|4|4|4|4|4|4|4|4|1|4|3.5|14.29|3|4|4|4|4|4|3.83|2|2|2|2|3|2|2.17|76.5|4|3|3|3.33|3|3|3|3|11|4|4|4|3|3.75|3|3|5|5|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|3|4|4|3.67|-18.26|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Asian||28|28203|Bachelors Degree|Single|Consultant|28202|1|1|Current/Previous Big|Other Big|Big|General Community|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500008321|504312569|504314787|31|0|2|504208036|4|0|2|500833808|2||-2||2|1|500014681|500014681|-2|500014505, 500015184|-2|0|4|||17159|12|||1|918957|917230|4|3|45|237874676114443178
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-28|2016-05-26|Baseline|2015-07-10|2015-07-28|Complete|Done|3|1|4|2|4|3|2.83|||||||||2|4|3|1|3|3|2.67|||||||||4|3|4|3.67||||||3|5|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2||||4|4||||Yellow|PERL 2014-2016|Changing Match Type|10||1|3|1|3|F|Black||15|No|Mother|28208|8|One Parent: Female|$10,000 to $14,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|Multi-race (Black & White)||41|28216||Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community|mentor2.0|Match Support|277|60|598|500000170|500008321|504308876|504311094|31|0|2|504215512|36|0|2|500833533|2||-2||4|2|500014681|500014681|-2|500014505|-2|34|2|||46|2|||1|914712|-1|4|3|44|2806833304218536184
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-28|2017-02-26|Followup|2016-07-28|2016-08-25|Declined|Done||||||||1|1|3|1|2|3|1.83|||||||||1|1|3|2|3|3|2.17||||||2|4|2|2.67|||||||3|5|4|3|3.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|4|3||||2|2||||4|4||Red||Volunteer: Lost contact with child/agency|19||1|2|1|2|F|Hispanic||13|No|Mother|28217|3|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|F|White||45|28273|Some College|Single|Business|28217|2|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503779471|503781448|3|0|2|503040015|1|0|2|500834596|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|919303|698543|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-28|2016-01-11|Baseline|2015-07-28|2015-07-28|Complete|Done|3|4|4|4|4|3|3.67|||||||||3|4|3|2|3|3|3|||||||||4|4|4|4||||||2|4|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|5.5||1|1|1|1|F|Black||13|No|Mother|28217|6|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Finance: Banking||2|2|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500018851|504230613|503065429|31|0|2|503995309|1|0|2|500834694|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|919515|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-28|NaT|Followup|2016-07-28|2016-07-31|Complete|Done|3|3|3|2|3|4|3|||||||||3|3|3|2|2|2|2.5|||||||||3|3|3|3||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|||19.3||1|1|1|1|M|Black||10||GrandMother|28213|2|Grandparents|Unknown|Y|Yes||Self|General Community||Match Support|M|White||28|28204||Single|Finance: Accountant|28277|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|503022461|501332937|31|0|1|504323998|1|0|1|500834322|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|980040||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-30|2016-01-07|Baseline|2015-07-30|2015-07-30|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|2|2|2|3|2.5|||||||||4|4|4|4||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|5.3||1|1|1|1|M|Black||14|No|Mother|28217|6|One Parent: Female|$10,000 to $14,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||31|28209|Bachelors Degree|Single|Human Services|28203|1|8|Current/Previous Big|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500018851|503063769|503065429|31|0|1|504299841|1|0|1|500834948|2||-2||4|2|||-2||-2|34|2|||17159|12|||1|920327|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-07-30|2016-02-02|Baseline|2015-07-30|2015-07-30|Complete|Done|2|4|4|4|4|4|3.67|||||||||3|3|3|3|2|3|2.83|||||||||4|4|4|4||||||2|3|4|4|3.25|||||||4|4|4|3|2|3|3|3.29||||||||||2|2|2|2||||||3|4|3.5|||||1|1||||4|4||||Green||Volunteer: Feels incompatible with child/family|6.1||1|1|1|1|M|Black||15|No|Mother|28215|7|One Parent: Female|$60,000 to $74,999||No||School|General Community||Match Support|M|Black||52|28273|Bachelors Degree|Single|Self-Employed, Entrepreneur||25|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501401583|501401868|31|0|1|504338671|31|0|1|500834950|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|920331|-1|4|3|44|3003539216843226222
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-04|NaT|Followup|2016-08-04|2016-08-10|Complete|Done|1|3|2|1|4|3|2.33|4|4|4|1|4|4|3.5|-33.43|3|3|4|2|2|4|3|2|4|4|1|4|4|3.17|-5.36|4|4|4|4|3|2|3|2.67|49.81|4|4|4|3|3.75|4|5|3|4|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3|3.71|7.82|4|4|4|4|4|3|4|3.67|8.99|3|3|3|1|2|1.5|100|2|2|1|1|100|4|4|4|4|0|Green|||19.1||2|2|1|1|M|Black||12|No|Mother|28212|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||27|28211|Bachelors Degree|Married|Finance: Banking|28211|0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|503565188|503567063|31|0|1|504265907|1|0|1|500831744|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|923934|725936|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-08-11|2015-11-30|Baseline|2015-08-06|2015-08-11|Complete|Done|4|4|2|2|4|4|3.33|||||||||3|4|3|3|4|3|3.33|||||||||3|3|4|3.33||||||2|4|5|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Feels incompatible with child/family|3.6||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28212|6|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community|PERL 2014-2016|Enrollment|F|White||47|28270|Some College|Married|Homemaker|29020|18|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|504280484|504282684|36|0|2|504226821|1|0|2|500835375|2||-2||4|3|500014681|500014681|-2||-2|0|3|||7464|9|||1|924522|-1|4|3|44|4694273237201497095
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-13|NaT|Baseline|2015-08-13|2015-08-13|Complete|Done|4|2|3|2|4|4|3.17|||||||||3|3|4|2|3|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|||18.8||1|1|1|1|F|Black||13|No|Mother|28214|6|One Parent: Female|$50,000 to $59,999||Yes||Self|General Community||Match Support|F|White||29|28273|Masters Degree|Married|Finance: Accountant|28210|3|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504328960|504331182|31|0|2|504215323|1|0|2|500836079|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|926159|-1|4|3|44|8503368421346667831
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-13|NaT|Followup|2016-08-13|2016-08-22|Complete|Done|4|3|3|2|4|4|3.33|4|2|3|2|4|4|3.17|5.05|3|4|4|4|4|4|3.83|3|3|4|2|3|4|3.17|20.82|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|5|5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|3|3|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Green|||18.8||1|1|1|1|F|Black||13|No|Mother|28214|6|One Parent: Female|$50,000 to $59,999||Yes||Self|General Community||Match Support|F|White||29|28273|Masters Degree|Married|Finance: Accountant|28210|3|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504328960|504331182|31|0|2|504215323|1|0|2|500836079|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|926293|926159|4|3|45|8503368421346667831
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-13|NaT|Followup|2016-08-13|2016-09-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||18.8||1|1|1|1|F|Black||10|No|Mother|28216|2|One Parent: Female|$30,000 to $34,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||34|28031||Single|Self-Employed, Entrepreneur||9|8|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504186133|504188242|31|0|2|504122609|1|0|2|500834256|2||-2||2|1|||-2||-2|34|2|||17159|12|||1|937690||4|1|45|8136849793711030748
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-14|NaT|Baseline|2015-07-22|2015-08-14|Complete|Done|2|3|3|3|3|2|2.67|||||||||4|4|4|2|2|4|3.33|||||||||4|4|4|4||||||5|4|4|2|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||3|3||||Green|||18.8||1|1|1|1|M|Black||13|No|Mother|28273|6|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|Black||56|28273|Some College|Married|Govt|28228|0|7|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|504284556|504286757|31|0|1|504260574|31|0|1|500834204|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|918085|-1|4|3|44|2392572474128905139
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-14|NaT|Followup|2016-08-14|2016-09-28|Complete|Done|4|4|4|2|3|3|3.33|2|3|3|3|3|2|2.67|24.72|2|4|3|3|4|3|3.17|4|4|4|2|2|4|3.33|-4.8|4|4|4|4|4|4|4|4|0|3|3|4|3|3.25|5|4|4|2|3.75|-13.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|3|3.33|4|4|3|3.67|-9.26|2|3|2.5|2|2|2|25|2|2|2|2|0|4|4|3|3|33.33|Green|||18.8||1|1|1|1|M|Black||13|No|Mother|28273|6|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|Black||56|28273|Some College|Married|Govt|28228|0|7|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|504284556|504286757|31|0|1|504260574|31|0|1|500834204|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|926429|918085|4|3|45|2392572474128905139
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-08-20|2015-12-30|Baseline|2015-06-11|2015-08-20|Complete|Done|2|2|4|1|4|4|2.83|||||||||1|3|2|1|1|3|1.83|||||||||3|2|2|2.33||||||3|4|3|3|3.25|||||||4|2|4|4|4|2|2|3.14||||||||||3|3|2|2.67||||||1|4|2.5|||||1|1||||3|3||||Green||Child/Family: Moved|4.3||1|1|1|1|F|Black||15|No|Mother|28215|8|Two Parent|Unknown||Yes||Self|General Community||Match Support|F|Multi-race (Black & Asian)||23|28206|High School Graduate|Single|Business|28273|1|6|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|277|60|598|500000170|500020990|504207073|504025357|31|0|2|504201268|39|0|2|500829987|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|903693|-1|4|3|44|6720484407795402036
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-20|NaT|Followup|2016-08-20|2016-10-11|Declined|Late||||||||4|4|4|4|4|4|4|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||4|5|3|4|4||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||2|1|1.5||||1|1||||4|4||Green|||18.6||2|2|3|3|M|American Indian or Alaska Native||14|No|Mother|28269|7|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Asian||27|28202|Bachelors Degree|Single|Finance|28202|0|1|Current/Previous Big|Other Big|Big|General Site||Match Support|277|60|598|500000170|500020752|504150667|504152735|6|0|1|504242094|4|0|1|500836074|2||-2||2|1||500014681|-2||-1|0|4|||17159|12|||1|927866|886556|4|1|45|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-08-22|2016-05-17|Baseline|2015-07-24|2015-08-22|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Volunteer: Lost contact with child/agency|8.8||1|1|1|1|F|Black||12|No|Mother|28214|4|One Parent: Female|Unknown|Y|Yes||School|General Community|Amachi|Match Support|F|Asian||33|28205|Bachelors Degree|Single|Consultant|60654|2|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|504166613|504168697|31|0|2|503823941|4|0|2|500834370|2||-2||4|1|500000294|500000294|-2||-2|0|4|||7464|9|||1|918534|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-25|NaT|Followup|2016-08-25|2016-10-19|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||18.4||1|1|1|1|M|Black||9|No|Mother|28262|2|One Parent: Female|$30,000 to $34,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||40|28202|Bachelors Degree|Single|Self-Employed, Entrepreneur||7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|503967629|503969639|31|0|1|504276405|1|0|1|500834265|2||-2||2|1|||-2||-2|34|2|||46|2|||1|1040735||4|1|45|6619197389800008587
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-08-30|2015-12-30|Baseline|2015-08-10|2015-08-30|Complete|Done|3|1|4|1|1|3|2.17|||||||||2|1|3|1|2|4|2.17|||||||||1|2|2|1.67||||||3|4|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016|Child/Family: Moved|4||1|1|1|1|F|Black||12|No|Mother|28212|4|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||33|28270|Some College|Single|Business|28262|1|3|Other|BBBS Board/Staff|Big|General Community||Enrollment|277|60|598|500000170|500017732|504343306|504345530|31|0|2|504109000|31|0|2|500835668|2||-2||4|1|500014681|500014681|-2||-2|0|10|||7671|13|||1|925217|-1|4|3|44|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-08|NaT|Followup|2016-09-08|2016-09-12|Complete|Done|2|3|3|3|4|4|3.17|1|4|4|4|3|4|3.33|-4.8|2|||3|2|||2|3|4|4|2|3|3||||||4|4|4|4||3|3|3|4|3.25|3|3|3|4|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|||||3|4|2|3||3|3|3|2|4|3|0|2|2|2|2|0|4|4|4|4|0|Green|||17.9||1|2|1|2|F|Black||16|No|Mother|28205|9|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|F|Black||46|28214|Associate Degree|Married|Business|28202|2|10|Duke Energy|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500018851|503633704|503635645|31|0|2|503604638|31|0|2|500835662|2||-2||2|1|||-2||-2|0|4|||16705|3|||1|932233|663231|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-10|NaT|Baseline|2015-08-24|2015-09-10|Complete|Done|4|1|2|1|4|4|2.67|||||||||2|4|4|1|1|3|2.5|||||||||4|4|4|4||||||4|5|2|2|3.25|||||||4|1|4|4|2|4|4|3.29||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016||17.9||1|1|1|1|M|Black||11|No|Mother|28203|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28202|Bachelors Degree|Single|Retail: Sales|28209|4|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504039192|504041210|31|0|1|504344501|1|0|1|500837420|2||-2||2|1|500014681|500014681|-2||-2|0|4|||17159|12|||1|928481|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-10|NaT|Followup|2016-09-10|2016-11-09|Complete|Late|4|1|3|2|4|4|3|4|1|2|1|4|4|2.67|12.36|3|4|3|2|2|2|2.67|2|4|4|1|1|3|2.5|6.8|4|4|4|4|4|4|4|4|0|4|3|2|4|3.25|4|5|2|2|3.25|0|4|4|4|4|4|4|4|4|4|1|4|4|2|4|4|3.29|21.58|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||17.9||1|1|1|1|M|Black||11|No|Mother|28203|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28202|Bachelors Degree|Single|Retail: Sales|28209|4|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504039192|504041210|31|0|1|504344501|1|0|1|500837420|2||-2||2|1|500014681|500014681|-2||-2|0|4|||17159|12|||1|932966|928481|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-13|NaT|Followup|2016-09-13|2016-10-12|Complete|Done|4|2|3|1|4|3|2.83|4|1|2|1|3|4|2.5|13.2|1|4|4|2|2|4|2.83|1|3|4|2|3|2|2.5|13.2|4|4|4|4|3|4|4|3.67|8.99|4|4|3|5|4|3|4|5|4|4|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|2|1|1.5|100|2|2|2|2|0|4|4|4|4|0|Green|||17.8||3|3|1|1|F|Black||14|No|GrandMother|28215|8|Grandparents|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|F|White||23|28202||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|502583662|502584168|31|0|2|504286292|1|0|2|500836763|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|933630|621292|4|3|45|3959612471441160400
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-16|NaT|Baseline|2015-09-10|2015-09-16|Complete|Done|4|4|4|4|3|4|3.83|||||||||3|4|4|2|4|4|3.5|||||||||3|3|4|3.33||||||4|3|4|2|3.25|||||||4|4|4|3|4|4|4|3.86||||||||||1|1|3|1.67||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016||17.7||1|1|1|1|M|Some Other Race||13|No|Mother|28217|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||38|28205|Masters Degree|Married|Human Services: Social Worker|28204|5|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504155180|501093096|41|0|1|502462446|1|0|1|500839295|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7464|9|||1|932973|-1|4|3|44|358434295995756137
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-16|NaT|Followup|2016-09-16|2016-09-19|Complete|Done|4|4|4|4|4|4|4|4|4|4|4|3|4|3.83|4.44|4|4|4|4|2|4|3.67|3|4|4|2|4|4|3.5|4.86|4|2|2|2.67|3|3|4|3.33|-19.82|5|4|5|4|4.5|4|3|4|2|3.25|38.46|4|4|4|4|4|4|3|3.86|4|4|4|3|4|4|4|3.86|0|4|4|1|3|1|1|3|1.67|79.64|3|3|3|4|4|4|-25|1|1|2|2|-50|4|4|4|4|0|Green|PERL 2014-2016||17.7||1|1|1|1|M|Some Other Race||13|No|Mother|28217|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||38|28205|Masters Degree|Married|Human Services: Social Worker|28204|5|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504155180|501093096|41|0|1|502462446|1|0|1|500839295|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7464|9|||1|934749|932973|4|3|45|358434295995756137
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-21|NaT|Followup|2016-09-21|2016-09-19|Complete|Done|4|4|4|2|4|4|3.67|3|3|4|2|3|4|3.17|15.77|2|4|3|2|2|3|2.67|3|3|4|3|4|3|3.33|-19.82|4|4|4|4|4|3|3|3.33|20.12|5|4|5|5|4.75|4|4|3|3|3.5|35.71|4|4|4|4|3|4|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|2|3|3|2.67|37.45|3|3|3|3|3|3|0|2|2|1|1|100|4|4|4|4|0|Green|||17.5||1|2|1|2|F|Black||12|Yes|Mother|28217|4|One Parent: Female|Unknown||Yes||School|General Community|Amachi|Match Support|F|Black||78|28273|Masters Degree|Widowed|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503807530|503809507|31|0|2|503381588|31|0|2|500841214|2||-2||2|1||500000294|-2||-2|0|4|||7464|9|||1|935881|713201|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-22|NaT|Followup|2016-09-22|2016-10-31|Declined|Done||||||||3|1|3|1|4|4|2.67|||||||||2|4|3|1|2|2|2.33||||||4|4|4|4|||||||2|5|3|2|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4||||1|1||||4|4||Green|PERL 2014-2016||17.5||2|2|1|1|F|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||Yes||School|General Community|PERL 2014-2016|Match Support|F|White||26|28202|Bachelors Degree|Single|Finance: Banking|28262|1|7|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|504013056|504015071|31|0|2|504219921|1|0|2|500839610|2||-2||2|1|500014681|500014681|-2||-2|0|4|||17159|12|||1|936088|793476|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-09-23|2015-12-29|Baseline|2015-09-11|2015-09-23|Complete|Done|4|2|4|2|4|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|Amachi|Child: Lost interest|3.2||1|1|1|1|F|Black||10|Yes|GrandMother|28217|4|Grandparents|Less than $10,000|Y|Yes||School|General Community|Amachi|Match Support|F|White||32|28277|Masters Degree|Divorced|Tech: Computer/Programmer|28277|0|3|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|504195472|504197572|31|0|2|504222207|1|0|2|500839514|2||-2||4|1|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|933343|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-23|NaT|Followup|2016-09-23|2016-10-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|PERL 2014-2016||17.4||2|2|1|1|M|Black||10|No|Mother|28214|2|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||25|28227|Bachelors Degree|Single|Insurance|28277|1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|503779386|503781363|31|0|1|504333970|31|0|1|500839160|2||-2||2|1|500014681|500014681|-2||-2|0|4|||7464|9|||1|936510||4|1|45|1546374315672654438
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-28|NaT|Followup|2016-09-28|2016-10-26|Complete|Done|1|2|4|2|3|3|2.5|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4||4|||||||||4|4|4|4|3|4|3|3.71||||||||||2|3|2|2.33||||||3|4|3.5|||||2|2||||4|4||||Green|||17.3||3|3|1|1|F|Black||14|No|Mother|28216|7|Two Parent|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|White||43|28269|Masters Degree|Single|Business: Mgt, Admin||0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|502186245|501610196|31|0|2|504248899|1|0|2|500836970|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|938163||4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-29|NaT|Baseline|2015-09-23|2015-09-29|Complete|Done|4|1|4|4|2|4|3.17|||||||||1|3|3|1|1|3|2|||||||||3|2|2|2.33||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||17.2||1|1|1|1|M|Black||11|No|Mother|28214|4|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28273|Bachelors Degree|Single|Insurance|28226|7|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|504153965|504156015|31|0|1|504372591|1|0|1|500841770|2||-2||2|1|500014681|500014681|-2||-2|0|4|||7464|9|||1|936574|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-29|NaT|Followup|2016-09-29|2016-11-28|Declined|Late||||||||4|1|4|4|2|4|3.17|||||||||1|3|3|1|1|3|2||||||3|2|2|2.33|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||4|3|3.5||||2|2||||4|4||Green|PERL 2014-2016||17.2||1|1|1|1|M|Black||11|No|Mother|28214|4|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28273|Bachelors Degree|Single|Insurance|28226|7|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|504153965|504156015|31|0|1|504372591|1|0|1|500841770|2||-2||2|1|500014681|500014681|-2||-2|0|4|||7464|9|||1|938480|936574|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Baseline|2015-09-24|2015-10-05|Complete|Done|3|2|3|2|4|4|3|||||||||2|4|4|3|3|4|3.33|||||||||3|3|4|3.33||||||5|4|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|||||||2|2||||4|4||||Green|||17.1||1|1|1|1|F|Black||12|No|Mother|28215|6|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Multi-Race (None of the above)||27|28269|Bachelors Degree|Single|Transport: Flight Attendant|28208|1|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504358312|504320644|31|0|2|504048355|7|0|2|500842174|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|937130|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Baseline|2015-09-28|2015-10-05|Complete|Done|4|2|4|1|2|4|2.83|||||||||4|4|3|1|2|2|2.67|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||1|1||||4|4||||Green|||17.1||1|1|1|1|M|Black||10|No|Mother|28213|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Consultant|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504179804|504181918|31|0|1|504337207|1|0|1|500842586|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|937970|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Followup|2016-10-05|2016-12-20|Expired|Late||||||||4|2|4|1|2|4|2.83|||||||||4|4|3|1|2|2|2.67||||||4|4|4|4|||||||3|5|5|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|1|1.5||||1|1||||4|4||Green|||17.1||1|1|1|1|M|Black||10|No|Mother|28213|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Consultant|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504179804|504181918|31|0|1|504337207|1|0|1|500842586|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|940706|937970|4|0|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Followup|2016-10-05|2016-11-18|Complete|Done|3|3|3|2|4|4|3.17|3|2|3|2|4|4|3|5.67|3|4|4|4|4|3|3.67|2|4|4|3|3|4|3.33|10.21|4|4|4|4|3|3|4|3.33|20.12|4|4|3|4|3.75|5|4|4|3|4|-6.25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|4|4|-8.25|3|3|3|3||||2|2|2|2|0|3|3|4|4|-25|Green|||17.1||1|1|1|1|F|Black||12|No|Mother|28215|6|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Multi-Race (None of the above)||27|28269|Bachelors Degree|Single|Transport: Flight Attendant|28208|1|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504358312|504320644|31|0|2|504048355|7|0|2|500842174|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|940717|937130|4|3|45|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-09|NaT|Followup|2016-10-09|2016-10-08|Complete|Done|3|1|4|2|4|3|2.83|||||||||4|4|4|4|4|4|4|||||||||4|3|3|3.33||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||16.9||2|3|3|3|F|American Indian or Alaska Native||13|No|Aunt|28027|3|Other Relative|Unknown||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||50|28075|Bachelors Degree|Married|Education: Admin|28083|0|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|503012569|504347632|6|0|2|502949193|1|0|2|500841835|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||7671|13|||1|943030||4|3|45|1791051703918408849
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-13|NaT|Followup|2016-10-13|2016-10-11|Complete|Done|3|4|2|2|3|4|3|1|1|1|4|4|4|2.5|20|2|3|3|2|2|3|2.5|2|2|3|3|3|4|2.83|-11.66|4|4|4|4|4|4|4|4|0|3|4|3|4|3.5|5|5|5|3|4.5|-22.22|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|1|4|1|2|83.5|3|2|2.5|4|1|2.5|0|2|2|2|2|0|4|4|4|4|0|Green|||16.8||2|2|1|1|F|Black||11|No|Mother|28269|5|One Parent: Female|$50,000 to $59,999|Y|No||School|General Community||Match Support|F|Black||41|28216|Bachelors Degree|Single|Business|28282|2|11|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|504243465|504245581|31|0|2|504365625|31|0|2|500844251|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|944405|873076|4|3|45|2806833304218536184
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-10-19|2016-10-21|Baseline|2015-10-05|2015-10-19|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|4|3|3|4|3|3.33|||||||||3|3|3|3||||||4|2|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Feels incompatible with child/family|12.1||2|2|1|1|F|Black||11|No|Mother|28203|6|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|F|White||33|28210|PHD|Single|Medical|28105|1|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|504388136|504390375|31|0|2|504360253|1|0|2|500844373|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|940908|-1|4|3|44|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-10-20|2016-11-17|Baseline|2015-09-15|2015-10-20|Complete|Done|4|1|4|4|4|4|3.5|||||||||3|3|4|4|4|3|3.5|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow||Volunteer: Moved|12.9||1|1|1|1|M|Black||12|No|Mother|28273|7|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||RTBM|M|Black||29|28273|High School Graduate|Married|Military|28078|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|504290756|504292957|31|0|1|504315689|31|0|1|500844152|2||-2||4|2|||-2||-2|0|10|||46|2|||1|934222|-1|4|3|44|2763237020791144915
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-10-20|2016-11-17|Followup|2016-10-20|2016-10-27|Complete|Done|4|4|4|4|4|4|4|4|1|4|4|4|4|3.5|14.29|2|4|4|4|4|4|3.67|3|3|4|4|4|3|3.5|4.86|4|4|4|4|4|4|4|4|0|4|5|4|5|4.5|5|4|3|4|4|12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3|3.71|7.82|4|4|4|4|4|4|4|4|0|3|2|2.5|4|4|4|-37.5|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Moved|12.9||1|1|1|1|M|Black||12|No|Mother|28273|7|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||RTBM|M|Black||29|28273|High School Graduate|Married|Military|28078|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|504290756|504292957|31|0|1|504315689|31|0|1|500844152|2||-2||4|2|||-2||-2|0|10|||46|2|||1|947550|934222|4|3|45|2763237020791144915
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-10-21|2016-03-04|Baseline|2015-10-01|2015-10-21|Complete|Done|2|4|4|4|4|4|3.67|||||||||1|4|2|2|2|3|2.33|||||||||4|4|4|4||||||2|3|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||1|1||||4|4||||Green|PERL 2014-2016|Child/Family: Moved|4.4||1|1|2|2|M|Black||14|No|Mother|28212|5|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|Amachi, PERL 2014-2016|Enrollment|M|White||30|28209|Bachelors Degree|Married|Real Estate: Realtor|28217|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|503863366|503865360|31|0|1|504322037|1|0|1|500843765|2||-2||4|1|500014681|500000294, 500014681|-2||-2|0|5|||46|2|||1|939888|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-23|NaT|Followup|2016-10-23|2016-10-25|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|2|3|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||16.5||3|3|1|1|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28083|2|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|M|White||39|28027|Masters Degree|Married|Business|28269|9|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|502234905|502777258|38|0|1|504334608|1|0|1|500843097|2||500016307||2|1|500014681, 500016374|500000294, 500014681, 500016374|-2|500014681, 500016374|-2|0|10|||17159|12|||1|949913||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-28|NaT|Followup|2016-10-28|2016-10-20|Complete|Done|4|2|2|1|4|4|2.83|||||||||2|4|4|2|1|4|2.83|||||||||3|4|4|3.67||||||5|5|5|5|5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|Cabarrus County||16.3||1|1|2|2|M|Black||9|No|Mother|28027|4|One Parent: Female|$75,000 to $99,999||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|Black||34|28269|Some College|Married|Business|28025|5|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County, mentor2.0 2014|Match Support|277|60|598|500000170|500022817|503911799|503913806|31|0|1|503956879|31|0|1|500849358|2||500016307||2|2|500016374|500016374|-2|500014506, 500016374|-2|34|2|||7671|13|||1|1001945||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-29|NaT|Followup|2016-10-29|2016-10-10|Complete|Early|3|4|4|2|3|3|3.17|||||||||2|4|3|3|2|4|3|||||||||4|4|4|4||||||2|5|5|4|4|||||||3|4|4|4|4|4|3|3.71||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||16.3||4|4|1|1|F|White||18|No|Father|28025||One Parent: Male|Unknown||No||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||68|28027|Associate Degree|Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|500341548|500341682|1|0|2|504323327|1|0|2|500844725|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|3|||17159|12|||1|953186||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Baseline|2015-09-21|2015-10-30|Complete|Done|4|1|4|2|3|4|3|||||||||1|3|3|2|2|3|2.33|||||||||4|4|4|4||||||1|1|2|2|1.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|||16.2||1|1|1|1|F|Black||10|No|Mother|28216|4|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|F|Black||31|28216|Bachelors Degree|Single|Arts, Entertainment, Sports|28202|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504345626|504347850|31|0|2|504373316|31|0|2|500845709|2||-2||2|1|||-2||-2|0|10|||46|2|||1|935912|-1|4|3|44|1712849328738258411
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Baseline|2015-10-08|2015-10-30|Complete|Done|2|4|3|2|4|3|3|||||||||2|3|4|4|3|3|3.17|||||||||3|4|3|3.33||||||4|5|2|3|3.5|||||||4|3|2|2|3|4|4|3.14||||||||||3|4|2|3||||||3|3|3|||||2|2||||4|4||||Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016||16.2|Y|1|1|1|1|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28204|Masters Degree|Married|Consultant||0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504254978|504257111|3|0|1|504379733|1|0|1|500845639|2||-2||2|1|500011312, 500014681|500014681|-2|500014681|-2|0|5|||46|2|||1|942403|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Followup|2016-10-30|2016-12-14|Complete|Done|3|2|4|2|3|3|2.83|4|1|4|2|3|4|3|-5.67|2|3|2|2|3|3|2.5|1|3|3|2|2|3|2.33|7.3|4|4|4|4|4|4|4|4|0|2|2|3|2|2.25|1|1|2|2|1.5|50|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|2|2|3|1|2|0|2|2|2|2|0|4|4|4|4|0|Green|||16.2||1|1|1|1|F|Black||10|No|Mother|28216|4|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|F|Black||31|28216|Bachelors Degree|Single|Arts, Entertainment, Sports|28202|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504345626|504347850|31|0|2|504373316|31|0|2|500845709|2||-2||2|1|||-2||-2|0|10|||46|2|||1|953778|935912|4|3|45|1712849328738258411
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Followup|2016-10-30|2016-10-27|Complete|Done|2|2|2|2|3|4|2.5|2|4|3|2|4|3|3|-16.67|4|2|3|2|2|3|2.67|2|3|4|4|3|3|3.17|-15.77|4|4|4|4|3|4|3|3.33|20.12|3|2|3|3|2.75|4|5|2|3|3.5|-21.43|4|4|4|4|4|4|3|3.86|4|3|2|2|3|4|4|3.14|22.93|4|4|3|3.67|3|4|2|3|22.33|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016||16.2|Y|1|1|1|1|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28204|Masters Degree|Married|Consultant||0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504254978|504257111|3|0|1|504379733|1|0|1|500845639|2||-2||2|1|500011312, 500014681|500014681|-2|500014681|-2|0|5|||46|2|||1|953996|942403|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-04|NaT|Baseline|2015-10-27|2015-11-04|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||16.1||1|1|1|1|F|Multi-race (Hispanic & Asian)||10|No|Mother|28081|5|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||40|28025||Married|Self-Employed, Entrepreneur||11|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504432726|504434981|40|0|2|504430061|1|0|2|500852606|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7464|9|||1|951286|-1|4|3|44|3993797463174785246
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-04|NaT|Followup|2016-11-04|2016-10-31|Complete|Done|3|4|4|2|4|4|3.5|4|4|4|4|4|4|4|-12.5|2|4|4|2|3|4|3.17|4|4|4|1|4|4|3.5|-9.43|4|4|4|4|4|4|4|4|0|4|4|4|4|4|5|4|5|5|4.75|-15.79|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|2|3.71|4.04|4|4|4|4|4|4|4|4|0|4|4|4|4|2|3|33.33|1|1|2|2|-50|4|4|4|4|0|Green|PERL 2014-2016, Cabarrus County||16.1||1|1|1|1|F|Multi-race (Hispanic & Asian)||10|No|Mother|28081|5|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||40|28025||Married|Self-Employed, Entrepreneur||11|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504432726|504434981|40|0|2|504430061|1|0|2|500852606|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7464|9|||1|956252|951286|4|3|45|3993797463174785246
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-11|NaT|Baseline|2015-10-13|2015-11-11|Complete|Done|4|1|4|1|3|4|2.83|||||||||2|3|4|4|3|4|3.33|||||||||4|4|4|4||||||1|1|1|1|1|||||||4|4|4|3|1|4|3|3.29||||||||||4|3|1|2.67||||||4|1|2.5|||||1|1||||4|4||||Green|||15.8||1|1|1|1|M|Black||10|Yes|Mother|28216|5|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community|Amachi|Match Support|M|Black||41|28214|Some College|Married|Business|28287|0|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504207638|504209750|31|0|1|504357457|31|0|1|500850393|2||-2||2|1||500000294|-2||-2|0|4|||17159|12|||1|944553|-1|4|3|44|7674215580094440446
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-11|NaT|Followup|2016-11-11|2017-01-26|Expired|Late||||||||4|1|4|1|3|4|2.83|||||||||2|3|4|4|3|4|3.33||||||4|4|4|4|||||||1|1|1|1|1||||||||||4|4|4|3|1|4|3|3.29||||||4|3|1|2.67|||||4|1|2.5||||1|1||||4|4||Green|||15.8||1|1|1|1|M|Black||10|Yes|Mother|28216|5|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community|Amachi|Match Support|M|Black||41|28214|Some College|Married|Business|28287|0|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504207638|504209750|31|0|1|504357457|31|0|1|500850393|2||-2||2|1||500000294|-2||-2|0|4|||17159|12|||1|959794|944553|4|0|45|7674215580094440446
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-11|NaT|Followup|2016-11-11|2016-11-22|Complete|Done|4|2|3|2||4||||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|2|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016||15.8||1|1|1|1|F|Black||10|No|Mother|28216|3|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Hispanic||26|28031|Bachelors Degree|Single|Tech: Research/Design|28117|0|8|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504390954|504393193|31|0|2|504231700|3|0|2|500853984|2||-2||2|1|500014681||-2||-2|0|10|||17159|12|||1|962340||4|3|45|3650724132819756420
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-11-13|2017-02-27|Baseline|2015-10-14|2015-11-13|Complete|Done|3|4|4|1|1|3|2.67|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||4|2|5|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|3|2|3||||||4|4|4|||||1|1||||4|4||||Green||Volunteer: Time constraint|15.5||1|1|1|1|F|Black||16|No|Mother|28216|9|Two Parent|Unknown||Yes||School|General Community||Match Support|F|White||31|28203|Bachelors Degree|Married|Business: Mgt, Admin|28255|0|9|Other|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500018851|504269922|504272121|31|0|2|504285435|1|0|2|500847702|2||-2||4|1|||-2||-2|0|4|||18267|3|||1|944945|-1|4|3|44|3260639349613832803
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-11-13|2017-02-27|Followup|2016-11-13|2016-11-22|Complete|Done|3|2|1|2|1|1|1.67|3|4|4|1|1|3|2.67|-37.45|2|4|4|2|2|4|3|4|4|4|4|2|4|3.67|-18.26|4|4|4|4|4|4|4|4|0|4|3|5|5|4.25|4|2|5|3|3.5|21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|2|2|2.33|4|3|2|3|-22.33|4|3|3.5|4|4|4|-12.5|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Time constraint|15.5||1|1|1|1|F|Black||16|No|Mother|28216|9|Two Parent|Unknown||Yes||School|General Community||Match Support|F|White||31|28203|Bachelors Degree|Married|Business: Mgt, Admin|28255|0|9|Other|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500018851|504269922|504272121|31|0|2|504285435|1|0|2|500847702|2||-2||4|1|||-2||-2|0|4|||18267|3|||1|961096|944945|4|3|45|3260639349613832803
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-16|NaT|Followup|2016-11-16|2016-11-30|Complete|Done|3|3|3|2|3|3|2.83|4|4|4|1|4|4|3.5|-19.14|3|4|4|4|4|4|3.83|4|4|3|1|2|4|3|27.67|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|5|5|4.25|-5.88|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|4|4|3|4|4|3.67|8.99|4|4|4|3|1|2|100|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||15.7||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28216|Bachelors Degree|Married|Business|28202|0|10|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504378557|1|0|1|500856483|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|961771|905704|4|3|45|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Baseline|2015-11-10|2015-11-17|Complete|Done|3|1|1|1|3|1|1.67|||||||||1|1|2|1|1|4|1.67|||||||||4|4|4|4||||||2|5|1|1|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016, Cabarrus County||15.6||1|1|1|1|M|White||15|Yes|Mother|28025|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28025|High School Graduate|Single|Business: Sales|28025|5|0|Local TV|Media|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821678|503823656|1|0|1|504468148|1|0|1|500858177|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7438|1|||1|959176|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Baseline|2015-11-10|2015-11-17|Complete|Done|3|1|1|1|1|1|1.33|||||||||1|3|4|2|1|4|2.5|||||||||1|1|1|1||||||4|3|5|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|2|4|3||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016, Cabarrus County||15.6||1|1|1|1|M|White||12|Yes|Mother|28025|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||32|28025|Bachelors Degree||Business: Sales||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821686|503823656|1|0|1|504460050|1|0|1|500858397|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7496|10|||1|959399|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Followup|2016-11-17|2016-11-14|Complete|Done|4|4|1|1|1|4|2.5|3|1|1|1|3|1|1.67|49.7|4|4|4|4|4|4|4|1|1|2|1|1|4|1.67|139.52|2|4|4|3.33|4|4|4|4|-16.75|5|4|4|5|4.5|2|5|1|1|2.25|100|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|2|3.33|4|4|3|3.67|-9.26|2|4|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016, Cabarrus County||15.6||1|1|1|1|M|White||15|Yes|Mother|28025|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28025|High School Graduate|Single|Business: Sales|28025|5|0|Local TV|Media|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821678|503823656|1|0|1|504468148|1|0|1|500858177|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7438|1|||1|962415|959176|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Followup|2016-11-17|2016-11-14|Complete|Done|1|1|4|1|1|4|2|3|1|1|1|1|1|1.33|50.38|2|2|4|2|2|4|2.67|1|3|4|2|1|4|2.5|6.8|2|2|4|2.67|1|1|1|1|167|5|4|5|5|4.75|4|3|5|2|3.5|35.71|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|4|3.67|3|2|4|3|22.33|3|2|2.5|4|4|4|-37.5|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016, Cabarrus County||15.6||1|1|1|1|M|White||12|Yes|Mother|28025|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||32|28025|Bachelors Degree||Business: Sales||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821686|503823656|1|0|1|504460050|1|0|1|500858397|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7496|10|||1|962429|959399|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-18|NaT|Followup|2016-11-18|2016-11-21|Complete|Done|4|2|1|1|1|2|1.83|4|2|4|1|4|2|2.83|-35.34|4|4|4|4|3|4|3.83|4|4|3|1|4|4|3.33|15.02|4|4|4|4|4|4|4|4|0|4|5|5|2|4|5|4|4|5|4.5|-11.11|4|4|4|4|4|4|2|3.71|4|4|4|4|4|4|3|3.86|-3.89|4|3|4|3.67|4|2|4|3.33|10.21|2|1|1.5|4|4|4|-62.5|2|2|1|1|100|4|4|4|4|0|Green|Cabarrus County||15.6||2|2|1|1|M|White||12|No|Mother|28025|4|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||56|28269|Doctor of Medicine (MD)|Married|Medical: Doctor, Provider|28025|28|0|Agency Sponsored|Special Event|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503532014|503533889|1|0|1|504408440|1|0|1|500853427|2||500016307||2|1|500016374|500000294, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||16426|8|||1|963330|717073|4|3|45|1786514887916898235
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-11-19|2016-10-10|Baseline|2015-11-03|2015-11-19|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|2|3|2|1|3|2.17|||||||||2|2|2|2||||||1|3|1|1|1.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016|Volunteer: Moved|10.7||1|1|1|1|M|White||14|No|Mother|28209|7|One Parent: Female|$20,000 to $24,999||No||Self|General Community|PERL 2014-2016|Enrollment|M|White||27|28278|Masters Degree|Married|Business: Engineer|28278|2|8|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch Training Final Assessment|Match Support|277|60|598|500000170|500018851|504298668|504300882|1|0|1|504372921|1|0|1|500855505|2||-2||4|1|500014681|500014681|-2|500011316|-2|0|10|||17159|12|||1|955691|-1|4|3|44|2656293275676608966
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-19|NaT|Followup|2016-11-19|2017-01-17|Complete|Late|3|4|4|4|3|3|3.5|4|4|4|3|3|3|3.5|0|3|4|4|3|2|4|3.33|4|1|3|3|3|4|3|11|4|4|4|4|4|4|4|4|0|3|4|5|5|4.25|5|5|5|5|5|-15|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green|mentor2.0, mentor2.0 2014, mentor2.0 2015||15.6||1|2|1|2|M|Black||16|Yes|Mother|28208|9|One Parent: Female|Unknown|Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|M|White||26|28210|Bachelors Degree||Business|28281|0|5|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|277|60|598|500000170|500022907|504043128|504045146|31|0|1|503985272|1|0|1|500861533|2||500015511||2|1|500014505, 500014506, 500015184|500014505, 500014506|-2|500014506|-2|0|4|||7462|13|||1|963994|800113|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-11-23|2017-01-17|Baseline|2015-07-24|2015-11-23|Complete|Done|3|1|2|2|2|2|2|||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||2|5|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016|Volunteer: Lost contact with child/agency|13.8||1|1|1|1|M|Black||12|No|GrandMother|28215|6|Grandparents|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI, PERL 2014-2016|Enrollment|M|Black||30|28262|Some College|Married|Architect|28207|0|6|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment|Match Support|277|60|598|500000170|500021785|502458458|502458905|31|0|1|504387453|31|0|1|500855881|2||-2||4|1|500014681|500005291, 500014681|-2|500011316, 500014681|-2|0|5|||46|2|||1|918544|-1|4|3|44|3274057295643004474
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-23|NaT|Baseline|2015-11-06|2015-11-23|Complete|Done|3|4|1|4|4|4|3.33|||||||||2|4|3|1|2|3|2.5|||||||||3|4|4|3.67||||||3|4|2|2|2.75|||||||4|4|4|4|4|4|2|3.71||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016||15.4||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28208|3|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||30|28204|Some College|Single|Medical|28208|3|3|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504278828|504281028|38|0|2|504354967|35|0|2|500857068|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|957729|-1|4|3|44|2378213070582218846
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-23|NaT|Followup|2016-11-23|2016-11-25|Complete|Done|4|4|4|4|4|4|4|3|4|1|4|4|4|3.33|20.12|2|4|4|3|3|4|3.33|2|4|3|1|2|3|2.5|33.2|4|4|4|4|3|4|4|3.67|8.99|4|3|3|4|3.5|3|4|2|2|2.75|27.27|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|2|3.71|4.04|4|4|4|4|3|3|3|3|33.33|4|3|3.5|4|4|4|-12.5|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||15.4||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28208|3|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||30|28204|Some College|Single|Medical|28208|3|3|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504278828|504281028|38|0|2|504354967|35|0|2|500857068|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|965373|957729|4|3|45|2378213070582218846
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-24|NaT|Baseline|2015-09-22|2015-11-24|Complete|Done|4|3|4|4|3|4|3.67|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|2|4|3|3.57||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||15.4||1|1|1|1|M|Black||12|No|Mother|28211|5|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||48|28105||Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504227502|504229617|31|0|1|504460839|31|0|1|500859784|2||-2||2|1||500000294|-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1|936163|-1|4|3|44|2077565980961547475
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-24|NaT|Followup|2016-11-24|2016-12-27|Declined|Done||||||||4|3|4|4|3|4|3.67|||||||||2|4|4|2|3|4|3.17||||||4|4|4|4|||||||3|3|3|4|3.25||||||||||4|4|4|4|2|4|3|3.57||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Green|||15.4||1|1|1|1|M|Black||12|No|Mother|28211|5|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||48|28105||Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504227502|504229617|31|0|1|504460839|31|0|1|500859784|2||-2||2|1||500000294|-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1|966066|936163|4|1|45|2077565980961547475
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-30|NaT|Baseline|2015-11-17|2015-11-30|Complete|Done|2|2|1|2|2|3|2|||||||||2|3|3|2|3|4|2.83|||||||||2|3|2|2.33||||||4|4|5|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|VOL - Mentoring Hispanic Youth, PERL 2014-2016||15.2||1|1|2|2|F|Hispanic||13|No|Mother|28205|6|Two Parent|Unknown||Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504331538|504333760|3|0|2|503843020|3|0|2|500860738|2||-2||2|2|500011312, 500014681|500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|962816|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-30|NaT|Followup|2016-11-30|2016-11-29|Complete|Done|2|4|4|4|1|1|2.67|2|2|1|2|2|3|2|33.5|2|4|3|2|4|3|3|2|3|3|2|3|4|2.83|6.01|4|4|4|4|2|3|2|2.33|71.67|5|3|3|4|3.75|4|4|5|3|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|4|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Yellow|VOL - Mentoring Hispanic Youth, PERL 2014-2016||15.2||1|1|2|2|F|Hispanic||13|No|Mother|28205|6|Two Parent|Unknown||Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504331538|504333760|3|0|2|503843020|3|0|2|500860738|2||-2||2|2|500011312, 500014681|500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|967639|962816|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-02|NaT|Followup|2016-12-02|2016-12-10|Complete|Done|1|1|4|4|4|1|2.5|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||2|5|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||15.1||2|2|4|4|F|Black||17|Yes|GrandMother|28273|10|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501300013|500561354|31|0|2|500346193|31|0|2|500864495|2||-2||2|1||500000294|-2||-2|7294|13|||46|2|||1|968911||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-07|2016-05-24|Baseline|2015-11-06|2015-12-07|Complete|Done|3|4|2|2|3|4|3|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||2|3|4|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|5.6||1|1|1|1|M|Black||14|No|Mother|28027|7|One Parent: Female|$25,000 to $29,999||Yes||School|General Community||Match Support|M|White||24|28262||Single|Medical: Healthcare Worker|28025|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|502129820|502130249|31|0|1|504474407|1|0|1|500858150|2||-2||4|3|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|957862|-1|4|3|44|2881622112345502539
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-07|2017-01-12|Baseline|2015-11-20|2015-12-07|Complete|Done|1|1|4|1|1|2|1.67|||||||||3|2|2|2|3|2|2.33|||||||||4|4|4|4||||||5|3|1|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||1|1||||4|4||||Red|PERL 2014-2016, Cabarrus County|Volunteer: Lost contact with child/agency|13.2||2|2|1|1|M|Multi-race (Black & White)||13|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||No||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|Black||26|28262|Bachelors Degree|Single|Business: Sales|28025|0|1|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|504517520|504519821|36|0|1|504355611|31|0|1|500862169|2||500016307||4|3|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||17159|12|||1|964977|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-07|2017-01-12|Followup|2016-12-07|2016-12-18|Complete|Done|2|2|1|1|2|1|1.5|1|1|4|1|1|2|1.67|-10.18|1|4|2|2|3|2|2.33|3|2|2|2|3|2|2.33|0|4|4|4|4|4|4|4|4|0|5|4|2|2|3.25|5|3|1|3|3|8.33|4|4|4|4|2|4|4|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|2|3.33|4|4|4|4|-16.75|2|2|2|2|4|3|-33.33|1|1|1|1|0|4|4|4|4|0|Red|PERL 2014-2016, Cabarrus County|Volunteer: Lost contact with child/agency|13.2||2|2|1|1|M|Multi-race (Black & White)||13|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||No||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|Black||26|28262|Bachelors Degree|Single|Business: Sales|28025|0|1|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|504517520|504519821|36|0|1|504355611|31|0|1|500862169|2||500016307||4|3|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||17159|12|||1|970571|964977|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-08|NaT|Followup|2016-12-08|2017-02-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||14.9||1|1|1|1|M|Black||10|No|Mother|28208|2|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community||Match Support|M|White||27|28203|Bachelors Degree|Single|Insurance|21202|2|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504046908|504048929|31|0|1|504349113|1|0|1|500863535|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|56|1|||17159|12|||1|994081||4|0|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-14|2016-05-19|Baseline|2015-11-17|2015-12-14|Complete|Done|3|4|4|4|3|2|3.33|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|2|3|2.67||||||2|3|2.5||||||||||3|3||||Green|PERL 2014-2016|Volunteer: Moved|5.2||1|1|1|1|F|Black||16|No|Mother|28215|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||25|28205|Bachelors Degree|Single|Business|28031|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017777|503611723|503613600|31|0|2|504295160|1|0|2|500860670|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|10|||17159|12|||1|962728|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-14|NaT|Baseline|2015-11-20|2015-12-14|Complete|Done|3|3|2|1|2|3|2.33|||||||||2|3|3|3|2|4|2.83|||||||||4|4|3|3.67||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||2|3|1|2||||||4|3|3.5|||||2|2||||4|4||||Green|Amachi, PERL 2014-2016||14.8||1|1|1|1|F|Black||15|Yes|Mother|28215|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi, PERL 2014-2016|Match Support|F|White||30|28203|Bachelors Degree|Single|Business|60611|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|503611732|503613600|31|0|2|504421910|1|0|2|500862006|2||-2||2|1|500000294, 500014681|500000294, 500014681|-2|500014681|-2|0|10|||17159|12|||1|964751|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-14|NaT|Followup|2016-12-14|2016-12-12|Complete|Done|4|4|3|3|3|3|3.33|3|3|2|1|2|3|2.33|42.92|2|4|3|1|2|4|2.67|2|3|3|3|2|4|2.83|-5.65|4|2|2|2.67|4|4|3|3.67|-27.25|4|4|5|2|3.75|4|4|4|5|4.25|-11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|2|2.67|2|3|1|2|33.5|2|2|2|4|3|3.5|-42.86|2|2|2|2|0|4|4|4|4|0|Green|Amachi, PERL 2014-2016||14.8||1|1|1|1|F|Black||15|Yes|Mother|28215|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi, PERL 2014-2016|Match Support|F|White||30|28203|Bachelors Degree|Single|Business|60611|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|503611732|503613600|31|0|2|504421910|1|0|2|500862006|2||-2||2|1|500000294, 500014681|500000294, 500014681|-2|500014681|-2|0|10|||17159|12|||1|973924|964751|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-15|2017-02-28|Baseline|2015-11-30|2015-12-15|Complete|Done|4|1|4|1|4|4|3|||||||||1|1|4|4|1|4|2.5|||||||||4|4|4|4||||||1|4|3|4|3|||||||4|4|3|4|4|3|4|3.71||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Time constraint|14.5||1|1|1|1|M|Black||15||Mother|28209|8|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||31|28207|Masters Degree|Married|Finance: Accountant|28202|7|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504289347|504291548|31|0|1|504428167|1|0|1|500863609|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|967613|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-15|2017-02-28|Followup|2016-12-15|2016-12-01|Complete|Done|3|4|4|2|3|4|3.33|4|1|4|1|4|4|3|11|3|2|3|3|2|3|2.67|1|1|4|4|1|4|2.5|6.8|4|4|4|4|4|4|4|4|0|5|4|5|4|4.5|1|4|3|4|3|50|4|4|4|4|4|4|4|4|4|4|3|4|4|3|4|3.71|7.82|4|4|3|3.67|4|4|4|4|-8.25|4|4|4|3|4|3.5|14.29|1|1|2|2|-50|4|4|4|4|0|Red|PERL 2014-2016|Volunteer: Time constraint|14.5||1|1|1|1|M|Black||15||Mother|28209|8|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||31|28207|Masters Degree|Married|Finance: Accountant|28202|7|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504289347|504291548|31|0|1|504428167|1|0|1|500863609|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|974202|967613|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-15|NaT|Baseline|2015-11-30|2015-12-15|Complete|Done|2|2|2|3|3|2|2.33|||||||||4|2|4|4|4|4|3.67|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||1|1||||4|4||||Green|PERL 2014-2016||14.7||1|1|1|1|F|Black||15|No|Mother|28215|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||26|28213|Bachelors Degree|Single|Business: Mgt, Admin|28105|2|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500021785|504393421|504395660|31|0|2|504395484|31|0|2|500863556|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||46|2|||1|967546|-1|4|3|44|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-15|NaT|Followup|2016-12-15|2017-03-01|Expired|Late||||||||2|2|2|3|3|2|2.33|||||||||4|2|4|4|4|4|3.67||||||4|4|4|4|||||||4|3|3|3|3.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||2|2|2||||1|1||||4|4||Green|PERL 2014-2016||14.7||1|1|1|1|F|Black||15|No|Mother|28215|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||26|28213|Bachelors Degree|Single|Business: Mgt, Admin|28105|2|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500021785|504393421|504395660|31|0|2|504395484|31|0|2|500863556|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||46|2|||1|974242|967546|4|0|45|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-17|2016-08-29|Baseline|2015-12-07|2015-12-17|Complete|Done|4|2|4|2|4|4|3.33|||||||||2|4|2|2|2|2|2.33|||||||||4|3|3|3.33||||||3|4|2|4|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment, PERL 2014-2016|Volunteer: Lost contact with child/agency|8.4||1|1|1|1|M|Black||14|No|Mother|28269|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||RTBM|M|Black||40|28269|Bachelors Degree|Married|Tech: Support, Writing|28269|4|0|Local Radio|Media|Big|General Community|Amachi, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|504245120|504247236|31|0|1|504396885|31|0|1|500865817|2||-2||4|1|500007920, 500011315, 500011316, 500014681||-2|500000294, 500007920, 500011315, 500011316, 500014681|-2|0|4|||7437|1|||1|970842|-1|4|3|44|1546374315672654438
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2015-12-18|2016-01-08|Baseline|2015-12-08|2015-12-17|Complete|Done|3|3|3|3|4|4|3.33|||||||||2|4|3|3|4|4|3.33|||||||||4|4|4|4||||||2|4|3|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|0.7||1|1|1|1|F|Black||15|No|Mother|28269|8|One Parent: Female|$30,000 to $34,999||Yes||School|General Community|VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|F|White||26|28078|Masters Degree|Single|Business: Marketing|28269|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|277|60|598|500000170|500017777|504458036|504460294|31|0|2|504416792|1|0|2|500866388|2||-2||4|2||500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|971455|-1|4|3|44|3086452374500817499
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-22|NaT|Baseline|2015-12-04|2015-12-22|Complete|Done|3|2|2|2|3|4|2.67|||||||||2|3|3|3|4|3|3|||||||||3|3|3|3||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|2|2.5|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||14.5||1|1|2|2|M|White||12|No|Mother|28027|5|One Parent: Female|$30,000 to $34,999||Yes||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||58|28075|Masters Degree|Married|Business|32824|0|6|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504530586|504532918|1|0|1|503694720|1|0|1|500865400|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|3|||7464|9|||1|970132|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-22|NaT|Followup|2016-12-22|2017-01-12|Complete|Done|3|2|3|2|3|4|2.83|3|2|2|2|3|4|2.67|5.99|2|3|2|2|2|2|2.17|2|3|3|3|4|3|3|-27.67|3|3|3|3|3|3|3|3|0|3|4|3|4|3.5|3|3|4|3|3.25|7.69|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|3|3|3|3|3|3|0|3|3|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016, Cabarrus County||14.5||1|1|2|2|M|White||12|No|Mother|28027|5|One Parent: Female|$30,000 to $34,999||Yes||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||58|28075|Masters Degree|Married|Business|32824|0|6|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504530586|504532918|1|0|1|503694720|1|0|1|500865400|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|3|||7464|9|||1|977131|970132|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-28|NaT|Followup|2016-12-28|2017-02-09|Declined|Done||||||||4|1|3|1|4|4|2.83|||||||||1|4|4|4|4|4|3.5||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||1|1|1||||2|2||||4|4||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||14.3||2|2|1|1|M|Black||13|Yes|Mother|28204||One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community|Amachi|Match Support|M|White||24|28202|Bachelors Degree|Single|Finance: Banking|28202|0|5|Other|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|503663975|503665933|31|0|1|504468271|1|0|1|500868596|2||-2||2|1|500007920, 500011315, 500011316|500000294|-2|500007920, 500011315, 500011316|-2|0|10|||18267|3|||1|978234|736588|4|1|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-01-14|2016-08-29|Baseline|2015-11-09|2016-01-14|Complete|Done|3|3|3|1|2|3|2.5|||||||||2|3|3|4|3|4|3.17|||||||||4|4|4|4||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Green|PERL 2014-2016|Volunteer: Lost contact with child/agency|7.5||1|1|1|1|F|Black||10|No|Mother|28056|4|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||RTBM|F|White||30|28209|Bachelors Degree|Single|Finance: Banking|28211|3|2|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|504407275|504409521|31|0|2|504393547|1|0|2|500857377|2||-2||4|1|500014681||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|958346|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-01-14|NaT|Baseline|2015-11-24|2016-01-14|Complete|Done|1|1|3|3|2|1|1.83|||||||||1|1|4|4|4|4|3|||||||||4|4|4|4||||||2|5|2|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||13.7||1|1|1|1|F|Black||10|No|Mother|28203|3|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||25|28209|Bachelors Degree|Single|Business|28277|1|0|Bowl For Kids Sake|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504388295|504390534|31|0|2|504404378|1|0|2|500870013|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||132|8|||1|966128|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-01-14|NaT|Followup|2017-01-14|2017-02-20|Complete|Done|3|3|3|2|3|3|2.83|1|1|3|3|2|1|1.83|54.64|2|4|3|2|2|3|2.67|1|1|4|4|4|4|3|-11|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|2|5|2|5|3.5|-7.14|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|4|4|4|4|-16.75|2|3|2.5|4|3|3.5|-28.57|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||13.7||1|1|1|1|F|Black||10|No|Mother|28203|3|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||25|28209|Bachelors Degree|Single|Business|28277|1|0|Bowl For Kids Sake|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504388295|504390534|31|0|2|504404378|1|0|2|500870013|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||132|8|||1|982719|966128|4|3|45|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-01-21|2016-08-29|Baseline|2016-01-11|2016-01-21|Complete|Done|3|4|4|1|4|4|3.33|||||||||2|2|3|2|1|2|2|||||||||4|3|3|3.33||||||2|5|3|4|3.5|||||||1|1|2|4|3|3|4|2.57||||||||||2|4|3|3||||||2|4|3|||||1|1||||3|3||||Green|PERL 2014-2016|Volunteer: Feels incompatible with child/family|7.3||1|1|1|1|M|Black||15|No|Mother|28269|7|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Multi-race (Black & White)||27|28115|Bachelors Degree|Single|Business|28115|4|4|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500017777|504268284|504270481|31|0|1|503172653|36|0|1|500871097|2||-2||4|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|981397|-1|4|3|44|2378213070582218846
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-01-21|NaT|Followup|2017-01-21|2017-01-20|Complete|Done|3|4|4|2|3|4|3.33|3|4|4|2|4|4|3.5|-4.86|3|4|4|3|3|4|3.5|2|2|3|3|3|3|2.67|31.09|4|4|4|4|3|2|2|2.33|71.67|3|4|4|3|3.5|4|3|5|4|4|-12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||13.5||2|2|1|1|F|White||13|No|Father|28211|8|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||31|28205|Bachelors Degree|Single|Business: Mgt, Admin|28269|8|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|503405468|503407325|1|0|2|504322859|1|0|2|500870080|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|985022|611443|4|3|45|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-01-30|2017-02-27|Baseline|2015-12-22|2016-01-30|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|2|3|1|2|3|2.17|||||||||4|4|4|4||||||2|5|1|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|2|2.5|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment, PERL 2014-2016|Agency: Challenges with program/partnership|12.9||1|1|2|2|M|Black||15|No|Mother|28269|8|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||32|28202|Masters Degree|Single|Finance: Accountant|28202|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504397554|504399794|31|0|1|504206321|1|0|1|500869278|2||-2||4|1|500007920, 500011315, 500011316, 500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||17159|12|||1|977221|-1|4|3|44|5898021503604846505
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-01-30|2016-05-20|Baseline|2016-01-14|2016-01-30|Complete|Done|4|2|4|4|4|4|3.67|||||||||2|3|3|3|1|3|2.5|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|Volunteer: Moved|3.6||2|2|1|1|F|Black||12|No|Mother|28214|5|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||32|28208|Bachelors Degree|Single|Journalist/Media||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503976557|503978568|31|0|2|504365048|1|0|2|500871811|2||-2||4|1|500007920, 500011315, 500011316||-2||-2|34|2|||7464|9|||1|982536|-1|4|3|44|3198188609986797983
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-01-30|NaT|Baseline|2016-01-22|2016-01-29|Complete|Done|4|1|2|1|4|4|2.67|||||||||1|4|3|1|1|3|2.17|||||||||4|3|4|3.67||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||1|1|1|||||2|2||||4|4||||Green|Cabarrus County||13.2||1|1|1|1|F|Multi-race (Hispanic & White)||10|No|Mother|28025|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||25|28269||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504532725|504535058|35|0|2|503951023|1|0|2|500874940|2||500016307||2|1|500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||7496|10|||1|986043|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-01-30|NaT|Followup|2017-01-30|2017-01-26|Complete|Done|4|1|1|1|2|1|1.67|4|1|2|1|4|4|2.67|-37.45|1|4|4|1|1|3|2.33|1|4|3|1|1|3|2.17|7.37|1|4|4|3|4|3|4|3.67|-18.26|5|3|5|5|4.5|5|5|5|5|5|-10|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3.67|8.99|2|1|1.5|1|1|1|50|2|2|2|2|0|4|4|4|4|0|Green|Cabarrus County||13.2||1|1|1|1|F|Multi-race (Hispanic & White)||10|No|Mother|28025|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||25|28269||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504532725|504535058|35|0|2|503951023|1|0|2|500874940|2||500016307||2|1|500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||7496|10|||1|989056|986043|4|3|45|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-01-31|2016-06-06|Baseline|2016-01-15|2016-01-31|Complete|Done|4|1|4|2|4|4|3.17|||||||||3|2|3|4|4|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||2|2|2|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Feels incompatible with child/family|4.2||1|1|1|1|M|Black||14|No|Mother|28212|6|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Enrollment|M|White||38|28227|Some College|Single|Business: Sales||3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500013781|504076403|504078432|31|0|1|504415946|1|0|1|500872171|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||17159|12|||1|983125|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-02-09|2017-02-13|Baseline|2015-10-21|2016-02-09|Complete|Done|3|3|3|4|3|3|3.17|||||||||3|3|2|3|4|2|2.83|||||||||4|4|4|4||||||4|4|3|5|4|||||||4|4|4|3|3|2|3|3.29||||||||||4|4|3|3.67||||||2|4|3|||||1|1||||4|4||||Red|PERL 2014-2016|Volunteer: Moved|12.2||1|1|1|1|M|White||12|No|Mother|28214|7|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community|PERL 2014-2016|Match Support|M|White||56|28012|Some College|Married|Business: Mgt, Admin|33401|4|7|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|504231267|504233379|1|0|1|504379684|1|0|1|500871125|2||-2||4|3|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|3|||46|2|||1|948332|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-12|NaT|Baseline|2016-01-29|2016-02-11|Complete|Done|3|3|3|1|3|3|2.67|||||||||2|4|4|2|4|3|3.17|||||||||2|4|4|3.33||||||3|3|2|5|3.25|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|4|3.67||||||1|4|2.5|||||1|1||||4|4||||Green|PERL 2014-2016||12.8||1|1|1|1|M|Black||11|Yes|Mother|28215|5|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||29|28262|Some College|Single|Business|28204|0|4|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT, VOL - Thrive - Intro|Match Support|277|60|598|500000170|500020753|504230975|504233090|31|0|1|504284612|31|0|1|500876290|2||-2||2|1|500014681|500000294, 500014681|-2|500008492, 500011315, 500011316, 500014681|-2|0|4|||7462|13|||1|988696|-1|4|3|44|7327400833679234452
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-12|NaT|Followup|2017-02-12|2017-02-02|Complete|Done|3|2|3|3|1|2|2.33|3|3|3|1|3|3|2.67|-12.73|4|3|3|3|1|3|2.83|2|4|4|2|4|3|3.17|-10.73|4|4|4|4|2|4|4|3.33|20.12|4|3|5|4|4|3|3|2|5|3.25|23.08|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|2|4|2|2.67|3|4|4|3.67|-27.25|4|4|4|1|4|2.5|60|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||12.8||1|1|1|1|M|Black||11|Yes|Mother|28215|5|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||29|28262|Some College|Single|Business|28204|0|4|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT, VOL - Thrive - Intro|Match Support|277|60|598|500000170|500020753|504230975|504233090|31|0|1|504284612|31|0|1|500876290|2||-2||2|1|500014681|500000294, 500014681|-2|500008492, 500011315, 500011316, 500014681|-2|0|4|||7462|13|||1|993665|988696|4|3|45|7327400833679234452
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-13|NaT|Baseline|2016-02-01|2016-02-13|Complete|Done|4|1|1|3|4|2|2.5|||||||||2|2|3|1|1|4|2.17|||||||||3|4|3|3.33||||||3|5|2|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Cabarrus County||12.7||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28025|3|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||28|28027|Masters Degree|Single|Govt|28273|3|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504468562|504470835|36|0|1|504556956|31|0|1|500876668|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|989695|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-13|NaT|Followup|2017-02-13|2017-02-28|Complete|Done|3|1|3|2|1|3|2.17|4|1|1|3|4|2|2.5|-13.2|3|4|3|2|4|3|3.17|2|2|3|1|1|4|2.17|46.08|4|4|4|4|3|4|3|3.33|20.12|4|3|5|2|3.5|3|5|2|5|3.75|-6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|4|3.5|3|3|3|16.67|2|2|2|2|0|4|4|4|4|0|Green|Cabarrus County||12.7||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28025|3|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||28|28027|Masters Degree|Single|Govt|28273|3|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504468562|504470835|36|0|1|504556956|31|0|1|500876668|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|994031|989695|4|3|45|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-19|NaT|Baseline|2016-02-02|2016-02-19|Complete|Done|3|3|4|3|4|4|3.5|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||3|2|2.5|||||2|2||||4|4||||Red|PERL 2014-2016, Cabarrus County||12.6||1|1|2|2|F|Black||12|No|Mother|28083|5|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||41|28025|Some College|Single|Business|28217|4|0|LPL Financial|Workplace Partner|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504540553|504805582|31|0|2|503680923|31|0|2|500877015|2||500016307||2|3|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||11247|3|||1|990132|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-19|NaT|Followup|2017-02-19|2017-03-02|Complete|Done|3|2|3|2|3|4|2.83|3|3|4|3|4|4|3.5|-19.14|2|3|3|2|3|3|2.67|2|4|3|3|3|3|3|-11|4|4|4|4|4|4|4|4|0|3|3|3|3|3|4|3|4|3|3.5|-14.29|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|3|4|2|3|33.33|4|4|4|3|2|2.5|60|2|2|2|2|0|4|4|4|4|0|Red|PERL 2014-2016, Cabarrus County||12.6||1|1|2|2|F|Black||12|No|Mother|28083|5|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||41|28025|Some College|Single|Business|28217|4|0|LPL Financial|Workplace Partner|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504540553|504805582|31|0|2|503680923|31|0|2|500877015|2||500016307||2|3|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||11247|3|||1|995916|990132|4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-20|NaT|Baseline|2016-02-16|2016-02-20|Complete|Done|3|3|4|3|2|3|3|||||||||4|4|4|3|4|3|3.67|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|3|4|4|2|3.57||||||||||4|4|2|3.33||||||4|4|4|||||2|2||||4|4||||Green|Cabarrus County||12.5||1|1|2|2|M|Multi-race (Asian & White)||14|No|Mother|28027|9|One Parent: Female|$60,000 to $74,999|Y|No||Self|General Community|Cabarrus County|Match Support|M|Black||30|28213|Masters Degree|Single|Education|28217|0|7|Recruitment Event|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504545166|504547500|37|0|1|503788318|31|0|1|500879416|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7458|9|||1|994473|-1|4|3|44|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-20|NaT|Followup|2017-02-20|2017-02-20|Complete|Done|1|4|4|4|3|4|3.33|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||2|4|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||12.5||4|4|1|1|F|Hispanic||12|No|Mother|28027|4|Other/Unknown|Unknown||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||28|28075|Bachelors Degree|Single|Education: Teacher|28025|2|6|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|503270485|503272299|3|0|2|504574450|1|0|2|500880422|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||46|2|||1|996302||4|3|45|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-20|NaT|Followup|2017-02-20|2017-02-17|Complete|Done|3|3|4|4|3|3|3.33|3|3|4|3|2|3|3|11|2|4|2|1|3|2|2.33|4|4|4|3|4|3|3.67|-36.51|4|4|4|4|4|4|4|4|0|2|3|3|5|3.25|4|3|5|5|4.25|-23.53|4|3|4|4|4|3|3|3.57|4|4|4|3|4|4|2|3.57|0|1|2|3|2|4|4|2|3.33|-39.94|2|4|3|4|4|4|-25|1|1|2|2|-50|4|4|4|4|0|Green|Cabarrus County||12.5||1|1|2|2|M|Multi-race (Asian & White)||14|No|Mother|28027|9|One Parent: Female|$60,000 to $74,999|Y|No||Self|General Community|Cabarrus County|Match Support|M|Black||30|28213|Masters Degree|Single|Education|28217|0|7|Recruitment Event|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504545166|504547500|37|0|1|503788318|31|0|1|500879416|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7458|9|||1|996319|994473|4|3|45|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-22|NaT|Baseline|2016-01-14|2016-02-22|Complete|Done|3|2|3|4|3|3|3|||||||||3|2|4|3|3|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||12.5||1|1|1|1|F|Multi-race (Black & White)||10|Yes|Foster Parent|28216|4|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||45|28208|Bachelors Degree|Single|Education: Teacher|28208|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504498650|504500981|36|0|2|504131389|31|0|2|500878445|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1|982537|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-23|NaT|Baseline|2016-02-10|2016-02-23|Complete|Done|4|2|4|1|4|4|3.17|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||12.4||1|1|1|1|M|Black||11|No|Mother|28262|3|One Parent: Female|$30,000 to $34,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504295805|504298006|31|0|1|504337975|1|0|1|500878715|2||-2||2|1|500007920, 500011315, 500011316||-2||-2|34|2|||7464|9|||1|992976|-1|4|3|44|5923747279518652886
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-29|NaT|Baseline|2016-02-18|2016-02-29|Complete|Done|2|1|2|1|2|2|1.67|||||||||3|4|3|2|1|4|2.83|||||||||2|4|2|2.67||||||3|4|2|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|2|3.33||||||2|3|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||12.2||1|1|1|1|M|Black||15|No|Mother|28209|7|One Parent: Female|$25,000 to $29,999||Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||29|28209|Masters Degree|Single|Law: Lawyer|28202|0|4|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|500917189|500917459|31|0|1|504538036|1|0|1|500880191|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||7464|9|||1|995664|-1|4|3|44|2719955880210213907
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-03-10|NaT|Baseline|2015-06-24|2016-03-08|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|PERL 2014-2016||11.9||1|1|1|1|M|Black||13|No|Mother|28208|6|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28202|Bachelors Degree|Single|Law|28202|0|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504237243|504239358|31|0|1|504456306|1|0|1|500881682|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|909217|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-03-14|NaT|Baseline|2016-02-29|2016-03-14|Complete|Done|4|2|2|1|3|3|2.5|||||||||3|4|4|2|2|4|3.17|||||||||4|4|4|4||||||3|4|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green|||11.8||1|1|1|1|F|Black||13|No|Mother|28278|6|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|White||39|28134|Bachelors Degree|Single|Business: Marketing|28204|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504161470|504162947|31|0|2|504396335|1|0|2|500882097|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|999485|-1|4|3|44|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-03-23|NaT|Baseline|2016-03-09|2016-03-23|Complete|Done|4|4|1|2|1|4|2.67|||||||||2|1|3|4|1|3|2.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|Cabarrus County||11.5||1|1|1|1|M|Black||10|No|Mother|28027|3|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||35|28083|High School Graduate|Married|Medical||8|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504563369|504565703|31|0|1|504600175|1|0|1|500883737|2||500016307||2|2|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|1002382|-1|4|3|44|6200244613298520712
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Inactive|2016-03-24|NaT|Baseline|2016-03-14|2016-03-24|Complete|Done|3|4|4|3|3|3|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||11.4||1|1|1|1|F|Black||13|No|Mother|28213|6|One Parent: Female|$15,000 to $19,999|Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||38|28205|Bachelors Degree|Divorced|Business|28209|6|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504399552|504401793|31|0|2|504544485|1|0|2|500884475|2||-2||3|1|||-2|500007920, 500011315, 500011316|-2|0|5|||7464|9|||1|1003680|-1|4|3|44|458259588635328527
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-06|NaT|Baseline|2016-03-30|2016-04-06|Complete|Done|1|4|4|4|4|3|3.33|||||||||2|4|2|2|3|4|2.83|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||11||1|1|1|1|M|Black||12|No|Mother|28208|5|One Parent: Female|$30,000 to $34,999||Yes||Relative|General Community||Match Support|M|White||32|28203|Juris Doctorate (JD)|Single|Law: Lawyer|28277|1|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|503952082|503954090|31|0|1|504546069|1|0|1|500887070|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|0|3|||46|2|||1|1008663|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-19|NaT|Baseline|2016-04-08|2016-04-19|Complete|Done|3|2|3|4|3|3|3|||||||||4|1|4|4|3|4|3.33|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|||10.6||1|1|1|1|M|White||11|No|Mother|28277|4|One Parent: Female|$75,000 to $99,999||No||School|General Community||Match Support|M|White||53|28270|Masters Degree|Married|Self-Employed, Entrepreneur||15|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504581060|504583394|1|0|1|504503934|1|0|1|500888341|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1011466|-1|4|3|44|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Inactive|2016-04-22|NaT|Baseline|2016-04-13|2016-04-22|Complete|Done|3|2|3|2|2|4|2.67|||||||||2|3|4|2|2|3|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||10.5||1|1|2|2|M|Black||13|No|Mother|28269|6|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|M|White||42|28214|Bachelors Degree|Divorced|Business: Engineer||10|0|Self|Self|Big|General Community|Amachi, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504554067|504556401|31|0|1|503373934|1|0|1|500888917|2||-2||3|1|500007920, 500011315, 500011316||-2|500000294, 500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|1012748|-1|4|3|44|1962015587749138391
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-22|NaT|Baseline|2016-03-29|2016-04-19|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|1|4|2|4|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||1|4|2.5|||||2|2||||4|4||||Green|||10.5||1|1|1|1|F|Black||12|No|Mother|28217|4|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||35|28210|Masters Degree|Married|Finance||5|9|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504268884|504271081|31|0|2|504240747|1|0|2|500886770|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1|1008039|-1|4|3|44|20998188998147742
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-24|NaT|Baseline|2016-03-28|2016-04-24|Complete|Done|2|2|2|1|2|3|2|||||||||2|2|3|3|2|3|2.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|Cabarrus County, mentor2.0 2016||10.4||1|1|1|1|F|Black||13|No|Mother|28027|7|Two Parent|$60,000 to $74,999||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||30|28269|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|2|Recruitment Event|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504602680|504605091|31|0|2|504579649|1|0|2|500886605|2||500016307||2|1|500016374, 500016394|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7462|13|||1|1007638|-1|4|3|44|993637920138474088
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-25|NaT|Baseline|2016-04-08|2016-04-25|Complete|Done|4|2|3|2|3|4|3|||||||||3|3|3|3|2|3|2.83|||||||||4|3|4|3.67||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||10.4||1|1|1|1|M|White||11|No|Mother|28277|5|One Parent: Female|$60,000 to $74,999||No||School|General Community||Match Support|M|White||40|28173|Bachelors Degree|Married|Business: Mgt, Admin|33637|9|4|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504240231|504242346|1|0|1|504523981|1|0|1|500888425|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1011564|-1|4|3|44|7406803744350640674
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-28|NaT|Baseline|2016-04-07|2016-04-27|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|3|3|3|2|2|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|3|2.5|||||1|1||||4|4||||Green|PERL 2014-2016, Cabarrus County||10.3||1|1|1|1|M|White||10|No|GrandMother|28124|3|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||35|28027|Bachelors Degree|Single|Tech: Computer/Programmer|28202|2|6|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, mentor2.0, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504640447|504638197|1|0|1|504266263|1|0|1|500888255|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014505, 500016374|-2|0|4|||17159|12|||1|1011251|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-29|NaT|Baseline|2016-04-13|2016-04-26|Complete|Done|4|1|4|2|4|4|3.17|||||||||2|4|3|1|1|4|2.5|||||||||4|2|2|2.67||||||3|2|2|2|2.25|||||||4|3|4|4|4|4|3|3.71||||||||||4|4|4|4||||||3|4|3.5|||||1|1||||4|4||||Green|PERL 2014-2016||10.3||1|1|1|1|M|Black||14|No|Mother|28212|6|One Parent: Female|$35,000 to $39,999||Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|White||35|28215|Some College|Living w/ Significant Other|Tech: Engineer|11735|1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504129013|504131049|31|0|1|504577506|1|0|1|500888874|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|56|1|||7496|10|||1|1012689|-1|4|3|44|2197933814735019388
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-30|NaT|Baseline|2016-04-13|2016-04-30|Complete|Done|3|2||2|3|4||||||||||2|2|3|1|2|3|2.17|||||||||3|4|4|3.67||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|3|3|3.33||||||4|4|4|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||10.2||1|1|1|1|M|Black||15|No|Mother|28120|6|One Parent: Female|Less than $10,000||Yes||Relative|General Community|PERL 2014-2016|Match Support|M|White||28|28214|Bachelors Degree|Married|Business|28214|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|503782093|503784070|31|0|1|504545677|1|0|1|500888935|2||-2||2|1|500007920, 500011315, 500011316|500014681|-2|500007920, 500011315, 500011316|-2|0|3|||17159|12|||1|1012760|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-10|NaT|Baseline|2016-05-02|2016-05-09|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||9.9||1|1|3|3|M|Multi-race (Black & White)||12|Yes|Mother|28215|6|One Parent: Female|$35,000 to $39,999||No||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||57|28269|Bachelors Degree|Married|Finance: Accountant|28202|34|2|Omega Psi Phi|Fraternity/Sorority|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|502183411|502183840|36|0|1|500189229|31|0|1|500891295|2||-2||2|1|500014681|500000294, 500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||8694|14|||1|1019351|-1|4|3|44|4203557099934965158
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-17|NaT|Baseline|2016-04-13|2016-05-17|Complete|Done|3|3|3|4|2|3|3|||||||||3|3|4|2|2|4|3|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||9.7||1|1|1|1|M|Black||13|No|Mother|28213|8|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|Black||27|28215|Bachelors Degree|Single|Tech: Computer/Programmer|28270|2|1|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|503917550|503962680|31|0|1|504577899|31|0|1|500888953|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|1012788|-1|4|3|44|6084148439133243542
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-05-24|2017-02-23|Baseline|2016-05-10|2016-05-24|Complete|Done|2|1|1|2|1|1|1.33|||||||||3|2|3|3|3|2|2.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|2|1|2||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|9||1|1|1|1|M|Black||15|No|Mother|28208|9|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|PHD|Single|Self-Employed, Entrepreneur|30604|4|0|Local Print|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504347348|504349572|31|0|1|504566830|1|0|1|500892524|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|34|2|||7439|1|||1|1022954|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-24|NaT|Baseline|2016-03-15|2016-05-24|Complete|Done|4|3|3|4|3|3|3.33|||||||||4|3|3|4|4|3|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||9.4||1|1|1|1|F|Black||10|No|Mother|28208|4|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||29|28210|Bachelors Degree|Single|Business: Sales|28269|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020910|504556546|504558880|31|0|2|504283498|1|0|2|500889681|2||-2||2|1|500007920, 500011315, 500011316||-2||-2|0|4|||17159|12|||1|1004119|-1|4|3|44|6084148439133243542
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-05-27|2017-01-20|Baseline|2016-05-04|2016-05-27|Complete|Done|3|4|2|4|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|3|4|4|3.86||||||||||3|3|3|3||||||3|2|2.5|||||1|1||||4|4||||Red||Child: Severity of challenges|7.8||1|1|1|1|M|Black||14|No|Mother|28215|7|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|M|White||23|28205|Bachelors Degree|Single|Finance|28210|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500008321|504318423|504320644|31|0|1|504561410|1|0|1|500891770|2||-2||4|3|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1020756|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-05-31|2017-01-27|Baseline|2016-05-02|2016-05-31|Complete|Done|2|3|4|3|3|3|3|||||||||3|3|3|2|3|3|2.83|||||||||4|3|2|3||||||2|3|5|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|3|3|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|Volunteer: Lost contact with child/agency|7.9||1|1|2|2|M|White||14|No|Mother|28214|7|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community||Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|504231264|504233379|1|0|1|504230177|1|0|1|500891315|2||-2||4|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|0|3|||7462|13|||1|1019394|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-31|NaT|Baseline|2016-05-13|2016-05-31|Complete|Done|2|4|4|4|4|2|3.33|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|4|1|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||9.2||1|1|1|1|M|Black||13|No|Mother|28227|7|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|M|Black||27|28205|Some College|Single|Retail: Sales|28210|2|6|Local Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|504425160|504427415|31|0|1|504509415|31|0|1|500893007|2||-2||2|1|||-2||-2|0|4|||7437|1|||1|1024882|-1|4|3|44|5544164653861671456
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-31|NaT|Baseline|2016-05-16|2016-05-31|Complete|Done|2|2|4|2|3|1|2.33|||||||||4|2|2|4|4|4|3.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2||||4|4||||Green|||9.2||1|1|1|1|F|Black||15|No|Mother|28212|8|One Parent: Female|$40,000 to $44,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||48|28212|Associate Degree|Single|Finance||11|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504473782|504476056|31|0|2|504550297|1|0|2|500893115|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1|1025743|-1|4|3|44|2806833304218536184
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-14|NaT|Baseline|2016-06-14|2016-06-14|Complete|Done|3|3|1|2|2|4|2.5|||||||||3|3|4|3|3|3|3.17|||||||||4|3|4|3.67||||||2|5|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Cabarrus County||8.7||1|1|1|1|F|White||11|No|GrandMother|28124|5|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|Cabarrus County|Match Support|F|White||45|28025|Some College||Business|28262|1|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504635786|504638197|1|0|2|504662207|1|0|2|500896660|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|1048528|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-16|NaT|Baseline|2016-05-24|2016-06-16|Complete|Done|4|4|1|4|3|4|3.33|||||||||2|4|3|1|2|3|2.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||8.7||1|1|1|1|F|Black||11|No|Mother|28216|4|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|White||27|28209|Bachelors Degree|Single|Medical|28054|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504628520|504630931|31|0|2|504409458|1|0|2|500894207|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|1031243|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-16|NaT|Baseline|2016-05-27|2016-06-16|Complete|Done|3|3|4|3|3|4|3.33|||||||||1|4|3|3|4|4|3.17|||||||||4|4|4|4||||||2|3|3|4|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||8.7||1|1|1|1|F|Multi-Race (None of the above)||14|No|Mother|28215|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Black||26|28262|Bachelors Degree|Single|Journalist/Media|28206|2|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504507791|504510086|7|0|2|504650231|31|0|2|500895078|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|1034810|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-06-20|2016-11-03|Baseline|2016-05-11|2016-06-20|Complete|Done|2|2|3|2|3|2|2.33|||||||||3|3|3|2|3|4|3|||||||||4|4|4|4||||||5|3|1|3|3|||||||4|4|4|4|3|4|2|3.57||||||||||2|2|1|1.67||||||4|4|4|||||1|1||||3|3||||Green||Volunteer: Lost contact with child/agency|4.5||1|1|1|1|F|Black||14|No|GrandMother|28105|9|Grandparents|$45,000 to $49,999||Yes|BBBS National Site|Web Link|General Community||RTBM|F|Black||39|28105|Bachelors Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504631841|504634252|31|0|2|504167347|31|0|2|500892753|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|1023753|-1|4|3|44|5605796235524810842
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-20|NaT|Baseline|2016-05-23|2016-06-20|Complete|Done|3|2|3|2|2|3|2.5|||||||||3|2|3|4|3|2|2.83|||||||||4|4|4|4||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4||||||||3|3|3|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||8.5||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28213|7|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|Asian||25|28204|Bachelors Degree|Single|Finance|28215|0|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504691840|504694268|36|0|1|504535890|4|0|1|500894068|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1|1030379|-1|4|3|44|8773162532572605235
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-30|NaT|Baseline|2016-01-05|2016-06-30|Complete|Done|4|1|1|1|4|4|2.5|||||||||1|4|3|2|2|3|2.5|||||||||4|4|4|4||||||5|3|3|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|Cabarrus County||8.2||1|1|1|1|M|Multi-race (Hispanic & White)||10|No|Mother|28025|3|One Parent: Female|Unknown|Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28027|Bachelors Degree|Single|Business|28027|2|4|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504553935|504556269|35|0|1|504682974|1|0|1|500897234|2||500016307||2|1|500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|34|2|||7464|9|||1|979891|-1|4|3|44|8216069172157856234
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-30|NaT|Baseline|2016-06-16|2016-06-30|Complete|Done|3|1|1|1|2|2|1.67|||||||||1|1|2|1|1|1|1.17|||||||||4|4|4|4||||||1|1|5|1|2|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||8.2||1|1|1|1|F|Black||12|No|Mother|28211|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||27|28205|Some College||Medical|28269|0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020910|504471617|504473895|31|0|2|504458762|31|0|2|500897003|2||-2||2|1|500007920, 500011315, 500011316||-2||-2|0|10|||17159|12|||1|1049879|-1|4|3|44|1545381051186164660
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-07-06|NaT|Baseline|2016-07-05|2016-07-06|Complete|Done|4|4|4|4|1|4|3.5|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||5|2|2|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Cabarrus County||8||1|1|1|1|F|Hispanic||10|No|Mother|28027|3|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|F|White||47|28081||Married|Finance: Banking||18|5|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504724296|504726733|3|0|2|504746325|1|0|2|500898734|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|1056807|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-07-22|NaT|Baseline|2014-10-22|2016-07-22|Complete|Done|3|2|2|2|3|3|2.5|||||||||1|3|4|2|2|3|2.5|||||||||3|3|3|3||||||3|4|4|4|3.75|||||||4|4|4|3|4|4|4|3.86||||||||||2|3|3|2.67||||||2|2|2|||||1|1||||4|4||||Green|PERL 2014-2016||7.5||1|1|2|2|M|Black||14|No|GrandMother|28208|7|One Parent: Female|$20,000 to $24,999|Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||29|28209|Masters Degree|Single|Business|29707|0|8|Community Engagement|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|503711736|503713702|31|0|1|501121735|1|0|1|500898534|2||-2||2|1|500014681||-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||18809|8|||1|807303|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-07-25|NaT|Baseline|2016-06-02|2016-07-25|Complete|Done|3|3|2|4|4|4|3.33|||||||||1|4|3|1|1|3|2.17|||||||||4|4|4|4||||||4|5|3|2|3.5|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||1|1|1|||||1|1||||4|4||||Green|PERL 2014-2016||7.4||1|1|1|1|F|Black||12|No|Mother|28216|6|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||29|28269|Some College|Single|Business: Sales|28262|1|0|Community Engagement|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504628514|504630931|31|0|2|504599441|31|0|2|500899221|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||18809|8|||1|1041155|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-07-28|NaT|Baseline|2016-05-23|2016-07-27|Complete|Done|3|4|4|4||4||||||||||1|4|3|4|2|3|2.83|||||||||4|4|4|4||||||1|5|5|5|4|||||||||||||3|||||||||||4|4|3|3.67||||||4|1|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||7.3||1|1|1|1|F|Black||9|No|Mother|28217||One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Some Other Race||25|28208|Bachelors Degree|Single|Business: Sales|28278|0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504601619|504604030|31|0|2|504611053|41|0|2|500900279|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||46|2|||1|1030413|-1|4|3|44|727731964632783453
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-07-28|NaT|Baseline|2016-06-27|2016-07-27|Complete|Done|4|2|3|1|3|2|2.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|||7.3||1|1|1|1|F|Black||11|No|Mother|28215|6|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||30|28209|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28204|2|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504671571|504673998|31|0|2|504308223|1|0|2|500898271|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1|1054180|-1|4|3|44|20998188998147742
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-05|NaT|Baseline|2014-10-14|2016-08-05|Complete|Done|4|2|2|4|4|4|3.33|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|Cabarrus County||7||1|1|1|1|F|Black||11|No|Mother|28027|4|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||35|28027|Masters Degree|Married|Medical: Nurse||0|6|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504026659|504028677|31|0|2|504744796|31|0|2|500901331|2||500016307||2|1|500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|3|||7464|9|||1|803145|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-11|NaT|Baseline|2016-08-09|2016-08-11|Complete|Done|2|1|3|4|1|1|2|||||||||2|2|3|2|4|3|2.67|||||||||4|4|4|4||||||5|2|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||6.8||1|1|1|1|F|Black||11|No|Mother|28025|4|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||25|28027|Some College|Single|Business: Sales||0|6|Community Engagement|Special Event|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504711954|504714390|31|0|2|504718024|1|0|2|500902765|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||18809|8|||1|1068488|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-17|NaT|Baseline|2016-08-16|2016-08-17|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|4|3|2|2|4|2.83|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||6.6||1|1|1|1|M|Black||13|Yes|Mother|28025|6|One Parent: Female|$40,000 to $44,999||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||53|28027|Bachelors Degree|Married|Finance: Banking||11|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|502392338|502392776|31|0|1|504744814|1|0|1|500903717|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7464|9|||1|1070261|-1|4|3|44|2806833304218536184
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-23|NaT|Baseline|2016-02-22|2016-08-23|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||6.4||1|1|1|1|M|Black||10|No|Mother|28277|3|One Parent: Female|$40,000 to $44,999||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||45|28210|Masters Degree|Divorced|Finance: Banking|28202|10|11|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504022991|504025006|31|0|1|504545438|31|0|1|500903682|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1|996615|-1|4|3|44|5969614404793803539
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-30|NaT|Baseline|2015-11-17|2016-08-30|Complete|Done|3|2|4|3|3|4|3.17|||||||||2|3|3|3|2|3|2.67|||||||||4|3|4|3.67||||||3|4|3|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||1|1|1|||||1|1||||4|4||||Green|||6.2||1|1|1|1|F|Multi-race (Black & White)||13|No|Foster Parent|28214|6|Two Parent|$60,000 to $74,999||No||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||34|28209|Doctor of Medicine (MD)||Medical|28202|0|4|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504338170|504340392|36|0|2|504465810|31|0|2|500904260|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|5|||17159|12|||1|962749|-1|4|3|44|2806833304218536184
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-30|NaT|Baseline|2016-08-03|2016-08-30|Complete|Done|4|3|4|4|4|4|3.83|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||4|3|3|1|2.75|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||6.2||1|1|3|3|M|Black||12|No|Mother|28262|6|One Parent: Female|$20,000 to $24,999||Yes||School|General Community||Match Support|M|Black||25|28269|Masters Degree|Single|Finance|28202|0|1|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504275306|504277506|31|0|1|504359606|31|0|1|500901552|2||-2||2|1|||-2|500014681|-1|0|4|||12831|3|||1|1067176|-1|4|3|44|7674215580094440446
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-30|NaT|Baseline|2016-08-10|2016-08-30|Complete|Done|4|1|3|3|4|4|3.17|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||2|4|3|3||||||4|4|4|||||2|2||||4|4||||Green|||6.2||1|1|2|2|M|Black||10|No|Mother|28277|3|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||51|28277|Bachelors Degree|Married|Finance|28277|0|0|Igniting Breakfast|Special Event|Big|General Community|mentor2.0, mentor2.0 2014|Match Support|277|60|598|500000170|500017732|504660516|504662943|31|0|1|503922166|1|0|1|500902981|2||-2||2|1|||-2|500014505, 500014506|-2|0|10|||17266|8|||1|1068870|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-08-30|NaT|Baseline|2016-08-15|2016-08-26|Complete|Done|2|4|4|4|4|3|3.5|||||||||2|4|4|4|1|4|3.17|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|1|2.33||||||3|3|3|||||2|2||||4|4||||Green|||6.2||1|1|1|1|M|Multi-race (Black & Hispanic)||15|No|Mother|28269|8|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|M|White||33|28203|Juris Doctorate (JD)|Married|Law: Lawyer|28202|2|7|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504148143|504125727|38|0|1|504559007|1|0|1|500903465|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1069856|-1|4|3|44|887254134148570071
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-01|NaT|Baseline|2016-08-30|2016-09-01|Complete|Done|3|2|1|1|1|2|1.67|||||||||2|4|4|2|3|4|3.17|||||||||3|4|4|3.67||||||3|5|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||6.1||1|1|1|1|M|Black||12|No|Mother|28215|4|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28203|Bachelors Degree|Single|Business: Sales|28202|0|3|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504280334|504282534|31|0|1|504556921|1|0|1|500905599|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|4|||18809|8|||1|1073776|-1|4|3|44|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-06|NaT|Baseline|2016-08-18|2016-09-06|Complete|Done|3|1|4|2|1|3|2.33|||||||||2|4|2|4|1|4|2.83|||||||||3|3|2|2.67||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|2|3.71||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Green|||6||1|1|1|1|M|Black||10|Yes|Mother|28212|2|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||24|28202|Bachelors Degree|Single|Finance: Banking|28202|0|2|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504260162|504262304|31|0|1|504639207|1|0|1|500903992|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1070814|-1|4|3|44|4802885652788112046
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-09|NaT|Baseline|2016-09-02|2016-09-09|Complete|Done|3|4|4|4|3|3|3.5|||||||||3|3|4|1|4|4|3.17|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Red|Cabarrus County||5.9||1|1|1|1|F|Black||13|No|Mother|28025|7|One Parent: Female|$40,000 to $44,999||No||Self|General Community|Cabarrus County|Match Support|F|Black||47|28075|Masters Degree|Married|Finance: Banking|28282|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504633835|504636246|31|0|2|504775410|31|0|2|500906055|2||500016307||2|3|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7496|10|||1|1074821|-1|4|3|44|7410064544211008071
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-15|NaT|Baseline|2016-09-01|2016-09-13|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||5.7||1|1|2|2|M|Black||12|No|Mother|28215|5|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|Black||54|28262|Bachelors Degree|Married|Business||7|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504310625|504312843|31|0|1|503442370|31|0|1|500905889|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||7464|9|||1|1074516|-1|4|3|44|7399582438680751686
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-19|NaT|Baseline|2016-09-07|2016-09-19|Complete|Done|3|4|4|2|1|3|2.83|||||||||1|4|3|4|2|3|2.83|||||||||2|2|2|2||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||2|4|4|3.33||||||3|4|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||5.6||1|1|1|1|F|Black||9|No|Mother|28216|3|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|Black||42|28105|Bachelors Degree|Married|Business|28277|0|2|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504604960|504607371|31|0|2|504374080|31|0|2|500906296|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||46|2|||1|1075377|-1|4|3|44|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-20|NaT|Baseline|2016-08-23|2016-09-20|Complete|Done|4|1|2|2|3|3|2.5|||||||||2|4|3|1|2|3|2.5|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||5.5||1|1|1|1|M|Black||12|No|Mother|28212|4|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||28|28205|Bachelors Degree|Married|Business: Sales|28209|0|10|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504260159|504262304|31|0|1|504639152|1|0|1|500904577|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1071886|-1|4|3|44|4802885652788112046
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-21|NaT|Baseline|2016-06-23|2016-09-21|Complete|Done|3|2|3|2|4|3|2.83|||||||||1|2|2|2|2|2|1.83|||||||||4|2|2|2.67||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|||5.5||1|1|1|1|M|White||10|No|Mother|28226|3|One Parent: Female|$35,000 to $39,999|Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||30|28226|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|1|Other|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504379951|504382189|1|0|1|504736110|1|0|1|500905929|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|10|||7671|13|||1|1052656|-1|4|3|44|1706608681384859512
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-22|NaT|Baseline|2016-09-01|2016-09-22|Complete|Done|3|3|3|2|2|3|2.67|||||||||3|4|3|2|2|4|3|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||5.5||1|1|1|1|M|Black||9|No|Mother|28273|3|One Parent: Female|$35,000 to $39,999||Yes||School|General Community||Match Support|M|White||41|28226|Bachelors Degree|Married|Business: Sales|28273|4|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504403567|504405809|31|0|1|504689704|1|0|1|500905927|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1074565|-1|4|3|44|4318803846885526429
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-23|NaT|Baseline|2015-10-07|2016-09-21|Complete|Done|3|1|4|3|4|4|3.17|||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||4|4|3|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||5.4||1|1|1|1|F|Black||11|No|Mother|28212|5|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||37|28227|Bachelors Degree|Married|Business: Mgt, Admin|28173|10|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504357732|504359958|31|0|2|504576046|1|0|2|500909829|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1|941865|-1|4|3|44|6692528426538080183
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-28|NaT|Baseline|2016-09-13|2016-09-27|Complete|Done|3|3|4|3|3|4|3.33|||||||||2|4|4|3|4|4|3.5|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|PERL 2014-2016||5.3||1|1|1|1|F|Black||12|No|Mother|28269||One Parent: Female|$25,000 to $29,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||28|28203|Bachelors Degree|Single|Finance: Banking|28203|0|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504489376|504491661|31|0|2|504604779|1|0|2|500907166|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||7464|9|||1|1076882|-1|4|3|44|7341607196510895077
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-09-29|NaT|Baseline|2016-09-14|2016-09-27|Complete|Done|4|2|1|1|4|4|2.67|||||||||2|4|3|2|3|4|3|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||5.2||1|1|1|1|F|Black||11|No|Mother|28031|4|Two Parent|$15,000 to $19,999|Y|No||School|General Community|PERL 2014-2016|Match Support|F|White||44|28031|Masters Degree|Married|Education||0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500017732|504577421|504579758|31|0|2|504771021|1|0|2|500907629|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|1077436|-1|4|3|44|7137064858903755892
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-03|NaT|Baseline|2016-09-07|2016-10-03|Complete|Done|4|3|4|2|3|4|3.33|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||3|2|5|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green|||5.1||1|1|1|1|M|Black||10|No|GrandMother|28212|4|One Parent: Female|$10,000 to $14,999|Y|No||School|General Community|PERL 2014-2016|Match Support|M|White||48|28211|Masters Degree|Married|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504592676|504595050|31|0|1|504742988|1|0|1|500906468|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|1075490|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-03|NaT|Baseline|2016-09-16|2016-09-28|Complete|Done|3|1|2|1|4|4|2.5|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green|||5.1||1|1|1|1|M|Black||10|No|Mother|28273|3|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||33|28273|Bachelors Degree|Married|Tech: Computer/Programmer|28262|9|4|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504391010|504393249|31|0|1|504614273|1|0|1|500908114|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1078158|-1|4|3|44|703802826159951755
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-10|NaT|Baseline|2016-09-06|2016-10-10|Complete|Done|3|2|1|1|2|3|2|||||||||3|3|4|3|4|4|3.5|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016||4.9||1|1|1|1|M|Black||11|No|Mother|28210|5|One Parent: Female|$50,000 to $59,999||No||Self|General Community|PERL 2014-2016|Match Support|M|Native Hawaiian or Other Pacific Islander||26|28209|Bachelors Degree|Single|Business: Engineer|28202|1|8|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504714089|504716526|31|0|1|504679648|5|0|1|500906166|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|1075177|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-10|NaT|Baseline|2016-09-20|2016-10-10|Complete|Done|3|1|1|1|1|1|1.33|||||||||4|1|3|4|4|3|3.17|||||||||4|4|4|4||||||5|5|3|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||1|1||||4|4||||Green|||4.9||1|1|2|2|M|Black||10|Yes|Mother|28214|4|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||30|28209|Bachelors Degree|Married|Real Estate: Realtor|28217|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020910|504759201|504761658|31|0|1|504322037|1|0|1|500908756|2||-2||2|1||500014681|-2||-2|0|10|||46|2|||1|1079039|-1|4|3|44|7105699653014118193
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-15|NaT|Baseline|2015-12-15|2016-10-15|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|Cabarrus County||4.7||1|1|1|1|M|Black||13|No|Mother|28027|7|One Parent: Female|$50,000 to $59,999||Yes||Self|General Community|Cabarrus County|Match Support|M|White||32|28027|Some College|Married|Business: Sales|28216|5|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504507408|504509703|31|0|1|504651211|1|0|1|500913035|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|974325|-1|4|3|44|4173153455025080196
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-10-17|2017-02-23|Baseline|2016-02-10|2016-10-11|Complete|Done||1|1|1|2|2||||||||||2|4|4|3|1|4|3|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||2|2|2|2|3|3|1|2.14||||||||||3|4|4|3.67||||||4|3|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|4.2||1|1|1|1|M|Black||15|No|Mother|28211|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||34|28209||Married|Business: Sales||0|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504039275|504041293|31|0|1|504461897|1|0|1|500908017|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|992934|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-19|NaT|Baseline|2016-09-21|2016-10-19|Complete|Done|3|4|3|4|3|3|3.33|||||||||2|4|3|3|2|3|2.83|||||||||4|3|3|3.33||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Green|||4.6||1|1|1|1|M|Black||9|No|Mother|28262|2|One Parent: Female|$50,000 to $59,999||No||School|General Community||Match Support|M|Black||35|28269|Masters Degree|Married|Business: Sales|29708|2|3|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504203765|504205876|31|0|1|504766376|31|0|1|500909175|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||4748|14|||1|1079634|-1|4|3|44|3402014428779854546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-20|NaT|Baseline|2016-09-13|2016-10-19|Complete|Done|3|4|4|4|3|4|3.67|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|3|3.67||||||4|2|3|||||1|1||||4|4||||Green|PERL 2014-2016||4.5||1|1|1|1|M|Black||10|No|Mother|28216|4|One Parent: Female|Less than $10,000|Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28203|Bachelors Degree|Single|Finance: Banking|28281|3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504647175|504649586|31|0|1|504759286|1|0|1|500907299|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|1076979|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-20|NaT|Baseline|2016-09-16|2016-10-19|Complete|Done|3|4|4|3|4|3|3.5|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||2|5|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|||4.5||1|1|1|1|M|Black||12|No|GrandMother|28212|6|One Parent: Female|$10,000 to $14,999|Y|No||School|General Community||Match Support|M|White||26|28210|Bachelors Degree|Married|Business: Sales|28277|0|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504592666|504595050|31|0|1|504625671|1|0|1|500908174|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1078208|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-21|NaT|Baseline|2016-09-20|2016-10-21|Complete|Done|3|4|4|3|4|4|3.67|||||||||2|3|3|2|3|3|2.67|||||||||4|3|3|3.33||||||2|4|5|4|3.75|||||||4|4|4|3|3|3|3|3.43||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||3|3||||Green|||4.5||1|1|1|1|M|White||14|No|Mother|28212|7|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|M|White||28|28205|Bachelors Degree|Single|Tech: Sales, Mktg|28202|3|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504574961|504577295|1|0|1|504676344|1|0|1|500908810|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1079095|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-23|NaT|Baseline|2016-10-16|2016-10-23|Complete|Done|2|1|1|2|1|1|1.33|||||||||3|3|4|2|2|4|3|||||||||3|4|4|3.67||||||3|2|3|5|3.25|||||||4|4|4|4|4|3|4|3.86||||||||||3|4|4|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||4.4||1|1|1|1|F|White||12|No|Non-Relative: Other|28205|5|Two Parent|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|F|White||25|28207|Bachelors Degree|Single|Tech: Computer/Programmer|28202|1|5|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500021785|504536121|504538455|1|0|2|504562411|1|0|2|500916158|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|1089554|-1|4|3|44|2082620892288628337
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-24|NaT|Baseline|2016-09-20|2016-10-24|Complete|Done|4|1|3|1|3|4|2.67|||||||||3|3|3|1|4|4|3|||||||||4|4|4|4||||||4|3|2|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||4.4||1|1|1|1|M|Multi-race (Black & White)||11|No|Mother|28212|6|One Parent: Female|$50,000 to $59,999||Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||22|28202|Bachelors Degree|Single|Tech: Sales, Mktg|28202|0|2|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|503623886|503625775|36|0|1|504803107|1|0|1|500915035|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|1078937|-1|4|3|44|5499465424599250965
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-10-26|2017-02-23|Baseline|2016-10-12|2016-10-25|Complete|Done|3|3|4|3|4|3|3.33|||||||||2|2|4|2|2|3|2.5|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|2|1.5|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|3.9||1|1|1|1|M|Black||10|No|Mother|28208|3|One Parent: Female|$35,000 to $39,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business|28203|2|9|BBBS National Site|Web Link|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|503401421|503403278|31|0|1|504818783|1|0|1|500916185|2||-2||4|1|||-2|500007920, 500011315, 500011316|-1|34|2|||46|2|||1|1087576|-1|4|3|44|5096023753338979088
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-28|NaT|Baseline|2016-10-20|2016-10-28|Complete|Done|2|2|3|2|4|3|2.67|||||||||4|4|4|3|4|3|3.67|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||4.3||1|1|1|1|M|White||12|No|Mother|28226|6|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community||Match Support|M|White||31|28205|Bachelors Degree|Single|Real Estate: Realtor|28202|1|6|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504436181|504438437|1|0|1|504741299|1|0|1|500921121|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1091915|-1|4|3|44|6694016660882153370
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-28|NaT|Baseline|2016-10-21|2016-10-28|Complete|Done|4|4|4|2|4|4|3.67|||||||||3|3|4|3|4|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red|PERL 2014-2016, Cabarrus County||4.3||1|1|4|4|F|Black||14|No|Mother|28027|6|Two Parent|$60,000 to $74,999|Y|No|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Multi-race (Black & White)||23|28273|Some College|Single|Student: College|28227|0|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504655474|504657901|31|0|2|503853917|36|0|2|500918496|2||500016307||2|3|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||7464|9|||1|1092531|-1|4|3|44|7048951337647301192
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-31|NaT|Baseline|2016-09-21|2016-10-31|Complete|Done|4|2|3|3|3|4|3.17|||||||||3|3|3|4|4|3|3.33|||||||||4|4|4|4||||||4|2|2|4|3|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|3|3.67||||||3|2|2.5|||||1|1||||4|4||||Green|||4.2||1|1|1|1|M|White||12|No|Mother|28031|6|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||28|28031|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|7|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504417121|504419373|1|0|1|504579745|1|0|1|500909172|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|1079633|-1|4|3|44|458920933571351085
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-31|NaT|Baseline|2016-09-28|2016-10-31|Complete|Done|3|3|4|4|3|3|3.33|||||||||4|3|3|3|4|3|3.33|||||||||4|4|4|4||||||5|3|4|2|3.5|||||||3|4|4|3|3|4|4|3.57||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||4.2||1|1|1|1|M|Black||15|No|Mother|28105|9|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|Black||30|28105|Bachelors Degree|Married|Business|28078|0|7|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504698283|504700711|31|0|1|504765309|31|0|1|500918562|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|56|1|||7464|9|||1|1082280|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-31|NaT|Baseline|2016-10-07|2016-10-31|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|3|4|3|3|4|3.33|||||||||4|4|3|3.67||||||5|5|4|5|4.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|||||||2|2||||4|4||||Green|||4.2||1|1|1|1|M|Black||13|No|Mother|28215|7|One Parent: Female|$40,000 to $44,999||Yes||Self|General Community||Match Support|M|Multi-race (Hispanic & White)||28|28205|Bachelors Degree|Married|Finance: Banking|28202|1|4|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504564027|504566361|31|0|1|504766711|35|0|1|500913521|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1085878|-1|4|3|44|2806833304218536184
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-31|NaT|Baseline|2016-10-12|2016-10-31|Complete|Done|4|3|4|1|3|4|3.17|||||||||2|1|2|4|4|4|2.83|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|2|3.71||||||||||4|3|4|3.67||||||4|4|4|||||2|2||||4|4||||Green|||4.2||1|1|1|1|M|Black||9|No|Mother|28212|3|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|White||32|28209||Single|Finance|28202|2|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504392725|504394964|31|0|1|504697126|1|0|1|500914996|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1087780|-1|4|3|44|3727915399477748546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-31|NaT|Baseline|2016-10-12|2016-10-31|Complete|Done|4|2|4|2|3|4|3.17|||||||||2|4|4|3|3|4|3.33|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||1|1||||4|4||||Green|||4.2||1|1|1|1|M|Black||9|No|Mother|28212||One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||33|28202|PHD|Single|Real Estate: Realtor|28269|3|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504399529|504394964|31|0|1|504803637|1|0|1|500915028|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1087843|-1|4|3|44|3727915399477748546
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-31|NaT|Baseline|2016-10-13|2016-10-26|Complete|Done|3|2|3|2|3|4|2.83|||||||||4|4|4|4|4|4|4|||||||||3|4|2|3||||||5|4|2|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5||||||||||4|4||||Green|||4.2||1|1|1|1|M|Multi-race (Black & White)||12|No|Mother|28078|5|One Parent: Female|$40,000 to $44,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||31|28078|Some College|Married|Business: Sales|28078|0|5|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504416044|504418296|36|0|1|504623074|1|0|1|500918304|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1088445|-1|4|3|44|7269080898586176194
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-10-31|NaT|Baseline|2016-10-17|2016-10-31|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|3|4|3|3|4|3.5|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|||4.2||1|1|1|1|M|Black||10|Yes|Mother|28208|3|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community||Match Support|M|Black||46|28277|Some College|Married|Business|28277|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504401349|504403590|31|0|1|504856770|31|0|1|500921965|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1089892|-1|4|3|44|4309014537710246316
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-12|NaT|Baseline|2016-10-17|2016-11-12|Complete|Done|2|2|2|2|2|2|2|||||||||3|3|3|2|3|3|2.83|||||||||4|4|4|4||||||3|4|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|Cabarrus County||3.8||1|1|1|1|F|Black||13|No|Mother|28025|7|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|Cabarrus County|Match Support|F|White||41|28027|Masters Degree|Married|Homemaker||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504792692|504795152|31|0|2|504760167|1|0|2|500916273|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|1089720|-1|4|3|44|3918615128866826495
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-14|NaT|Baseline|2016-09-16|2016-11-14|Complete|Done|4|2|4|1|4|4|3.17|||||||||2|3|4|2|2|4|2.83|||||||||4|4|4|4||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green|||3.7||1|1|1|1|F|Black||11|No|Mother|28269|6|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||39|28269|Bachelors Degree|Single|Govt|28202|1|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504628103|504630514|31|0|2|504469742|31|0|2|500922796|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1|1078161|-1|4|3|44|4825213036474521167
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-14|NaT|Baseline|2016-10-21|2016-11-14|Complete|Done|4|1|1|1|3|4|2.33|||||||||1|3|3|1|4|4|2.67|||||||||4|4|4|4||||||5|2|4|3|3.5|||||||4|4|4|4|4|4|3|3.86|||||||||||||||||||4|3|3.5|||||2|2|||||||||Green|||3.7||1|1|1|1|M|Black||11|Yes|Mother|28217|4|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||27|28278||Single|Business|28208|0|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504456498|504458770|31|0|1|504766383|1|0|1|500918854|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|1092391|-1|4|3|44|5597049740348738
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-16|NaT|Baseline|2016-10-23|2016-11-15|Complete|Done|4|2|3|4|4|4|3.5|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green|||3.6||1|1|1|1|F|Black||10|No|Mother|28211|5|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||39|28277|Masters Degree|Married|Education||3|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504835647|504838149|31|0|2|504545759|31|0|2|500918758|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1|1092977|-1|4|3|44|8726431331992650796
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-16|NaT|Baseline|2016-11-14|2016-11-16|Complete|Done|2|2|2|2|2|1|1.83|||||||||2|3|4|4|2|3|3|||||||||4|4|4|4||||||4|2|5|4|3.75|||||||3|3|3|3|3|3|3|3||||||||||1|3|3|2.33||||||3|4|3.5|||||1|1||||4|4||||Green|PERL 2014-2016, Cabarrus County||3.6||1|1|1|1|M|White||13|No|Foster Parent|28027|6|One Parent: Male|$100,000 to $124,999|Y|No|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||28|28269|Bachelors Degree|Single|Medical|46250|0|7|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504748250|504750703|1|0|1|504885284|1|0|1|500927298|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||17159|12|||1|1104179|-1|4|3|44|71389706163855294
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-16|NaT|Baseline|2016-11-15|2016-11-16|Complete|Done|4|4|4|3|2|4|3.5|||||||||4|4|4|2|2|4|3.33|||||||||3|3|2|2.67||||||4|5|2|5|4|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||3.6||1|1|1|1|M|White||10|No|Mother|28081|5|One Parent: Female|$10,000 to $14,999|Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||25|28027||Married|Medical: Healthcare Worker||0|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504862022|504864541|1|0|1|504930361|1|0|1|500927996|2||-2||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|34|2|||7671|13|||1|1105162|-1|4|3|44|2036270106764562772
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-21|NaT|Baseline|2016-11-18|2016-11-21|Complete|Done|3|3|4|3|3|3|3.17|||||||||2|3|3|3|3|3|2.83|||||||||4|3|3|3.33||||||2|4|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|3|3|3.33||||||2|3|2.5|||||1|1||||4|4||||Green|Cabarrus County||3.5||1|1|1|1|M|Black||13|No|Mother|28025|7|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|Cabarrus County|Match Support|M|Black||29|28027|Bachelors Degree|Married|Business||0|10|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504732530|504734976|31|0|1|504893030|31|0|1|500929513|2||-2||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|5|||7464|9|||1|1107317|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-28|NaT|Baseline|2016-11-11|2016-11-22|Complete|Done|3|2|3|2|2|3|2.5|||||||||4|4|4|2|4|3|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||3.3||1|1|1|1|M|White||13|No|Mother|28277|8|One Parent: Female|$60,000 to $74,999||No||Self|General Community|PERL 2014-2016|Match Support|M|White||26|28207|Masters Degree|Living w/ Significant Other|Tech: Engineer|28203|1|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504808434|504810913|1|0|1|504557160|1|0|1|500926948|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|1103507|-1|4|3|44|5571803589598086587
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-29|NaT|Baseline|2016-09-16|2016-11-29|Complete|Done|3|2|1|1|2|2|1.83|||||||||2|3|2|2|2|2|2.17|||||||||3|3|3|3||||||1|2|4|5|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||1|1||||4|4||||Green|||3.2||1|1|1|1|F|Black||15|No|Mother|28211|9|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||47|28215|Masters Degree|Married|Education|28202|5|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504471621|504473895|31|0|2|504580592|31|0|2|500925801|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|1078193|-1|4|3|44|1545381051186164660
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-29|NaT|Baseline|2016-10-24|2016-11-29|Complete|Done|3|2|3|2|1|4|2.5|||||||||3|3|3|2|2|3|2.67|||||||||4|4|4|4||||||3|4|1|4|3|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||3.2||1|1|1|1|F|Black||11|No|Mother|28209|5|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||23|28203|Bachelors Degree||Finance: Accountant|28031|0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504662612|504665039|31|0|2|504595097|1|0|2|500918825|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1093147|-1|4|3|44|2719955880210213907
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-30|NaT|Baseline|2016-10-20|2016-11-10|Complete|Done|3|1|1|1|1|1|1.33|||||||||1|3|1|||||||||||||4|4|4|4||||||2|1|5|4|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4||||||||||4|4||||Green|||3.2||1|1|1|1|F|White||12|Yes|Non-Relative: Other|28205|5|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|F|White||28|28202|Bachelors Degree|Single|Finance|28202|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504539986|504538455|1|0|2|504793129|1|0|2|500926111|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1092039|-1|4|3|44|2082620892288628337
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-04|NaT|Baseline|2016-11-22|2016-12-04|Complete|Done|3|3|3|3|3|2|2.83|||||||||2|3|2|2|3|2|2.33|||||||||4|3|3|3.33||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||1|4|2.5|||||2|2||||4|4||||Green|Cabarrus County||3.1||1|1|1|1|F|Black||12|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||24|28262|Masters Degree|Single|Human Services: Social Worker|28027|0|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504937152|504939686|31|0|2|504797758|31|0|2|500930335|2||500016307||2|1|500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|1108671|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-06|NaT|Baseline|2016-11-11|2016-12-06|Complete|Done|4|4|4|2|4|4|3.67|||||||||2|4|3|3|4|4|3.33|||||||||4|3|3|3.33||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||3||1|1|1|1|M|Black||12|No|Mother|28213|5|One Parent: Female|$20,000 to $24,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||33|28203|Bachelors Degree|Married|Business|32207|9|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|502383218|502383656|31|0|1|504867282|1|0|1|500926962|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|6854|8|||46|2|||1|1103521|-1|4|3|44|20998188998147742
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-21|NaT|Baseline|2016-09-16|2016-12-19|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||2.5||1|1|1|1|M|Black||15|No|Mother|28227|8|One Parent: Female|$25,000 to $29,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||25|28277|Bachelors Degree|Single|Business|28208|1|8|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504662357|504664784|31|0|1|504791469|31|0|1|500933117|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1|1078180|-1|4|1|44|3557919386369667257
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-21|NaT|Baseline|2016-10-21|2016-12-21|Complete|Done|4|1|1|1|4|4|2.5|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3||||||||||4|4||||Green|||2.5||1|1|1|1|M|Black||12|No|Mother|28210|5|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community||Match Support|M|Black||30|28210|Bachelors Degree|Married|Military||1|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504565095|504567429|31|0|1|504860995|31|0|1|500932205|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1092382|-1|4|3|44|6156547733130613405
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Completed|2016-12-22|2017-02-28|Baseline|2016-12-01|2016-12-19|Complete|Done|4|1|4|4|4|4|3.5|||||||||4|4|4|1|4|1|3|||||||||4|4|4|4||||||1|1|5|5|3|||||||4|4|4|3|3|3|4|3.57||||||||||4|4|4|4||||||1|1|1|||||1|1||||4|4||||Red||Child/Family: Moved|2.2||1|1|1|1|M|Black||14|No|Mother|28215|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Black||32|28213|Masters Degree|Married|Finance: Auditor|28202|0|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500020753|504851045|504853547|31|0|1|504774982|31|0|1|500932246|2||-2||4|3||500014681|-2|500007920, 500011315, 500011316|-2|0|5|||46|2|||1|1112091|-1|4|3|44|2141487034287122220
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-01-11|NaT|Baseline|2016-12-13|2017-01-11|Complete|Done|3|2|1|1|3|1|1.83|||||||||1|1|2|4|2|4|2.33|||||||||4|4|4|4||||||1|4|1|3|2.25|||||||4|4|4|4|4|4|3|3.86||||||||||1|4|1|2||||||3|2|2.5|||||1|1||||4|4||||Green|||1.8||1|1|1|1|F|Black||11|No|Mother|28208|4|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||24|28203|Bachelors Degree|Single|Finance|28255|0|6|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504617847|504620258|31|0|2|504580008|1|0|2|500935128|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||7462|13|||1|1116525|-1|4|3|44|8408514790530965815
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-01-30|NaT|Baseline|2016-12-06|2017-01-30|Complete|Done|2|2|4|2|3|4|2.83|||||||||4|4|4|2|4|3|3.5|||||||||3|3|4|3.33||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|2|3|||||1|1||||4|4||||Green|||1.2||1|1|1|1|M|Black||11|No|Mother|28202|4|One Parent: Female|$20,000 to $24,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||50|28210|Bachelors Degree|Married|Finance|28202|15|0|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504700175|504702604|31|0|1|504649796|1|0|1|500933583|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||18809|8|||1|1113991|-1|4|3|44|6761707515712559257
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-01-30|NaT|Baseline|2017-01-10|2017-01-30|Complete|Done|3|4|4|2|4|4|3.5|||||||||3|4|3|2|4|3|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||1.2||1|1|1|1|F|Multi-race (Black & White)||10|No|Mother|28213|5|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||38|28202|Bachelors Degree|Single|Business|28202|0|2|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504888357|504890877|36|0|2|504850919|1|0|2|500939317|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1|1124563|-1|4|3|44|4855845956679832355
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-01-30|NaT|Baseline|2017-01-11|2017-01-23|Complete|Done|2|2|3|2|1|2|2|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|2|3.33||||||4|4|4|||||1|1||||4|4||||Green|||1.2||1|1|1|1|M|Black||12|No|Mother|28217|6|One Parent: Female|$25,000 to $29,999|Y|No|BBBS National Site|Web Link|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|M|White||37|28203|Masters Degree|Single|Business: Mgt, Admin|28226|0|1|Radio|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504736266|504738712|31|0|1|504634630|1|0|1|500940290|2||-2||2|1||500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|34|2|||131|1|||1|1124975|-1|4|3|44|2876415545463317777
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-01-30|NaT|Baseline|2017-01-11|2017-01-30|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|3|2|1|3|2.83|||||||||4|4|1|3||||||3|5|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|2|3||||||2|2|2|||||1|1||||4|4||||Green|||1.2||1|1|4|4|M|Black||12|No|Mother|28134|5|One Parent: Female|$50,000 to $59,999|Y|Yes||Self|General Community||Match Support|M|Black||43|28173|Masters Degree|Married|Finance: Banking|28281|7|0|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504675071|504677498|31|0|1|500353496|31|0|1|500942748|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1|1124998|-1|4|3|44|3894730386800788938
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-04|NaT|Baseline|2017-01-27|2017-02-04|Complete|Done|3|4|4|4|3|4|3.67|||||||||3|4|3|1|2|4|2.83|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||2|3|2.5|||||2|2||||4|4||||Green|Cabarrus County||1||1|1|1|1|M|Black||10|No|Mother|28027|5|One Parent: Female|$15,000 to $19,999||Yes||School|General Community|Cabarrus County|Match Support|M|Black||34|28227|Juris Doctorate (JD)|Separated|Law: Lawyer|28227|9|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504937135|504939686|31|0|1|504694440|31|0|1|500942634|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1130620|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-08|NaT|Baseline|2017-01-11|2017-02-08|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4||4|4|4||||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||0.9||1|1|1|1|M|Black||10|No|Mother|28211|2|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|M|Black||38|28227|Bachelors Degree|Single|Business: Marketing|28202|4|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504417080|504419332|31|0|1|504872445|31|0|1|500939553|2||-2||2|1||500007920, 500011315, 500011316, 500014681|-2|500007920, 500011315, 500011316|-2|0|5|||46|2|||1|1124976|-1|4|3|44|2763237020791144915
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-11|NaT|Baseline|2017-02-02|2017-02-11|Complete|Done|2|1|1|1|1|3|1.5|||||||||1|1|3|1|2|2|1.67|||||||||4|4|4|4||||||1|3|1|4|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|2|1.5|||||1|1||||4|4||||Green|Cabarrus County||0.8||1|1|1|1|F|White||13|No|Mother|28025|8|Two Parent|Unknown|Y|Yes||Therapist/Counselor|General Community|Cabarrus County|Match Support|F|White||31|28025||Separated|Business||0|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|504999127|505001687|1|0|2|504999362|1|0|2|500944301|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|5|||17159|12|||1|1133206|-1|4|3|44|6915279604152465197
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-17|NaT|Baseline|2017-02-06|2017-02-16|Complete|Done|3|4|1|1|3|1|2.17|||||||||1|4|4|4|1|3|2.83|||||||||4|4|4|4||||||5|4|5|3|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||0.6||1|1|1|1|M|Black||10|No|Mother|28269|3|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community||Match Support|M|White||24|28208|Bachelors Degree|Single|Tech: Management|28203|0|5|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504811851|504814332|31|0|1|504883582|1|0|1|500944658|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|3|||7464|9|||1|1134028|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-19|NaT|Baseline|2017-02-09|2017-02-19|Complete|Done|4|3|4|3|3|4|3.5|||||||||3|3|3|3|2|3|2.83|||||||||4|2|2|2.67||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|Cabarrus County||0.5||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28027|5|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|Black||54|28075|Masters Degree|Married|Business||0|9|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|504819474|504821973|36|0|1|505001672|31|0|1|500945474|2||500016307||2|1|500016374||-2|500016374|-2|0|10|||7464|9|||1|1135320|-1|4|3|44|0
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-19|NaT|Baseline|2017-02-14|2017-02-19|Complete|Done|3|1|2|3|3|4|2.67|||||||||2|4|4|3|4|3|3.33|||||||||4|4|4|4||||||5|2|4|5|4|||||||1|4|4|3|4|4|3|3.29||||||||||4|3|2|3||||||4|4|4|||||1|1||||4|4||||Green|Cabarrus County||0.5||1|1|2|2|M|Black||9|No|Mother|28081|3|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||24|28081|Some High School|Single|Service: Hotel||4|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|504902017|504904537|31|0|1|501028238|31|0|1|500946229|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|10|||17159|12|||1|1136700|-1|4|3|44|2544020271035850193
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-20|NaT|Baseline|2016-11-11|2017-02-17|Complete|Done|3|3|4|2|3|3|3|||||||||2|3|3|2|2|2|2.33|||||||||4|3|3|3.33||||||3|4|2|2|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||2|3|2|2.33||||||2|3|2.5|||||1|1||||4|4||||Green|||0.5||1|1|1|1|F|Hispanic||13|No|Mother|28226|7|One Parent: Female|$10,000 to $14,999||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Hispanic|Mexican|22|28227|Bachelors Degree|Single|Tech: Management|28202|0|4|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504672339|504674766|3|0|2|504870474|3|10|2|500941713|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|1103515|-1|4|3|44|5081726734274569781
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-23|NaT|Baseline|2017-01-10|2017-02-23|Complete|Done|4|4|4|3|1|4|3.33|||||||||1|4|4|2|1|4|2.67|||||||||4|3|2|3||||||3|3|5|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||2|2||||4|4||||Green|||0.4||1|1|2|2|M|Black||10|No|Mother|28214|2|One Parent: Female|$25,000 to $29,999||No|BBBS National Site|Web Link|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|504486089|504488364|31|0|1|502643791|3|0|1|500944356|2||-2||2|1|||-2||-2|34|2|||7496|10|||1|1124567|-1|4|3|44|6570326659017849719
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-23|NaT|Baseline|2017-01-11|2017-02-23|Complete|Done|4|2|3|2|4|2|2.83|||||||||4|4|3|3|2|4|3.33|||||||||4|3|4|3.67||||||3|4|5|5|4.25|||||||4|4|4|4|2|4|3|3.57||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|||0.4||1|1|1|1|M|Black||12|No|Foster Parent|28215|6|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|M|Black||25|28223|Bachelors Degree|Single|Business|28202|1|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500013781|504463138|504465396|31|0|1|504819424|31|0|1|500947979|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|1124991|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-23|NaT|Baseline|2017-02-08|2017-02-23|Complete|Done|4|2|3|2|4|4|3.17|||||||||3|4|2|3|3|3|3|||||||||4|4|3|3.67||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|1|1.5|||||2|2||||3|3||||Green|||0.4||1|1|1|1|M|Black||13|Yes|GrandMother|28214|7|Grandparents|$75,000 to $99,999|Y|Yes||Self|General Community||Match Support|M|White||31|28078|Bachelors Degree|Single|Business: Sales|28202|4|9|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504910266|504912793|31|0|1|504829494|1|0|1|500945213|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1|1134834|-1|4|3|44|5163136606149365864
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-27|NaT|Baseline|2017-02-06|2017-02-20|Complete|Done|3|2|1|2|2|2|2|||||||||3|3|2|4|2|3|2.83|||||||||4|4|4|4||||||3|3|3|5|3.5|||||||4|4|4||4|4|2|||||||||||3|4|2|3||||||1|3|2|||||1|1||||4|4||||Green|||0.3||1|1|1|1|F|Black||9|No|Mother|28269|3|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Multi-race (Black & White)||21|28213|Some College|Single|Business: Sales|28211|0|9|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504673056|504675483|31|0|2|504845407|36|0|2|500944794|2||-2||2|1||500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1134179|-1|4|3|44|7044657180546140448
BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2017-02-28|NaT|Baseline|2017-02-07|2017-02-27|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|2|2|3|3|2|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||0.2||1|1|1|1|M|Black||10|No|Mother|28277|5|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|M|White||31|28277|Masters Degree|Married|Finance: Accountant|28273|0|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504838542|504838321|31|0|1|504930064|1|0|1|500945724|2||-2||2|1||500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|1134613|-1|4|3|44|2742327884002010428
