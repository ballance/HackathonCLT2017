ChildPartKey|AgencyName|TeamName|MatchType|MatchStatus|MatchOpenDate|MatchCloseDate|SurveyType|YOSScheduledDate|YOSCompletionDate|YOSCompletionType|YOSStatus|Q1|Q2Neg|Q3Neg|Q4Neg|Q5|Q6|SocAccept|Q1b|Q2b|Q3b|Q4b|Q5b|Q6b|SocAcceptB|SocAcceptPrcnt|Q7Neg|Q8|Q9|Q10Neg|Q11Neg|Q12|SchComp|Q7b|Q8b|Q9b|Q10b|Q11b|Q12b|SchCompB|SchCompPrcnt|Q13|Q14|Q15|EdExpect|Q13b|Q14b|Q15b|EdExpectb|EdExpectPrcnt|Q16|Q17|Q18|Q19|Grades|Q16b|Q17b|Q18b|Q19b|Gradesb|GradesPrcnt|Q20Neg|Q21Neg|Q22Neg|Q23Neg|Q24Neg|Q25Neg|Q26Neg|RiskAtt|Q20b|Q21b|Q22b|Q23b|Q24b|Q25b|Q26b|RiskAttb|RiskAttPrcnt|Q27|Q28|Q29|PTrust|Q27b|Q28b|Q29b|PTrustb|PTrustPrcnt|Q30Neg|Q31Neg|Truancy|Q30b|Q31b|Truancyb|TruancyPrcnt|Q32|SpAdult|Q32b|SpAdultb|SpAdultPrcnt|Q33Neg|JJustice|Q33b|JJusticeB|JJusticePrcnt|MatchSupportLevel|MatchReportSources|MatchClosureReasons|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildLivingSituation|ChildIncomeLevel|ChildFamilyAssistance|ChildFreeReducedLunch|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolPartKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|MatchKey|MatchTypeKey|SiteTypeKey|MatchActivityKey|SiteKey|StatusKey|MatchSupportLevelKey|MatchReportSourceKey|ChildReportSourceKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|YOSSurveyKey|PriorBaselineYOSSurveyKey|YOSStatusKey|YOSCompletionTypeKey|SurveyTypeKey
500897083|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-13|2012-11-19|Baseline|2009-11-06|2009-11-13|Complete|Done|4|1|4|1|3|4|2.83|||||||||3|3|3|4|4|4|3.5|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red|Amachi|Child/Family: Infraction of match rules/agency policies|36.2||1|1|1|1|M|Black||21|Yes|Mother|28269|One Parent: Female|Unknown|Y|No||Service Organization|General Community|Amachi|Match Support|M|White||54|28210||Married|Self-Employed, Entrepreneur||0|0|Holy Comforter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|500897335|31|0|1|501862348|1|0|1|500407273|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|11|||9216|7|||1|268|-1|4|3|44
501086649|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-20|2013-01-09|Baseline|2009-10-23|2009-11-20|Complete|Done|4|3|4|2|3|4|3.33|||||||||4|4|4|4|3|3|3.67|||||||||4|3|3|3.33||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||2|2|||||||||Red||Volunteer: Feels incompatible with child/family|37.7||1|1|1|1|M|Black||21|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Relative|General Community||Match Support|M|White||39|28205|Bachelors Degree|Single|Transport: Pilot|30320|2|0|Other Church Partner|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500004169|501086923|31|0|1|501833794|1|0|1|500399391|2||-2||4|3|||-2||-2|0|3|||7453|7|||1|385|-1|4|3|44
501313839|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-11|2013-06-18|Baseline|2009-10-19|2009-11-11|Complete|Done|3|2|3|3|4|4|3.17|||||||||2|3|4|4|2|4|3.17|||||||||3|4|4|3.67||||||4|5|5|5|4.75|||||||4|4|4|3|2|2|1|2.86||||||||||3|4|3|3.33||||||3|3|3|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|43.2||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||36|28204|Bachelors Degree|Single|Consultant||4|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501314117|31|0|1|501788563|1|0|1|500396680|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|590|-1|4|3|44
501702616|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-20|2010-10-22|Baseline|2009-11-03|2009-11-20|Complete|Done|2|4|2|1|2|2|2.17|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|3|4|2|3.57||||||||||3|3|4|3.33||||||3|3|3|||||2|2|||||||||Green||Child/Family: Moved|11||1|1|1|1|M|Black||17|No|Mother|28134|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||58|29710|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501702954|31|0|1|501849169|1|0|1|500405205|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|1183|-1|4|3|44
501670169|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2012-04-04|Baseline|2009-09-30|2009-09-30|Complete|Done|4|4|4|4|4|4|4|||||||||2||4|||4||||||||||4|4|3|3.67||||||4|2|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||4|2|3|||||1|1|||||||||Green||Volunteer: Time constraint|30.1||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|F|Black||32|28269||Single|Consultant|28209|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501670507|31|0|2|501466072|31|0|2|500379969|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|2678|-1|4|3|44
501386394|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2011-03-25|Baseline|2009-09-30|2009-09-30|Complete|Done|2|3|2|3|4|3|2.83|||||||||1|4|4|2|2|4|2.83|||||||||4|4|4|4||||||2|4|4|4|3.5|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||2|1|1.5|||||1|1|||||||||Yellow||Volunteer: Time constraint|17.8||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||RTBM|M|Black||45|28215||Married|Tech: Research/Design||0|0|Mayfield Memorial|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500001281|501386675|31|0|1|501818567|31|0|1|500388796|2||-2||4|2|||-2||-2|34|2|||9212|7|||1|3316|-1|4|3|44
501376516|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2010-07-30|Baseline|2009-09-30|2009-09-30|Complete|Done|3|1|4|2|1|4|2.5|||||||||1|3|1|4|2|3|2.33|||||||||4|3|4|3.67||||||3|4|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||1|1|||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|10||1|1|1|1|M|Black||20|Yes|Mother|28205|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Enrollment|M|White||34|28209|||Consultant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010355|501376795|31|0|1|501822933|1|0|1|500386771|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|4386|-1|4|3|44
501868921|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2010-12-21|Baseline|2009-10-30|2009-10-30|Complete|Done|3|1|1|1|1|2|1.5|||||||||3|2|4|4|4|4|3.5|||||||||4|3|3|3.33||||||4|5|5|4|4.5|||||||4|4|4|4|3|3|3|3.57||||||||||2|4|3|3||||||2|1|1.5|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|13.7||2|2|1|1|F|Black||19|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||34|28217|Juris Doctorate (JD)|Married|Law: Lawyer|28204|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501869291|31|0|2|501220647|31|0|2|500398441|2||-2||4|2||500005291|-2||-2|0|10|||7464|9|||1|4527|-1|4|3|44
501524313|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-22|2010-04-23|Baseline|2009-09-22|2009-09-22|Complete|Done|2|2|3|2|3|3|2.5|||||||||3|3|3|3|3|3|3|||||||||3|3|3|3||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Green||Child/Family: Moved|7||2|2|2|2|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||36|28278|Bachelors Degree|Single|Retail: Sales|30071|5|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500009242|501524605|31|0|1|501508941|1|0|1|500381084|2||-2||4|1||500005291|-2||-2|0|10|||7464|9|||1|4772|-1|4|3|44
501201068|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2012-08-29|Baseline|2009-10-30|2009-10-30|Complete|Done|3|2|3|2|4|4|3|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|4|5|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||1|1|||||||||Green||Child/Family: Lost contact with volunteer/agency|34||1|1|1|1|M|Black||21|No|Mother|28215|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||60|28262|Masters Degree|Single|Tech: Engineer||5|0|AA Task Force|Service Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501201342|31|0|1|501771844|31|0|1|500396764|2||-2||4|1|||-2|500000294|-2|6854|8|||9226|6|||1|5730|-1|4|3|44
501766666|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-02|2010-08-03|Baseline|2009-10-02|2009-10-02|Complete|Done|4|2|2|1|4|4|2.83|||||||||2|2|4|4|1|4|2.83|||||||||4|4|4|4||||||5|2|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green|Amachi|Child/Family: Moved|10||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||31|28211|Bachelors Degree|Single|Unknown|28209|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|501765484|31|0|2|501541222|1|0|2|500386249|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|5882|-1|4|3|44
501796006|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-03|2011-12-20|Baseline|2009-11-03|2009-11-03|Complete|Done|3|4|4|2|3|4|3.33|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4|||||||3|3|5||||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|2|3|||||2|2|||||||||Green||Volunteer: Time constraint|25.5||3|3|1|1|F|Black||17|No|Mother|28031|Two Parent|Unknown|Y|Yes||School|General Community||Match Support|F|White||37|28078|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501489205|31|0|2|501621517|1|0|2|500396069|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|6008|-1|4|3|44
501820715|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-23|2010-11-30|Baseline|2009-10-23|2009-10-23|Complete|Done|4|1|1|2|3|3|2.33|||||||||3|4|1|4|4|3|3.17|||||||||4|3|4|3.67||||||4|3|3|1|2.75|||||||4|4|4|4|2|4|4|3.71||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Green||Volunteer: Health|13.2||1|1|2|2|M|Black||22|No|Mother|28227|One Parent: Female|Unknown|Y|Yes||Relative|General Community||Match Support|M|Black||68|28212|Associate Degree|Married|Craftsman||25|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501821070|31|0|1|501049119|31|0|1|500387870|2||-2||4|1|||-2|500000294|-2|0|3|||2238|7|||1|7575|-1|4|3|44
501788773|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-27|2012-06-28|Baseline|2009-10-27|2009-10-27|Complete|Done|3|2|2|1|4|4|2.67|||||||||2|4|3|4|4|3|3.33|||||||||4|4|3|3.67||||||3|4|4|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|2|2|||||2|2|||||||||Green|Amachi|Volunteer: Moved|32||1|1|1|1|M|Black||18|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|RTBM|M|White||33|28202|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501789128|31|0|1|501845020|1|0|1|500393644|2||-2||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|7735|-1|4|3|44
501724491|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2011-03-30|Baseline|2009-10-29|2009-10-29|Complete|Done|4|2|4|1|1|4|2.67|||||||||1|1|3|1|1|2|1.5|||||||||4|4|4|4||||||2|3|5|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|4|3.67||||||4|3|3.5|||||1|1|||||||||Green||Volunteer: Moved|17||1|1|1|1|M|Multi-race (Black & Asian)||19|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|M|White||42|28216||Divorced|Medical|28078|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501724831|39|0|1|501852487|1|0|1|500397005|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|7914|-1|4|3|44
501861660|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-06|2010-02-04|Baseline|2009-11-06|2009-11-06|Complete|Done|3|4|4|3|3|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||2|4|4|4|4|4|4|3.71||||||||||3|4|4|3.67||||||4|4|4|||||1|1|||||||||Green||Volunteer: Lost contact with child/agency|3||1|1|1|1|F|Hispanic||17||Mother|28273|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|White||35|28205|Bachelors Degree|Single|Business: Mgt, Admin|28255|4|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500009242|501862033|3|0|2|501588905|1|0|2|500405168|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|9549|-1|4|3|44
501776333|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-08|2013-07-25|Baseline|2009-09-08|2009-09-08|Complete|Done|3|2|3|2|4|4|3|||||||||3|3|3|2|3|3|2.83|||||||||3|3|3|3||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|46.5||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28210|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|501776688|31|0|1|501832599|31|0|1|500381636|2||-2||4|1|||-2|500000294|-2|34|2|||7464|9|||1|9814|-1|4|3|44
501831576|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2010-08-03|Baseline|2009-09-29|2009-09-29|Complete|Done|4|4|4|3|3|4|3.67|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|2|4|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Yellow|Amachi|Volunteer: Time constraint|10.1||3|3|1|1|F|Black||18|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|White||33|28211|Bachelors Degree|Single|Medical: Admin|28211|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010355|501831944|31|0|2|501427745|1|0|2|500387626|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|11655|-1|4|3|44
501792675|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2011-09-21|Baseline|2009-09-30|2009-09-30|Complete|Done|4|4|4|1|3|4|3.33|||||||||2|4|3|2|4|3|3|||||||||4|4|4|4||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2|||||||||Green||Volunteer: Moved|23.7||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|19085|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501793030|31|0|1|501664548|1|0|1|500386328|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|12540|-1|4|3|44
501771253|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2011-04-21|Baseline|2009-09-29|2009-09-29|Complete|Done|4|1|4|1|4|4|3|||||||||2|4|4|3|3|4|3.33|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|4|3|||||||||||||||Yellow||Volunteer: Feels incompatible with child/family|18.7||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||34|28269|Bachelors Degree|Single|Medical: Nurse|28054|3|6|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500009007|501741899|31|0|2|501322818|31|0|2|500383563|2||500003586||4|2|||-2|500000294|-2|0|10|||7462|13|||1|13780|-1|4|3|44
501250109|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-11|2013-02-27|Baseline|2009-09-11|2009-09-11|Complete|Done|3|1|3|1|3|3|2.33|||||||||3|3|3|3|4|3|3.17|||||||||3|3|3|3||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Red||Volunteer: Lost contact with child/agency|41.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28227|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501250385|31|0|1|501790515|31|0|1|500381167|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|13945|-1|4|3|44
501686310|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2013-03-13|Baseline|2009-10-30|2009-10-30|Complete|Done|3|4|4|4|3|4|3.67|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1|||||||||Red||Child/Family: Lost contact with volunteer/agency|40.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28211|One Parent: Female|Unknown||No|Radio|Media|General Community||Match Support|M|Black||34|28202|Juris Doctorate (JD)|Single|Law: Lawyer||1|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501686648|36|0|1|501818631|31|0|1|500392214|2||-2||4|3|||-2||-2|55|1|||7446|3|||1|14832|-1|4|3|44
501725162|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2016-10-14|Baseline|2009-10-29|2009-10-29|Complete|Done|4|1|2|1|4|4|2.67|||||||||3|4|2|3|3|3|3|||||||||1|4|4|3||||||5|1|5|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|2|3.33||||||4|3|3.5|||||2|2|||||||||Green||Agency: Challenges with program/partnership|83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501724831|39|0|1|501833178|1|0|1|500394157|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|16143|-1|4|3|44
501375940|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-10|2010-04-06|Baseline|2009-11-12|2009-12-10|Complete|Done|4|2|4|2|3|4|3.17|||||||||2|4|4|3|4|3|3.33|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1|||||||||Green||Volunteer: Moved|3.8||1|1|1|1|M|Black||18|No|Mother|28215|One Parent: Female|Unknown||No||Service Organization|General Community||Match Support|M|White||33|28211|Bachelors Degree|Single|Business: Marketing|28213|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500009007|501376219|31|0|1|501857916|1|0|1|500410007|2||-2||4|1|||-2||-2|0|11|||7464|9|||1|17849|-1|4|3|44
501777213|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-15|2011-01-19|Baseline|2009-12-02|2009-12-15|Complete|Done|4|1|3|1|2|4|2.5|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||5|1|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|2|3.33||||||2|2|2|||||2|2|||||||||Green||Volunteer: Moved|13.1||2|2|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||37|28217|Bachelors Degree|Single|Unemployed||0|0|Yahoo!|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500011639|501777568|31|0|1|501897253|31|0|1|500417596|2||-2||4|1||500005291|-2||-2|0|10|||32|2|||1|21893|-1|4|3|44
501872495|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-14|2010-10-26|Baseline|2009-12-03|2009-12-10|Complete|Done|4|1|2|1|3|3|2.33|||||||||1|3|3|3|2|3|2.5|||||||||4|4|4|4||||||1|5|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red||Child/Family: Moved|10.4||1|1|1|1|M|Black||19|No|Non-Relative: Other|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|Some Other Race||37|28209|PHD|Single|Medical: Doctor, Provider||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500009007|501872868|31|0|1|501891059|41|0|1|500418064|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|22175|-1|4|3|44
501831955|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-11|2010-10-27|Baseline|2009-12-04|2009-12-11|Complete|Done|3|4|3|2|2|2|2.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1|||||||||Green||Child/Family: Feels incompatible with volunteer|10.5||1|1|1|1|M|White||16||Mother|28027|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||37|28025|High School Graduate|Divorced|Unknown||1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|501832323|1|0|1|501972975|1|0|1|500418296|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|22305|-1|4|3|44
501904094|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-15|2013-06-19|Baseline|2009-12-11|2010-01-12|Complete|Done|4|1|4|2|4|4|3.17|||||||||2|4|4|3|4|4|3.5|||||||||4|4|4|4||||||3|4|2|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red||Volunteer: Lost contact with child/agency|41.1||1|1|1|1|F|Black||16|No|Mother|28214|One Parent: Female|Unknown|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||56|28208|Some College|Single|Finance: Accountant|28203|19|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500004169|501904482|31|0|2|501342148|31|0|2|500420809|2||-2||4|3|||-2|500000294|-2|34|2|||7446|3|||1|23717|-1|4|3|44
501860404|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-21|2012-07-31|Baseline|2010-01-11|2010-01-21|Complete|Done|3|1|4|2|4|4|3|||||||||2|4|2||4|3||||||||||4|4|4|4||||||5|3|2|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|1|2.5|||||2|2|||||||||Green||Volunteer: Moved|30.3||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Enrollment|M|White||30|28202||Single|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501860777|31|31|1|501893096|1|0|1|500425993|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|26821|-1|4|3|44
501955313|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-29|2011-08-16|Baseline|2010-01-19|2010-01-29|Complete|Done|4|2|3|2|4|4|3.17|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||1|3|3|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|18.5||2|2|1|1|F|Black||16||Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28270||Single|Business: Clerical||10|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500010765|501955711|31|0|2|500915390|1|0|2|500427542|2||-2||4|1||500005291|-2||-2|0|10|||130|1|||1|27768|-1|4|3|44
501936316|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-28|2016-08-29|Baseline|2010-01-21|2010-01-28|Complete|Done|3|3|3|2|2|2|2.5|||||||||3|3||3|3|3||||||||||3|3|3|3||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child/Family: Lost contact with volunteer/agency|79||1|1|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||54|28203|||Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|501936714|31|0|1|501872326|1|0|1|500428557|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|28181|-1|4|3|44
501877268|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2011-10-13|Baseline|2010-01-22|2010-01-26|Complete|Done|4|3|4|4|3|4|3.67|||||||||2|3|2|2|1|3|2.17|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||2|2|||||||||Red||Child/Family: Lost contact with volunteer/agency|20.5||1|1|1|1|M|Black||19|No|Mother|28213|One Parent: Female|Unknown|Y|Yes|Radio|Media|General Community||Match Support|M|White||33|28269|||Construction||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011639|501877641|31|0|1|501942543|1|0|1|500429020|2||-2||4|3|||-2||-2|55|1|||7447|3|||1|28469|-1|4|3|44
501588821|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-10|2012-05-23|Baseline|2010-01-22|2010-02-10|Complete|Done|4|1|2|1|3|3|2.33|||||||||1|4|3|1|1|4|2.33|||||||||4|4|4|4||||||5|1|1|2|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|27.4||1|1|2|2|F|Black||16||Mother|28208|Two Mothers|Unknown||Yes||Self|General Community||Match Support|F|Black||34|28273|Masters Degree|Living w/ Significant Other|Consultant|28273|1|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501589141|31|0|2|501359582|31|0|2|500429105|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|28524|-1|4|3|44
501434147|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Baseline|2010-02-01|2010-03-31|Complete|Done|3|1|4|3|1|3|2.5|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4|5|2|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|||83.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||26|28215|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501434432|31|0|1|501926474|31|0|1|500441566|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|29966|-1|4|3|44
501716763|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-07|2016-11-11|Baseline|2010-02-02|2010-05-07|Complete|Done|1|1|1|1|1|1|1|||||||||2|1|2|2|3|2|2|||||||||3|3|3|3||||||2|3|2|2|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1|||||||||Red||Child/Family: Lost contact with volunteer/agency|78.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Amachi, Cabarrus County|Match Support|F|Black||39|28269||Single|Self-Employed, Entrepreneur|28027|7|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501716992|31|0|2|502112513|31|0|2|500449029|2||-2||4|3||500000294, 500016374|-2|500016374|-2|6854|8|||7458|9|||1|30228|-1|4|3|44
501957505|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-25|2012-03-31|Baseline|2010-02-03|2010-02-22|Complete|Done|4|1|1|1|3|4|2.33|||||||||2|3|4|3|3|3|3|||||||||4|3|4|3.67||||||5|2|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|3|3|||||1|1|||||||||Green|Amachi|Volunteer: Moved|25.1||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||55|28078|||Business: Marketing|28070|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501957903|31|0|1|501718938|1|0|1|500432245|2||-2||4|1|500000294||-2||-2|0|10|||7464|9|||1|30477|-1|4|3|44
501852702|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-25|2011-08-30|Baseline|2010-02-25|2010-06-25|Complete|Done|3|2|2|2|2|2|2.17|||||||||3|3|2|3|3|3|2.83|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||1|1|||||||||Red||Volunteer: Lost contact with child/agency|14.2||1|1|1|1|F|Black||19|No|Mother|28216|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||33|28205||Single|Consultant|28205|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501853073|31|0|2|501637271|1|0|2|500458675|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|33507|-1|4|3|44
502117432|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-03|2011-03-21|Baseline|2010-03-03|2010-03-03|Complete|Done|4|4|4|1|1|3|2.83|||||||||1|1|3|2|2|3|2|||||||||4|4|4|4||||||4|3|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|1|2.5|||||2|2|||||||||Green||Child/Family: Moved|12.6||1|1|4|4|F|Black||17|No|Father|28027|One Parent: Male|Unknown||Yes||BBBS Board/Staff|General Community||Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500011639|502117859|31|0|2|500189709|31|0|2|500438904|2||-2||4|1|||-2|500000294, 500016374|-2|0|13|||2230|7|||1|34304|-1|4|3|44
501877080|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-31|2010-09-02|Baseline|2010-03-10|2010-03-31|Complete|Done|1|4|4|2|4|4|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||1|1|||||||||Green||Volunteer: Feels incompatible with child/family|5.1||1|1|3|3|M|Black||17|No|Mother|28215|One Parent: Female|Unknown||Yes|Radio|Media|General Community||Enrollment|M|White||36|28202|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010765|501877453|31|0|1|501811850|1|0|1|500440340|2||-2||4|1|||-2||-2|55|1|||7464|9|||1|35176|-1|4|3|44
501741559|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-13|2011-10-13|Baseline|2010-03-16|2010-08-13|Complete|Done|3|3|3|4|3|3|3.17|||||||||3|3|3|3|2|3|2.83|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||4|2|3|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|14||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||32|28208|Bachelors Degree|Married|Tech: Production Line||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501741899|31|0|1|502213067|31|0|1|500464036|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|35898|-1|4|3|44
501919423|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-24|NaT|Baseline|2010-03-18|2010-03-24|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|3|3.5|||||1|1|||||||||Green|Project Big||83.7||1|1|1|1|M|Multi-race (Black & Hispanic)||17|No|Mother|28214|One Parent: Female|Unknown||No|TV|Media|General Community|Project Big|Match Support|M|White||34|28164|Masters Degree||Finance|28210|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501919819|38|0|1|502034798|1|0|1|500442066|2||500004641||2|1|500004640|500004640|-2||-2|56|1|||7464|9|||1|36152|-1|4|3|44
501765404|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-20|2013-08-29|Baseline|2010-03-22|2010-04-20|Complete|Done|3|3|3|1|4|3|2.83|||||||||2|3|3|2|3|3|2.67|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|3|2|3|1|3||||||||||4|3|4|3.67||||||4|3|3.5|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|40.3||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Multi-race (Black & White)||28|28262||Single|Student: College|28262|3|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501765751|31|0|1|501958658|36|0|1|500443642|2||-2||4|2|||-2||-2|0|10|||9221|5|||1|36416|-1|4|3|44
502076679|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2012-09-06|Baseline|2010-04-13|2010-04-30|Complete|Done|4|2|3|2|3|4|3|||||||||3|3||3|3|3||||||||||3|3|3|3||||||2|4|4|4|3.5|||||||4|4|4|4||4|4|||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red||Volunteer: Time constraint|28.3||1|1|1|1|M|Black||17|No|Mother|28273|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||37|28278|||Finance: Banking||0|0|AA Task Force|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502077103|31|0|1|502003579|1|0|1|500446859|2||-2||4|3|||-2||-2|0|4|||9228|10|||1|38100|-1|4|3|44
501938887|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2011-10-26|Baseline|2010-04-14|2010-04-30|Complete|Done|4|3|4|3|4|4|3.67|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Red||Child/Family: Lost contact with volunteer/agency|17.9||1|1|1|1|M|Black||18|No|Mother|28205|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|M|White||34|28205|||Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|501939285|31|0|1|502014005|1|0|1|500447313|2||-2||4|3|||-2||-2|0|8|||7496|10|||1|38283|-1|4|3|44
501877073|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2010-09-01|Baseline|2010-04-15|2010-04-30|Complete|Done|2|4|4|4|4|3|3.5|||||||||2|2|2|2|4|2|2.33|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||1|1|||||||||Yellow||Child/Family: Lost contact with volunteer/agency|4.1||1|1|2|2|M|Black||18|No|Mother|28215|One Parent: Female|Unknown||Yes|Radio|Media|General Community||Enrollment|M|Black||40|28215|Some College|Married|Transport: Driver||3|0|Michael Baisden|Media|Big|General Community||Match Support|277|60|598|500000170|500010765|501877446|31|0|1|502035292|31|0|1|500447499|2||-2||4|2|||-2||-2|55|1|||11146|1|||1|38363|-1|4|3|44
501990745|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-14|2012-08-29|Baseline|2010-04-19|2010-05-14|Complete|Done|2|2|3|1|1|2|1.83|||||||||3|3|3|3|4|3|3.17|||||||||3|3|3|3||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||1|1|||||||||Red||Child: Severity of challenges|27.5||1|1|1|1|M|Black||16||Mother|28269|One Parent: Female|Unknown||Yes||BBBS Board/Staff|General Community||Match Support|M|Black||35|28213||Married|Human Services: Youth Worker||0|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500011746|501991144|31|0|1|502098002|31|0|1|500447817|2||-2||4|3|||-2||-2|0|13|||4748|14|||1|38490|-1|4|3|44
501749652|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-01|2013-11-07|Baseline|2010-04-20|2010-09-01|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Moved|38.2||1|1|2|2|M|Black||18||Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|Black||52|28107|Some College|Divorced|Tech: Engineer|28262|3|0|Local Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500012459|501749994|31|0|1|501645507|31|0|1|500464305|2||-2||4|2|||-2||-2|0|10|||7437|1|||1|38597|-1|4|1|44
502088477|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-24|2010-08-24|Baseline|2010-05-05|2010-05-24|Complete|Done|3|3|3|3|3|3|3|||||||||2|3|3|2|2|3|2.5|||||||||3|2|2|2.33||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|2|2.5|||||1|1|||||||||Green||Child/Family: Moved|3||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Black||35|28210|||Personal Trainer/Coach||0|0|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500010355|502070907|31|0|1|502013648|31|0|1|500451408|2||500003586||4|1||500000294|-2|500000294|-2|0|10|||7464|9|||1|39523|-1|4|3|44
502083450|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-20|2011-08-26|Baseline|2010-05-05|2010-05-20|Complete|Done|4|4|4|4|3|4|3.83|||||||||4|2|3|2|4|3|3|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Amachi|Volunteer: Time constraint|15.2||2|2|1|1|M|Black||16|No|Mother|28027|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||44|28262||Divorced|Service: Restaurant|28027|0|10|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|502083874|31|0|1|502104415|31|0|1|500453680|2||500003586||4|1|500000294|500005291|-2||-2|7016|11|||7464|9|12|3|1|39542|-1|4|3|44
502114586|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2011-08-30|Baseline|2010-05-13|2010-08-27|Complete|Done|2|1|4|1|3|4|2.5|||||||||1|4|3|4|1|3|2.67|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||1|1|||||||||Green||Volunteer: Time constraint|12.1||1|1|1|1|M|Black||18|No|Mother|28211|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||RTBM|M|White||40|28277|Bachelors Degree|Married|Construction||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|502115013|31|0|1|502081755|1|0|1|500462278|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|40059|-1|4|3|44
502106926|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-25|2012-06-28|Baseline|2010-05-20|2010-05-25|Complete|Done|4|4|4|1|2|4|3.17|||||||||1|2|4|3|3|3|2.67|||||||||4|4|4|4||||||5|1|5|1|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red||Volunteer: Time constraint|25.1||2|2|1|1|M|Black||17|No|Mother|28031|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28031||Single|Govt||0|0|AA Task Force|Special Event|Big|General Community||Match Support|277|60|598|500000170|500011746|502107353|31|0|1|502072628|1|0|1|500453665|2||-2||4|3|||-2||-2|0|10|||11098|8|||1|40460|-1|4|3|44
502083495|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-26|2011-10-20|Baseline|2010-05-20|2010-05-26|Complete|Done|4|4|4|1|4|4|3.5|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red|Amachi|Volunteer: Lost contact with child/agency|16.8||1|1|2|2|M|Black||18|Yes|Mother|28025|One Parent: Female|Unknown||Yes||Service Organization|General Community|Amachi|Match Support|M|Black||52|28027||Married|Business: Human Resources|28273|0|0|Big Champions|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|502083919|31|0|1|502089653|31|0|1|500453681|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|11|||7461|12|||1|40468|-1|4|3|44
502102857|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-05|2010-10-28|Baseline|2010-05-20|2010-08-05|Complete|Done|4|4|3|1|4|4|3.33|||||||||3|4|3|3|1|4|3|||||||||4|4|2|3.33||||||4|4|5|1|3.5|||||||4|4|4|4|2|4|3|3.57||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Red||Volunteer: Unrealistic expectations|2.8|Y|2|2|1|1|M|Black||18|No|Mother|28278|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||63|28278|Some College|Married|Business: Engineer||25|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500009007|502103284|31|0|1|502240743|1|0|1|500463814|2||-2||4|3||500005291|-2|500000294|-2|0|4|||7464|9|||1|40474|-1|4|3|44
500185534|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-13|2012-12-20|Followup|2011-05-13|2011-06-28|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Family structure changed|79.3||1|1|3|5|M|Black||18||Mother|28204|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||63|28206|Some College|Married|Self-Employed, Entrepreneur|28206|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187159|31|0|1|500189461|31|0|1|500093294|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|81705||4|1|45
500185571|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-02|2015-07-14|Followup|2011-05-02|2011-05-16|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|4|2|2|3|2.67|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red||Child: Graduated|110.4||1|1|1|1|M|Black||19||Mother|28215|Other/Unknown|Unknown||No|Other|Faith Organization|General Community||Match Support|M|Black||49|28213|Bachelors Degree|Married|Finance: Banking|28288|4|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187198|31|0|1|500188438|31|0|1|500089543|2||-2||4|3|||-2||-2|5635|9|||7464|9|||1|81707||4|3|45
500185593|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-05|2011-04-27|Followup|2010-12-05|2011-02-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|64.7||1|1|2|2|M|Black||21||Mother|28262|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||34|28213|Bachelors Degree|Single|Finance: Banking|28202|0|2|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500187227|31|0|1|500234684|31|0|1|500062071|2||-2||4|2|||-2||-2|0|8|||7458|9|||1|81708||4|1|45
500185596|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-19|2011-05-05|Followup|2010-12-19|2011-03-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|64.5||1|1|1|1|M|Black||22||Mother|28205|Other/Unknown|Unknown||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|500187230|31|0|1|500310736|31|0|1|500068627|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81709||4|0|45
500185601|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-28|2015-07-23|Followup|2011-01-28|2011-02-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|89.8||2|2|1|1|M|Black||20||Mother|28210|Other/Unknown|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28078|High School Graduate|Single|Finance: Accountant|28202|0|4|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500187235|31|0|1|501082220|1|0|1|500236473|2||-2||4|1|||-2||-2|6854|8|||7458|9|||1|81710||4|1|45
500185624|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-28|2013-02-26|Followup|2010-06-28|2010-06-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Moved|68||1|1|1|1|M|Black||16|Yes|Mother|28213|Other/Unknown|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||61|28205||Married|Tech: Management||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|500187258|31|0|1|500923420|31|0|1|500182113|2||500003586||4|2|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|81711||4|1|45
500185628|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-09|2012-08-30|Followup|2010-08-09|2010-10-24|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|72.7||2|2|2|2|M|American Indian or Alaska Native||22||Mother|28031|Other/Unknown|Unknown||No||Neighbor/Friend|General Community||Match Support|M|White||51|28078|Bachelors Degree|Married|Business: Sales|28269|0|6|Igniting Breakfast|Special Event|Big|General Community|mentor2.0, mentor2.0 2015|RTBM|277|60|598|500000170|500008321|500187262|6|0|1|500190654|1|0|1|500117464|2||||4|3|||-2|500014505, 500015184|-2|0|8|||17266|8|||1|81712||4|0|45
500185630|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-26|2012-09-06|Followup|2010-09-26|2010-11-10|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Time constraints|71.4||3|3|2|2|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||39|28211|High School Graduate|Single|Finance: Banking|28208|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008629|500187264|31|0|2|500542491|31|0|2|500122710|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|81713||4|1|45
500185637|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-29|2014-12-11|Followup|2010-12-29|2011-02-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|107.4||1|1|2|2|M|Black||20||Mother|28206|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Black||55|28297|Masters Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500187271|31|0|1|500189284|31|0|1|500073080|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|81714||4|1|45
500185644|BBBS of Greater Charlotte|Main Office|C|Completed|2002-03-12|2011-06-17|Followup|2011-03-12|2011-05-27|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|111.2||1|1|1|1|M|Black||23||Mother|28269|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||46|28213|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008062|500187279|31|0|1|500188593|31|0|1|500036593|2||-2||4|3|||-2||-2|0|8|||7496|10|||1|81715||4|0|45
500185647|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-09|2013-10-31|Followup|2010-07-09|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|123.8||1|2|1|2|F|Black||21|Yes|Mother|28217|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||38|28269|Bachelors Degree|Married|Unknown|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187284|31|0|2|500188649|31|0|2|500038124|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|81716||4|1|45
500185675|BBBS of Greater Charlotte|Main Office|C|Completed|2003-06-04|2010-08-03|Followup|2010-06-04|2010-06-16|Complete|Done|4|3|3|3|4|4|3.5|||||||||2|3|3|2|3|3|2.67|||||||||4|4|4|4||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|2|1.5|||||2|2|||||||||Green||Child: Graduated|86||1|1|1|1|F|Black||24||Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||43|28278|Juris Doctorate (JD)|Single|Law: Lawyer|28205|0|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|500187557|31|0|2|500188632|31|0|2|500036632|2||-2||4|1|||-2||-2|0|10|||7459|10|||1|81717||4|3|45
500185678|BBBS of Greater Charlotte|Main Office|C|Completed|2003-02-23|2012-07-31|Followup|2011-02-23|2011-04-18|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|113.2||1|1|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28277|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500187309|31|0|1|500188619|31|0|1|500036619|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81718||4|1|45
500185706|BBBS of Greater Charlotte|Main Office|C|Completed|2000-07-28|2011-07-22|Followup|2010-07-28|2010-07-20|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Green||Child: Graduated|131.8||1|1|1|1|M|White||23||Mother|28226|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||46|28078|Bachelors Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500187480|1|0|1|500188657|1|0|1|500036657|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81720||4|3|45
500185721|BBBS of Greater Charlotte|Main Office|C|Completed|2003-12-03|2012-05-25|Followup|2010-12-03|2010-12-06|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|101.7||1|1|1|1|M|Black||22||Mother|28054|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||43|28207||Single|Unknown||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500187333|31|0|1|500188678|1|0|1|500036678|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81721||4|1|45
500185723|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-05|2015-06-25|Followup|2010-09-05|2010-11-20|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|81.6||2|2|1|1|M|Black||19||Mother|28214|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|M|Black||36|28214|Bachelors Degree|Single|Tech: Computer/Programmer|28147|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187335|31|0|1|501310677|31|0|1|500284133|2||-2||4|3|||-2||-2|6855|8|||7464|9|||1|81722||4|0|45
500185729|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-26|2012-09-05|Followup|2010-11-26|2011-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|57.3||2|2|2|2|M|Black||22||Relative: Other|28208|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||35|2109||Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500187496|31|0|1|500188672|1|0|1|500223221|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81723||4|1|45
500185734|BBBS of Greater Charlotte|Main Office|C|Completed|2003-10-15|2013-08-15|Followup|2010-10-15|2010-10-26|Complete|Done|3|3|2|3|3|3|2.83|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Red||Child: Graduated|118||1|1|1|1|F|Black||21||Mother|28203|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|White||45|28202|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187476|31|0|2|500188688|1|0|2|500036688|2||-2||4|3|||-2||-2|0|8|||7464|9|||1|81724||4|3|45
500185752|BBBS of Greater Charlotte|Main Office|C|Completed|2004-03-16|2012-10-17|Followup|2011-03-16|2011-05-24|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|103.1||1|2|1|2|M|Black||22|Yes|Mother|28227|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||51|28212|Some College|Single|Clergy||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500012459|500187343|31|0|1|500188744|31|0|1|500038128|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|81725||4|1|45
500185758|BBBS of Greater Charlotte|Main Office|C|Completed|2000-10-30|2011-06-17|Followup|2010-10-30|2011-01-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|127.5||1|1|1|1|F|Black||24||Mother|28205|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||46|28078|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008062|500187350|31|0|2|500188703|1|0|2|500036703|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81726||4|0|45
500185778|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-17|2016-06-23|Followup|2010-06-17|2010-06-30|Complete|Done|4|4|4|3|3|3|3.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||4|3|5|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|144.2||1|1|1|1|M|Black||18||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||42|27514||Married|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187368|31|0|1|500188776|1|0|1|500036776|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81727||4|3|45
500185781|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-13|2012-04-30|Followup|2011-02-13|2011-04-06|Complete|Late|3|2|3|2|3|3|2.67|||||||||2|3|3|2|2|3|2.5|||||||||4|3|3|3.33||||||3|2|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2|||||||||Red||Child: Graduated|50.5||2|2|2|2|M|Black||23||Mother|28262|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||34|28105||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013709|500187370|31|0|1|500188751|1|0|1|500244796|2||||4|3|||-2||-2|6854|8|||7464|9|||1|81728||4|3|45
500185815|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-17|2011-08-24|Followup|2010-12-17|2011-02-11|Blank|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|20.2||5|5|2|2|F|Black||21|No|Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||44|28211|Bachelors Degree|Single|Transport: Flight Attendant||10|0|Other|Service Organization|Big|General Site||Match Support|277|60|598|500000170|500001281|500187403|31|0|2|501356152|1|0|2|500419960|2||-2||4|1|||-2||-1|0|10|||7452|6|||1|81730||4|3|45
500185842|BBBS of Greater Charlotte|Main Office|C|Completed|2004-12-02|2012-02-08|Followup|2010-12-02|2011-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|86.2||1|1|1|1|M|Black||20||Mother|28206|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Site||Match Support|277|60|598|500000170|500008629|500187428|31|0|1|500188911|31|0|1|500036911|2||-2||4|1|||-2||-1|0|10|||7464|9|||1|81731||4|1|45
500185846|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-28|2014-10-23|Followup|2010-09-28|2010-11-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|120.8||1|2|1|2|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||65|28256|Bachelors Degree||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187437|31|0|2|500188764|31|0|2|500038142|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|81732||4|1|45
500185863|BBBS of Greater Charlotte|Main Office|C|Completed|2005-03-12|2014-05-15|Followup|2011-03-12|2011-03-18|Complete|Done|3|2|2|3|3|3|2.67|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|110.1||1|1|1|1|F|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||43|28202|Bachelors Degree|Married|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187435|31|0|2|500188915|1|0|2|500036915|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81735||4|3|45
500185865|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-15|2014-08-20|Followup|2010-12-15|2010-12-14|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow||Child/Family: Lost contact with volunteer/agency|68.1||2|2|2|2|F|Black||19||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187761|31|0|2|500189140|31|0|2|500326656|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|81736||4|3|45
500185897|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-05|2014-01-31|Followup|2011-02-05|2011-02-16|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|4|3.67||||||2|2|2|||||2|2|||||||||Red|Project Big|Child: Graduated|83.8||2|2|1|1|M|Black||21|No|Relative: Other|28208|Other Relative|Unknown||No||Self|General Community||Match Support|M|White||39|28277|Bachelors Degree|Single|Tech: Computer/Programmer||4|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500008321|500187458|31|0|1|500549520|1|0|1|500155451|2||500004641||4|3|500004640||-2||-2|0|10|||46|2|||1|81738||4|3|45
500185907|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2015-02-18|Followup|2010-10-29|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|99.7||2|3|1|1|F|Black||19|Yes|Mother|28262|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||48|28212||Single|Medical: Healthcare Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187470|31|0|2|500697782|31|0|2|500134557|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81739||4|1|45
500185972|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-01|2012-12-21|Followup|2010-09-01|2010-11-16|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|75.7||2|3|1|1|F|Black||22|Yes|Mother|28206|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|F|Black||38|28213|Bachelors Degree|Single|Education: Teacher|28202|2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187610|31|0|2|500492482|31|0|2|500120588|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81741||4|0|45
500186040|BBBS of Greater Charlotte|Main Office|C|Completed|2002-12-19|2011-06-17|Followup|2010-12-19|2011-03-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|101.9||1|1|1|1|F|Black||24|No|GrandMother|28208|Grandparents|Unknown||No||Self|General Community||Match Support|F|Black||48|28217|Bachelors Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008062|500187836|31|0|2|500188989|31|0|2|500036989|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81742||4|0|45
500186071|BBBS of Greater Charlotte|Main Office|C|Completed|2004-01-05|2014-04-30|Followup|2011-01-05|2011-02-28|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|123.8||1|1|1|1|M|White||21|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||40|28277|Masters Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187670|1|0|1|500189012|1|0|1|500037012|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81745||4|1|45
500186088|BBBS of Greater Charlotte|Main Office|C|Completed|2003-10-03|2011-10-26|Followup|2010-10-03|2010-12-18|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|96.8||1|1|1|1|M|Black||23|No|Mother|28203|Other/Unknown|Unknown||No||School|General Community||Match Support|M|White||44|28210|Bachelors Degree|Single|Finance: Banking|28211|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|277|60|598|500000170|500002335|500187606|31|0|1|500188966|1|0|1|500036966|2||-2||4|1|||-2||-1|0|4|||7496|10|||1|81746||4|0|45
500186092|BBBS of Greater Charlotte|Main Office|C|Completed|2000-06-20|2011-06-17|Followup|2010-06-20|2010-06-30|Complete|Done|3|3|4|4|4|4|3.67|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||2|5|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||1|2|1.5|||||2|2|||||||||Green||Child: Graduated|131.9||1|2|1|2|F|Black||23||Foster Parent|28203|Foster Home|Unknown||No||Self|General Community||Match Support|F|Black||47|28215|Bachelors Degree||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500187688|31|0|2|500189027|31|0|2|500038146|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81747||4|3|45
500186106|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-18|2015-08-13|Followup|2010-10-18|2010-12-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|93.8||2|2|1|1|F|Black||20||Mother|28217|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||35|28211|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187698|31|0|2|500778380|1|0|2|500202993|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|81748||4|1|45
500186107|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-22|2012-10-17|Followup|2010-06-22|2010-06-30|Complete|Done|4|1|4|2|3|2|2.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2|||||||||Green||Child: Graduated|75.9||2|2|1|1|M|Black||22||Mother|28206|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|Black||52|28210|Masters Degree|Married|Business: Mgt, Admin||0|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500012459|500187654|31|0|1|500392161|31|0|1|500102003|2||-2||4|1|||-2||-2|0|10|||2230|7|||1|81749||4|3|45
500186133|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-14|2016-06-28|Followup|2010-10-14|2010-10-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|140.5||1|1|1|1|M|White||18||Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||51|28262|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500187724|1|0|1|500188930|1|0|1|500036930|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|81750||4|1|45
500186141|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-02|2014-04-30|Followup|2011-04-02|2011-05-16|Complete|Done|4|3|4|1|4|4|3.33|||||||||2|4|4|3|4|3|3.33|||||||||4|4|4|4||||||4|3|4|2|3.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|72.9||3|3|1|1|F|Black||20|No|Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||45|28269|Bachelors Degree|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|500187731|31|0|2|501046739|31|0|2|500254296|2||-2||4|1|||-2|500000294|-2|0|10|||46|2|||1|81751||4|3|45
500186174|BBBS of Greater Charlotte|Main Office|C|Completed|2005-07-28|2012-10-31|Followup|2010-07-28|2010-10-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|87.1||2|2|2|2|F|Black||18||Mother|28208|One Parent: Female|Unknown||No||Self|General Community||Enrollment|F|Black||48|29715|Some College|Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500187758|31|0|2|500189225|31|0|2|500038037|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|81752||4|0|45
500186190|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-13|2014-08-20|Followup|2010-10-13|2010-11-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|118.2||1|1|2|2|F|Black||20||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187761|31|0|2|500189140|31|0|2|500037140|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|81754||4|1|45
500186191|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-21|2011-05-24|Followup|2010-10-21|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|79||1|2|1|2|F|Black||18|Yes|Mother|28213|One Parent: Female|Unknown|Y|No|Brochure|Media|General Community|Amachi|Match Support|F|Black||58|28269|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500187792|31|0|2|500189141|31|0|2|500038186|2||500003586||4|1|500000294|500000294|-2|500000294|-2|51|1|||2238|7|||1|81755||4|1|45
500186206|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-24|2013-09-30|Followup|2011-02-24|2011-03-15|Complete|Done|3|2|4|1|4|4|3|||||||||3|3|4|1|3|4|3|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|3|3|4|3|3.57||||||||||3|2|1|2||||||3|1|2|||||2|2|||||||||Red||Child/Family: Moved|103.2||1|1|1|1|M|Black||20||GrandMother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||44|28214|PHD|Married|Medical: Doctor, Provider||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187812|31|0|1|500189157|31|0|1|500037157|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|81756||4|3|45
500186247|BBBS of Greater Charlotte|Main Office|C|Completed|2005-06-30|2012-09-26|Followup|2010-06-30|2010-07-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|86.9||1|1|2|2|M|Black||21||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|M|Black||39|28269|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Site|mentor2.0 2014|RTBM|277|60|598|500000170|500008321|500187842|31|0|1|500189197|31|0|1|500037197|2||-2||4|3|||-2|500014506|-1|0|10|||7464|9|||1|81759||4|1|45
500186248|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-09|2011-07-29|Followup|2011-03-09|2011-03-18|Complete|Done|3|2|2|2|3|3|2.5|||||||||4|3|4|4|3|4|3.67|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|3|3|3.71||||||||||3|3|3|3||||||4|2|3|||||2|2|||||||||Yellow||Volunteer: Lost contact with child/agency|28.6||3|3|1|1|F|Black||17||Mother|28214|Other/Unknown|Unknown||No||Self|General Community||Enrollment|F|Black||40|28216||Single|Finance: Banking||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500001281|500187843|31|0|2|501470065|31|0|2|500340015|2||-2||4|2|||-2||-2|0|10|||7462|13|||1|81760||4|3|45
500186260|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-29|2015-12-17|Followup|2010-10-29|2011-01-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|133.6||3|3|1|1|M|Black||19|No|Mother|28025|One Parent: Female|Unknown||No||Self|General Site||Match Support|M|Black||42|28025|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|500187857|31|0|1|500189139|31|0|1|500037139|2||-2||4|2|||-1||-2|0|10|||7464|9|||1|81761||4|0|45
500186277|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2014-07-16|Followup|2010-07-08|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Moved|60.3||3|4|2|3|F|Black||18||Mother|28206|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||39|28210|Bachelors Degree|Married|Business: Sales||8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500187876|31|0|2|500188587|1|0|2|500373187|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|81762||4|1|45
500186291|BBBS of Greater Charlotte|Main Office|C|Completed|2004-11-30|2011-07-29|Followup|2010-11-30|2010-12-13|Complete|Done|3|3|4|3|4|3|3.33|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2|||||||||Green||Child: Graduated|79.9||1|1|2|2|F|Black||23||Foster Parent|28269|Other Relative|Unknown|Y|No||Self|General Community||Match Support|F|Black||49|28269|Bachelors Degree|Divorced|Finance|28282|0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500008629|500219859|31|0|2|500189241|31|0|2|500037241|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|81763||4|3|45
500186325|BBBS of Greater Charlotte|Main Office|C|Completed|2003-11-19|2012-11-29|Followup|2010-11-19|2011-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|108.4||2|2|2|3|M|Black||22||Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28202|Bachelors Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187951|31|0|1|500189265|1|0|1|500047102|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81765||4|1|45
500186327|BBBS of Greater Charlotte|Main Office|C|Completed|2003-01-11|2012-11-30|Followup|2011-01-11|2011-02-28|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|118.6||1|1|1|1|M|Black||22||Mother|28208|One Parent: Female|Unknown|Y|No||School|General Community||Match Support|M|White||63|28211|Some College|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|500187974|31|0|1|500189289|1|0|1|500037301|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|81766||4|1|45
500186336|BBBS of Greater Charlotte|Main Office|C|Completed|2002-09-20|2011-07-28|Followup|2010-09-20|2010-12-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|106.2||1|1|1|1|M|Black||24||Mother|28208|One Parent: Female|Unknown|Y|No||School|General Community||Match Support|M|White||57|28277|Bachelors Degree|Married|Business: Sales||0|0|Billboard|Media|Big|General Community||Match Support|277|60|598|500000170|500011184|500187974|31|0|1|500189301|1|0|1|500037314|2||-2||4|1|||-2||-2|0|4|||125|1|||1|81769||4|0|45
500186352|BBBS of Greater Charlotte|Main Office|C|Completed|2002-07-29|2014-01-02|Followup|2010-07-29|2010-07-30|Complete|Done|3|3|3|3|3|3|3|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||5|5|3|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|137.2||4|4|2|2|M|Black||21||Mother|28212|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|White||45|28226|Masters Degree|Married|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500187945|31|0|1|500189280|1|0|1|500037290|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|81770||4|3|45
500186355|BBBS of Greater Charlotte|Main Office|C|Completed|2005-05-02|2011-08-24|Followup|2011-05-02|2011-04-20|Complete|Done|3|3|3|3|3|3|3|||||||||2|3|3|3|3|3|2.83|||||||||4|3|3|3.33||||||3|3|3|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|75.7||2|3|1|2|M|Some Other Race||23||Father|28208|One Parent: Male|Unknown||No||Neighbor/Friend|General Community||Match Support|M|White||40|28205|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500187961|41|0|1|500189814|1|0|1|500038144|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|81771||4|3|45
500186374|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-28|2012-01-10|Followup|2010-06-28|2010-09-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|66.4||2|2|1|1|F|Black||22||Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||55|28269|High School Graduate|Single|Business: Human Resources|28202|5|0|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008629|500187968|31|0|2|500419439|31|0|2|500102160|2||-2||4|2|||-2||-2|0|10|||6247|12|||1|81772||4|0|45
500186385|BBBS of Greater Charlotte|Main Office|C|Completed|2003-02-11|2013-01-09|Followup|2011-02-11|2011-03-18|Complete|Done|3|2|4|3|4|4|3.33|||||||||2|4|4|4|3|4|3.5|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|118.9||1|1|1|1|M|Black||22||Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||43|28269|Bachelors Degree|Single|Finance: Accountant|28262|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|500187967|31|0|1|500189269|31|0|1|500037278|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|81773||4|3|45
500186428|BBBS of Greater Charlotte|Main Office|C|Completed|2005-10-03|2013-09-30|Followup|2010-10-03|2010-10-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|95.9||1|2|2|3|M|Black||21||Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||40|28211|Bachelors Degree|Single|Unknown||0|0|Brochure|Media|Big|General Community||Match Support|277|60|598|500000170|500004169|500187986|31|0|1|500189441|1|0|1|500044683|2||-2||4|1|||-2||-2|0|10|||127|1|||1|81774||4|1|45
500186435|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-23|2015-08-20|Followup|2010-07-23|2010-08-20|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|144.9||1|1|1|1|M|Black||20||Mother|28216|One Parent: Female|Unknown||No|Brochure|Media|General Community||Match Support|M|White||45|28226|Bachelors Degree|Married|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187988|31|0|1|500189358|1|0|1|500037395|2||-2||4|1|||-2||-2|51|1|||7496|10|||1|81776||4|3|45
500186436|BBBS of Greater Charlotte|Main Office|C|Completed|2003-08-07|2010-11-12|Followup|2010-08-07|2010-09-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|87.2||1|1|1|1|M|Black||24||Mother|28216|One Parent: Female|Unknown||No|Brochure|Media|General Community||Match Support|M|Black||42|28213|Bachelors Degree|Married|Finance: Banking||0|0|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500187988|31|0|1|500189444|31|0|1|500037500|2||-2||4|1|||-2||-2|51|1|||7458|9|||1|81777||4|1|45
500186570|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-05|2011-04-05|Followup|2010-10-05|2010-10-28|Complete|Done|3|4|4|4|2|4|3.5|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|4|3|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2|||||||||Yellow||Child/Family: Lost contact with volunteer/agency|78||2|2|1|1|F|Black||19||Mother|28269|Other/Unknown|Unknown||No||Self|General Community||RTBM|F|Black||37|28213|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|500188168|31|0|2|500189615|31|0|2|500037719|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|81780||4|3|45
500186615|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-09|2011-09-29|Followup|2011-05-09|2011-06-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|64.7||2|2|1|1|F|Black||22||Mother|28278|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||39|28269|PHD|Single|Medical: Doctor, Provider||0|8|Other|BBBS Board/Staff|Big|General Site|Amachi, mentor2.0 2014|Enrollment|277|60|598|500000170|500008629|500188023|31|0|2|500403330|31|0|2|500093132|2||-2||4|1|500000294|500000294|-2|500000294, 500014506|-1|0|10|||7671|13|||1|81781||4|1|45
500186636|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-27|2011-08-16|Followup|2010-06-27|2010-09-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|61.6||2|2|1|1|F|Black||20||Mother|28208|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|F|Black||48|28277|Masters Degree|Married|Business: Sales||0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188037|31|0|2|500452589|31|0|2|500102306|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|81782||4|0|45
500186645|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-03|2016-01-06|Followup|2010-06-03|2010-07-02|Complete|Done|4|2|3|2|3|3|2.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|Amachi|Child: Graduated|139.1||1|1|1|1|M|Black||18|Yes|Mother|28208|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28256|High School Graduate|Married|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500018987|500188043|31|0|1|500189545|31|0|2|500037636|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81783||4|3|45
500186646|BBBS of Greater Charlotte|Main Office|C|Completed|2005-10-20|2013-09-23|Followup|2010-10-20|2010-12-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|95.1||3|3|3|3|F|Some Other Race||21||Mother|28217|Other/Unknown|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||39|28216|Some College||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500188044|41|0|2|500189263|31|0|2|500047741|2||-2||4|2|||-2||-2|0|8|||7464|9|||1|81784||4|1|45
500186665|BBBS of Greater Charlotte|Main Office|C|Completed|2004-07-20|2013-02-28|Followup|2010-07-20|2010-10-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|103.3||1|1|1|1|M|Black||21||Mother|28202|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|Black||40|28207||Single|Medical: Nurse||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500188050|31|0|1|500189566|31|0|1|500037664|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|81785||4|0|45
500186675|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-23|2013-08-29|Followup|2010-08-23|2010-10-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|72.2||4|4|1|1|F|Black||20|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||38|28221||Single|Human Services: Youth Worker||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188055|31|0|2|500865601|31|0|2|500185332|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81786||4|1|45
500186682|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2015-07-22|Followup|2010-07-20|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|96.1||3|4|1|1|M|Black||20|Yes|Mother|28227|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|M|Black||57|28262||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|500887363|31|0|1|500184396|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81788||4|1|45
500186692|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-11|2012-06-30|Followup|2010-09-11|2010-11-26|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|33.6||7|8|1|1|F|Black||19|No|Mother|28270|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|White||50|28270|Some College|Single|Finance: Banking|28217|1|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500188059|31|0|2|501582415|1|0|2|500381441|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|81789||4|0|45
500186702|BBBS of Greater Charlotte|Main Office|C|Completed|2004-04-28|2014-11-25|Followup|2011-04-28|2011-04-20|Complete|Done|3|3|3|3|3|3|3|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|3|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||2|2|2|||||2|2|||||||||Green|Amachi|Child: Graduated|126.9||1|2|1|2|F|Black||20|Yes|GrandMother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||57|28212|Some College|Married|Unknown||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|RTBM|277|60|598|500000170|500017732|500188150|31|0|2|500189528|31|0|2|500038225|2||500003586||4|1|500000294|500000294|-2|500015184|-1|0|10|||7462|13|||1|81790||4|3|45
500186760|BBBS of Greater Charlotte|Main Office|C|Completed|2004-08-09|2010-10-26|Followup|2010-08-09|2010-09-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Family structure changed|74.5||1|1|1|1|M|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||No|TV|Media|General Community|Amachi|Match Support|M|Black||43|28269|Bachelors Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188154|31|0|1|500189588|31|0|1|500037690|2||500003586||4|1|500000294|500000294|-2|500000294|-2|56|1|||2238|7|||1|81792||4|1|45
500186765|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-05|2013-08-15|Followup|2010-09-05|2010-09-03|Complete|Done|2|3|3|3|3|3|2.83|||||||||3|3|4|3|3|4|3.33|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|107.3||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||46|28078|Masters Degree|Widowed|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500004169|500188083|31|0|2|500189359|31|0|2|500037396|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81793||4|3|45
500186788|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-21|2011-06-17|Followup|2010-09-21|2010-10-01|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|80.8||1|1|2|2|M|Black||24||Mother|28208|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||47|28204||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|500188098|31|0|1|500189605|1|0|1|500037707|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|81794||4|1|45
500186798|BBBS of Greater Charlotte|Main Office|C|Completed|2005-03-30|2015-10-20|Followup|2011-03-30|2011-04-05|Complete|Done|3|2|4|4|3|3|3.17|||||||||2|3|3|3|3|3|2.83|||||||||4|3|3|3.33||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child/Family: Time constraints|126.7||1|2|1|2|F|Multi-Race (None of the above)||19|No|Father|28208|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||45|28226|Bachelors Degree||Business: Human Resources||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500187961|7|0|2|500189825|1|0|2|500038158|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81795||4|3|45
500186800|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-06|2012-07-25|Followup|2010-10-06|2010-12-21|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|93.6||1|1|3|3|F|Black||22||Mother|28216|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|500188103|31|0|2|500189320|31|0|2|500037337|2||-2||4|1|||-2|500016374|-2|0|4|||7464|9|||1|81796||4|0|45
500186813|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-05|2011-04-21|Followup|2010-10-05|2010-12-20|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|78.5||1|1|2|2|M|Black||22||Mother|28273|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||46|28214|Bachelors Degree|Single|Finance: Economist|28217|14|0|Brochure|Media|Big|General Community||Match Support|277|60|598|500000170|500009007|500188094|31|0|1|500189600|31|0|1|500037702|2||-2||4|3|||-2||-2|0|8|||127|1|||1|81797||4|0|45
500186830|BBBS of Greater Charlotte|Main Office|C|Completed|2005-07-14|2011-06-17|Followup|2010-07-14|2010-07-09|Complete|Done|3|3|3|2|3|3|2.83|||||||||3|3|3|3|2|3|2.83|||||||||3|3|3|3||||||4|4|5|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|71.1||1|1|2|2|M|Black||22||Mother|28208|Other/Unknown|Unknown||No||Self|General Community||Match Support|M|White||47|28204||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|500188106|31|0|1|500189605|1|0|1|500037708|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|81798||4|3|45
500186853|BBBS of Greater Charlotte|Main Office|C|Completed|2004-11-04|2012-01-27|Followup|2010-11-04|2010-10-29|Complete|Done|4|2|3|3|4|4|3.33|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2|||||||||Yellow||Child/Family: Lost contact with volunteer/agency|86.7||1|1|1|1|M|Black||21||Mother|28210|Other/Unknown|Unknown||No||Self|General Community||Match Support|M|Black||36|28203|Bachelors Degree||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500264223|31|0|1|500189632|31|0|1|500037741|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|81799||4|3|45
500186905|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-10|2015-11-04|Followup|2011-02-10|2011-03-31|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Graduated|128.8||1|1|1|1|F|Black||19|Yes|Mother|28205|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|F|Black||50|28215|Some College|Single|Finance: Banking||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188151|31|0|2|500189677|31|0|2|500037790|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|81801||4|1|45
500186923|BBBS of Greater Charlotte|Main Office|C|Completed|2004-08-31|2011-05-24|Followup|2010-08-31|2010-11-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Family structure changed|80.7||1|2|1|2|M|Black||19|Yes|Mother|28215|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||54|28216|Bachelors Degree|Single|Unknown|28205|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188131|31|0|1|500189696|31|0|1|500038078|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6855|8|||2238|7|||1|81803||4|0|45
500186925|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-24|2011-12-21|Followup|2011-02-24|2011-03-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|81.8||1|1|1|1|M|Black||22|Yes|Mother|28205|One Parent: Female|Unknown|Y|No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||59|28269|Masters Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188151|31|0|1|500189697|31|0|1|500037810|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|81804||4|1|45
500186926|BBBS of Greater Charlotte|Main Office|C|Completed|2004-08-30|2011-12-21|Followup|2010-08-30|2010-11-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|87.7||1|1|1|1|M|Some Other Race||23|Yes|Mother|28213|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||60|28277|Bachelors Degree|Married|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188133|41|0|1|500189699|31|0|1|500037812|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|81805||4|0|45
500186938|BBBS of Greater Charlotte|Main Office|C|Completed|2004-08-24|2011-12-21|Followup|2010-08-24|2010-10-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Lost contact with child/agency|87.9||1|1|1|1|F|Black||21||Mother|28215|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||40|28217|Bachelors Degree|Single|Finance: Accountant|28277|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188131|31|0|2|500189708|31|0|2|500037821|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|81806||4|1|45
500186943|BBBS of Greater Charlotte|Main Office|C|Completed|2005-10-26|2011-08-16|Followup|2010-10-26|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|69.7||2|2|1|1|F|Black||21||Mother|28269|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||40|28297|||Human Services: Social Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188139|31|0|2|500224697|31|0|2|500048942|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|81807||4|1|45
500186946|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-20|2012-08-23|Followup|2010-06-20|2010-09-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Lost contact with child/agency|62.1||2|2|1|1|F|Black||19|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||36|28262||Single|Education: Teacher||4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188139|31|0|2|500865596|31|0|2|500181565|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81808||4|0|45
500186952|BBBS of Greater Charlotte|Main Office|C|Active|2004-07-15|NaT|Followup|2010-07-15|2010-07-26|Complete|Done|4|4|4|2|3|4|3.5|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|5|3|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|4|2.5|||||2|2|||||||||Green|Amachi||152||1|1|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||73|28203||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|500188132|31|0|2|500189723|1|0|2|500037836|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81810||4|3|45
500186953|BBBS of Greater Charlotte|Main Office|C|Completed|2004-05-25|2012-08-09|Followup|2010-05-25|2010-08-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.5||1|1|2|2|M|Black||18|Yes|GrandMother|28214|Other Relative|Unknown||No||Self|General Community|Amachi|Match Support|M|White||45|28207||Single|Unknown|28209|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188126|31|0|1|500189724|1|0|1|500037838|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81811||4|0|45
500186955|BBBS of Greater Charlotte|Main Office|C|Completed|2004-05-21|2014-02-19|Followup|2011-05-21|2011-06-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Lost contact with child/agency|117||1|1|1|1|F|Black||18|No|Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||55|28226|||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|2|500189726|1|0|2|500037840|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81812||4|1|45
500186956|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-21|2015-03-04|Followup|2010-06-21|2010-09-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|128.4||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28203|Bachelors Degree|Married|Law: Lawyer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|500189727|1|0|1|500037841|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81813||4|0|45
500186960|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-31|2013-08-15|Followup|2010-07-31|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Time constraint|72.5||2|2|1|1|M|White||19|Yes|Mother|28227|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||40|28105|Some College|Married|Military|28112|11|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188147|1|0|1|500738970|1|0|1|500186719|2||500003586||4|3|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|81814||4|1|45
500186990|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-17|2014-02-28|Followup|2011-02-17|2011-03-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|60.4||2|2|3|3|M|Black||19|Yes|Mother|28269|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||51|28269|Bachelors Degree|Married|Unknown|28202|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500188170|31|0|1|500189496|31|0|1|500339895|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81816||4|1|45
500187075|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-21|2014-01-16|Followup|2010-09-21|2010-09-16|Complete|Done|3|4|4|4|3|3|3.5|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|3|4|3|4|4|3.71||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|111.8||1|1|6|6|F|Black||21||Mother|28205|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||38|28209|Bachelors Degree|Single|Human Services: Non-Profit||0|0|Recruitment Event|Self|Big|General Site||Match Support|277|60|598|500000170|500012459|500188223|31|0|2|500189550|1|0|2|500037643|2||-2||4|1|||-2||-1|0|10|||7458|9|||1|81819||4|3|45
500187077|BBBS of Greater Charlotte|Main Office|C|Completed|2005-05-31|2013-04-02|Followup|2010-05-31|2010-06-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|94.1||2|2|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||41|28210|Bachelors Degree|Married|Medical: Pharmacist||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500188224|31|0|1|500189824|1|0|2|500037944|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81820||4|1|45
500187090|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-04|2013-08-29|Followup|2010-10-04|2010-12-19|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|82.8||2|2|3|3|F|Black||20||Mother|28216|Two Parent|Unknown||No||School|General Community||Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|500188103|31|0|2|500189320|31|0|2|500125754|2||-2||4|1|||-2|500016374|-2|0|4|||7464|9|||1|81821||4|0|45
500191327|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-07|2012-09-05|Followup|2010-12-07|2011-01-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Family structure changed|69||2|2|1|1|M|Black||19||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28212||Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008629|500191330|31|0|1|500547393|31|0|1|500144146|2||-2||4|1|||-2||-2|0|10|||46|2|||1|81823||4|1|45
500191820|BBBS of Greater Charlotte|Main Office|C|Completed|2005-09-30|2013-08-29|Followup|2010-09-30|2010-11-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|94.9|Y|2|2|2|2|M|Black||19||Mother|28227||Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||72|28214||Married|Retired||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500191823|31|0|1|500191501|31|0|1|500044434|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|81825||4|1|45
500234359|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-17|2011-06-17|Followup|2010-12-17|2011-03-03|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|66||1|1|1|1|M|Black||22||Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||33|28269|Bachelors Degree|Single|Finance: Banking|28262|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008062|500234368|31|0|1|500251451|31|0|1|500068942|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|81834||4|0|45
500237080|BBBS of Greater Charlotte|Main Office|C|Completed|2005-11-16|2012-01-12|Followup|2010-11-16|2011-01-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Severity of challenges|73.9||1|1|2|2|M|Black||18|Yes|Mother|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||40|28269||Married|Business: Marketing||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500237089|31|0|1|500220237|31|0|1|500057623|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81835||4|1|45
500252077|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-24|2016-01-20|Followup|2010-11-24|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|85.8||3|3|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Tech: Computer/Programmer||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501750989|31|0|1|501365749|1|0|1|500317108|2||500003586||4|3|500000294|500000294|-2||-2|7295|11|||46|2|||1|81838||4|1|45
500261295|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-21|2017-03-09|Followup|2010-12-21|2011-02-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|134.6||1|1|1|1|M|White||20||Mother|28104|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||60|28270|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500261310|1|0|1|500188435|1|0|1|500073081|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81839||4|1|45
500267459|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-19|2013-02-27|Followup|2010-09-19|2010-10-05|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|77.3||1|1|1|1|M|Black||16||Mother|28203|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28202|Bachelors Degree|Single|Finance: Accountant||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|500187395|31|0|1|500464544|1|0|1|500121193|2||-2||4|3|||-2||-2|0|10|||46|2|||1|81841||4|1|45
500271303|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-30|2015-08-03|Followup|2011-04-30|2011-06-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|75.1||2|2|1|1|F|Black||17|Yes|Mother|28227|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|White||31|28204|Bachelors Degree|Single|Business: Engineer|28269|0|2|TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500271368|31|0|2|501291358|1|0|2|500354049|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||130|1|||1|81842||4|1|45
500293140|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-05|2011-02-09|Followup|2010-12-05|2011-01-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|62.2||2|2|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28205|Some College|Single|Business: Clerical||0|10|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008629|500191330|31|0|1|500191399|1|0|1|500062178|2||-2||4|1||500005291|-2||-2|0|10|||46|2|||1|81843||4|1|45
500337327|BBBS of Greater Charlotte|Main Office|C|Active|2006-12-14|NaT|Followup|2010-12-14|2010-12-10|Complete|Done|4|1|4|1|3|3|2.67|||||||||2|3|3|3|2|3|2.67|||||||||3|3|3|3||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|||123||2|3|4|5|M|Black||16||GrandMother|28208|Grandparents|Unknown||No||School|General Site||Match Support|M|Black||49|28217|Associate Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site||Match Support|277|60|598|500000170|500017732|500251937|31|0|1|500189300|31|0|1|500148262|2||-2||2|1|||-1||-1|0|4|||7464|9|||1|81845||4|3|45
500340183|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-18|2013-08-30|Followup|2010-12-18|2010-12-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|44.4||3|3|1|1|M|Black||17|No|Relative: Other|28208|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction||0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|500340317|31|0|1|501933993|1|0|1|500419988|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|81847||4|1|45
500342076|BBBS of Greater Charlotte|Main Office|C|Completed|2006-02-14|2012-02-28|Followup|2011-02-14|2011-03-19|Complete|Done|3|1|3|1|3|3|2.33|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2|||||||||Green||Child: Graduated|72.4||1|1|1|1|M|Black||23||Mother|28216|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||35|28207|Bachelors Degree|Single|Business: Marketing||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|500342211|31|0|1|500188562|1|0|1|500080816|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|81848||4|3|45
500361200|BBBS of Greater Charlotte|Main Office|C|Active|2006-03-21|NaT|Followup|2011-03-21|2011-06-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Cabarrus County||131.8||2|2|1|1|F|White||17|No|Mother|28027|Two Parent|Unknown||No||Relative|General Community|Cabarrus County|Match Support|F|White||32|28115|Bachelors Degree|Single|Human Services: Social Worker||0|0|other|College Partner|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500361450|1|0|2|500368628|1|0|2|500085591|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|3|||7670|5|||1|81850||4|0|45
500363209|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-24|2010-12-30|Followup|2010-05-24|2010-08-08|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|55.2||1|1|1|1|F|Multi-Race (None of the above)||16|Yes|Mother|28025|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||57|28262||Married|Finance: Banking||0|9|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188099|7|0|2|500371073|31|0|2|500099752|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81851||4|0|45
500363212|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-24|2012-11-27|Followup|2010-05-24|2010-08-08|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Moved|66.2||2|2|1|1|F|Multi-Race (None of the above)||16||Mother|28025|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||34|28211|Associate Degree|Living w/ Significant Other|Business: Clerical|28211|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188099|7|0|2|500797130|1|0|2|500176231|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|81852||4|0|45
500378354|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-01|NaT|Followup|2011-05-01|2011-05-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||106.5||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$40,000 to $44,999||No|Big|Neighbor/Friend|General Community||Match Support|M|White||36|28270|Juris Doctorate (JD)|Married|Law: Lawyer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500378596|31|0|1|501181060|1|0|1|500264206|2||-2||2|1|||-2||-2|6854|8|||46|2|||1|81854||4|1|45
500382177|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-18|2015-08-25|Followup|2010-09-18|2010-10-20|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|4|4|4|3|3|3.5|||||||||4|4|4|4||||||3|3|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|2|3|2.67||||||4|4|4|||||2|2|||||||||Yellow||Volunteer: Lost contact with child/agency|107.2||1|1|2|2|M|Black||16||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||43|28215|Bachelors Degree|Single|Finance: Banking|28262|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|500382427|31|0|1|500188566|31|0|1|500122093|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|81857||4|3|45
500383915|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-20|2012-08-30|Followup|2010-06-20|2010-09-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|50.3||2|2|2|2|F|Black||20||GrandMother|28205|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||64|28269||Married|Finance: Economist||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|500384165|31|0|2|500540512|31|0|2|500274279|2||-2||4|1|||-2||-2|6855|8|||7464|9|||1|81858||4|0|45
500383923|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-30|2012-08-30|Followup|2010-08-30|2010-11-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|72||1|1|2|2|M|Black||18||GrandMother|28205|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||66|28269||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500384165|31|0|1|500540549|31|0|1|500118470|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|81859||4|0|45
500392419|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-06|2013-08-29|Followup|2011-03-06|2011-03-10|Complete|Done|4|4|4|2|3|3|3.33|||||||||4|3|4|3|4|3|3.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|4|3.5|||||2|2|||||||||Yellow||Child/Family: Moved|77.8||2|2|1|1|F|Black||21||Father|28105|One Parent: Male|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||32|28277||Single|Business: Sales||0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500392669|31|0|2|500746900|1|0|2|500162012|2||-2||4|2|||-2||-2|6855|8|||7464|9|||1|81860||4|3|45
500392858|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-15|2010-12-30|Followup|2010-12-15|2010-12-09|Complete|Done|3|3|4|3|4|3|3.33|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2|||||||||Green||Child/Family: Moved|24.5||3|3|2|2|M|Black||20||Aunt|28215|One Parent: Female|Unknown||No||Therapist/Counselor|General Community||Match Support|M|White||43|28227|High School Graduate|Married|Clergy||10|0|General|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|500393108|31|0|1|501064465|1|0|1|500326650|2||-2||4|1|||-2|500000294|-2|0|5|||6450|12|||1|81861||4|3|45
500392860|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-18|2011-07-29|Followup|2011-01-18|2011-02-16|Complete|Done|3|4|3|2|3|3|3|||||||||2|3|3|2|2|3|2.5||||||||||3|3|||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|42.3||2|2|2|2|M|Black||18||Aunt|28215|One Parent: Female|Unknown||No||Therapist/Counselor|General Community||Match Support|M|White||43|28227|High School Graduate|Married|Clergy||10|0|General|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|500393108|31|0|1|501064465|1|0|1|500236600|2||-2||4|1|||-2|500000294|-2|0|5|||6450|12|||1|81862||4|3|45
500393176|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-07|2012-06-21|Followup|2010-06-07|2010-08-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|72.5||1|1|1|1|F|Black||22||Relative: Other|28216|Other Relative|Unknown||No||Relative|General Community|Amachi|Match Support|F|Black||35|28213||Single|Tech: Engineer||2|0|Bellafonte Presbyter|Faith Organization|Big|General Site|Amachi|Enrollment|277|60|598|500000170|500013781|500187361|31|0|2|500415570|31|0|2|500101074|2||500003586||4|1|500000294|500000294|-2|500000294|-1|0|3|||2238|7|||1|81863||4|0|45
500395038|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-01|2015-02-20|Followup|2010-08-01|2010-08-03|Complete|Done|4|4|4|2|3|4|3.5|||||||||3|3|3|4|4|4|3.5|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Child: Graduated|102.7||1|1|1|1|M|White||20||Mother|28226|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|M|White||39|28211|Masters Degree|Married|Law: Lawyer|28204|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500395288|1|0|1|500392006|1|0|1|500104016|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|81864||4|3|45
500398853|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-16|2011-07-08|Followup|2011-02-16|2011-05-03|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|2010-2012 OJJDP JJI|Child: Lost interest|52.7||1|1|1|1|M|Black||21|No|Mother|28083|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||40|28269|Masters Degree|Married|Govt: Mgmt/Admin|28202|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500002335|500399103|31|0|1|500795095|31|0|1|500155431|2||-2||4|1|500005291||-2||-2|0|10|||2238|7|||1|81865||4|0|45
500399525|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-15|2012-08-29|Followup|2010-06-15|2010-08-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Agency: Challenges with program/partnership|74.5||1|1|1|1|F|Black||19||Mother|28214|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||46|28217|Some College|Single|Finance: Accountant|28208|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500399775|31|0|2|500416787|31|0|2|500099891|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|81866||4|0|45
500399844|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-20|2017-02-24|Followup|2010-08-20|2010-11-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|114.2||1|2|1|2|F|Black||16||Mother|28208|One Parent: Female|Unknown||No||School|General Site||Match Support|F|White||35|28210|Bachelors Degree|Single|Business: Mgt, Admin|29715|0|0|Radio|Media|Big|General Site||Match Support|277|60|598|500000170|500008321|500400094|31|0|2|500188569|1|0|2|500190707|2||-2||4|3|||-1||-1|0|4|||131|1|||1|81867||4|0|45
500402676|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-27|2012-02-29|Followup|2010-06-27|2010-09-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Graduated|68.1||1|1|1|1|M|White||24|||28211|One Parent: Female|Unknown||No||Therapist/Counselor|General Community|Amachi|Match Support|M|White||36|28208|Bachelors Degree|Single|Business: Mgt, Admin|28203|2|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500402926|1|0|1|500339569|1|0|1|500102368|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|5|||2238|7|||1|81869||4|0|45
500402978|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-29|2012-05-08|Followup|2010-06-29|2010-09-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Time constraints|70.3||1|1|1|1|M|White||22||Mother|28211|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||33|28203|Bachelors Degree|Single|Business: Sales|27609|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500402926|1|0|1|500414710|1|0|1|500103314|2||-2||4|2|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|81870||4|0|45
500402982|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-29|2011-05-24|Followup|2010-06-29|2010-09-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Moved|58.8||1|1|1|1|M|White||18||Mother|28211|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||37|28212||Single|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500402926|1|0|1|500467614|1|0|1|500103313|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|81871||4|0|45
500408135|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-25|2015-01-30|Followup|2010-05-25|2010-08-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|104.2||1|1|4|4|F|Black||19|Yes|Mother|28083|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500008321|500408385|31|0|2|500189709|31|0|2|500099932|2||500003586||4|1|500000294|500000294|-2|500000294, 500016374|-2|6854|8|||2230|7|||1|81872||4|0|45
500417281|BBBS of Greater Charlotte|Main Office|C|Completed|2006-07-31|2013-01-31|Followup|2010-07-31|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|78.1|Y|1|1|1|1|F|White||16||Mother|28211|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||48|28211|Masters Degree|Married|Finance: Banking|28202|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500402926|1|0|2|500349297|1|0|1|500112798|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|81876||4|1|45
500417525|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-17|2012-11-30|Followup|2011-01-17|2011-04-03|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Volunteer: Time constraint|70.4||1|1|1|1|M|Black||18||Mother|28208|One Parent: Female|Unknown||No|TV|Media|General Community|Project Big|Match Support|M|White||37|28202|||Medical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500417775|31|0|1|500755435|1|0|1|500151964|2||500004641||4|1|500004640|500004640|-2||-2|56|1|||46|2|||1|81877||4|0|45
500418050|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-12|2012-11-28|Followup|2011-05-12|2011-06-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|78.6||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||34|28273|High School Graduate|Single|Transport: Driver|28216|0|10|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188055|31|0|1|500417272|31|0|1|500093386|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81878||4|1|45
500432759|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-26|2010-09-29|Followup|2010-05-26|2010-08-10|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|52.1||1|1|1|1|F|Black||22||Mother|28205|One Parent: Female|Unknown||No||Faith Organization|General Community||Match Support|F|Black||37|28216|Bachelors Degree|Single|Human Services: Non-Profit|28205|2|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500433090|31|0|2|500415680|31|0|2|500099996|2||-2||4|2|||-2||-2|0|9|||7464|9|||1|81880||4|0|45
500433644|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-04|2011-11-30|Followup|2011-02-04|2011-02-16|Complete|Done|4|1|1|1|3|4|2.33|||||||||1|1|1|1|1|4|1.5|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||1|1|4|4|4|4|3|3||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Red||Volunteer: Time constraint|21.8||2|2|1|1|M|Black||17||Mother|28269|One Parent: Female|Unknown||No||Relative|General Community||Enrollment|M|Black||60|28078|Bachelors Degree|Married|Tech: Computer/Programmer|28202|25|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500433894|31|0|1|501882367|31|0|1|500430294|2||-2||4|3|||-2||-2|0|3|||7464|9|||1|81882||4|3|45
500463808|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-15|2010-11-02|Followup|2010-08-15|2010-09-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|50.6||1|1|1|1|M|Black||23||Mother|28269|One Parent: Female|$50,000 to $59,999||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28269|Juris Doctorate (JD)|Single|Law: Lawyer||0|8|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500001281|500464059|31|0|1|500498479|31|0|1|500117634|2||-2||4|2|||-2||-2|34|2|||6450|12|||1|81883||4|1|45
500465506|BBBS of Greater Charlotte|Main Office|C|Active|2006-08-21|NaT|Followup|2010-08-21|2010-10-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi||126.8||1|1|1|1|M|Black||16|Yes|Mother|28262|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||54|28226|Bachelors Degree|Married|Arts, Entertainment, Sports||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500496966|1|0|1|500118121|2||500003586||2|2|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|81884||4|1|45
500465511|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-21|2013-10-31|Followup|2010-08-21|2010-10-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Graduated|86.3||1|1|1|1|M|Black||21|Yes|Mother|28262|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|M|White||54|28210|Masters Degree|Married|Finance: Accountant||0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500527675|1|0|1|500118120|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|4|||2230|7|||1|81885||4|1|45
500465521|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-21|2012-05-31|Followup|2010-08-21|2010-10-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|69.3||1|1|1|1|F|Black||23|Yes|Mother|28262|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|F|White||42|28209|Masters Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|2|500542558|1|0|2|500118432|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|81886||4|1|45
500472874|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-06|2011-07-29|Followup|2010-08-06|2010-10-21|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|35.7||2|2|1|1|F|Black||20|No|Mother|28262|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||32|28262|Masters Degree|Single|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500008062|500473122|31|0|2|501179381|31|0|2|500278853|2||-2||4|3|||-2||-2|0|10|||46|2|||1|81887||4|0|45
500474486|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-23|2015-08-18|Followup|2010-08-23|2010-08-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|107.8||1|1|1|1|M|Black||20||Mother|28214|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||38|28209|Bachelors Degree|Single|Construction|28247|0|2|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500474735|31|0|1|500491064|31|0|1|500118168|2||-2||4|3|||-2||-2|34|2|||7447|3|||1|81888||4|1|45
500474841|BBBS of Greater Charlotte|Main Office|C|Completed|2006-11-18|2012-01-17|Followup|2010-11-18|2011-01-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|62||1|1|2|2|F|Black||15||Mother|28208|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Multi-Race (None of the above)||52|28227|Bachelors Degree|Single|Education: Admin||4|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500013709|500474737|31|0|2|500370830|7|0|2|500133665|2||-2||4|2|||-2||-2|34|2|||46|2|||1|81889||4|1|45
500477277|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2011-05-25|Followup|2010-10-29|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|54.8||1|1|1|1|F|Black||17||Mother|28213|One Parent: Female|Less than $10,000||No||Service Organization|General Community||Match Support|F|Black||47|28027|Bachelors Degree|Single|Retail: Sales|28145|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500003657|500477524|31|0|2|500491044|31|0|2|500134558|2||500003586||4|1|500000294||-2||-2|0|11|||2238|7|||1|81890||4|1|45
500478936|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-14|2013-11-11|Followup|2010-07-14|2010-07-26|Complete|Done|3|4|4|4|3|3|3.5|||||||||4|4|3|4|4|3|3.67|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2|||||||||Green||Child: Graduated|63.9||1|1|3|3|M|Black||21|No|Mother|28078|One Parent: Female|$25,000 to $29,999||No||Neighbor/Friend|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|500479187|31|0|1|501284751|31|0|1|500275964|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|8|||132|8|||1|81891||4|3|45
500480596|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-13|2014-01-16|Followup|2010-09-13|2010-11-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|88.1||1|1|1|1|M|Black||21|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Married|Business: Sales|28203|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500480847|31|0|1|500491267|1|0|1|500120915|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|81892||4|1|45
500483980|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-01|2014-03-24|Followup|2010-09-01|2010-09-02|Complete|Done|3|2|3|3|3|3|2.83|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||5|3|3|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|90.7||1|1|2|2|M|Black||21||Mother|28227|One Parent: Female|$10,000 to $14,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||71|28270||Single|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500484231|31|0|1|500423426|31|0|1|500120592|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|81893||4|3|45
500496598|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-23|NaT|Followup|2010-10-23|2011-01-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi, Cabarrus County||100.7||2|2|1|1|M|White||15|Yes|Mother|28083|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi, Cabarrus County|Match Support|M|White||35|28083|Masters Degree|Single|Business: Mgt, Admin|28027|2|3|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500496849|1|0|1|501383928|1|0|1|500299090|2||500003586||2|2|500000294, 500016374|500000294, 500016374|-2|500016374|-2|34|2|||7464|9|||1|81894||4|0|45
500539341|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-24|2012-01-27|Followup|2010-09-24|2010-09-14|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|4|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Amachi|Child: Family structure changed|64.1||1|1|2|2|M|White||19|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||44|28205||Single|Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|500539592|1|0|1|500191356|1|0|1|500123020|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|81895||4|3|45
500540847|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-02|2011-05-24|Followup|2010-07-02|2010-09-16|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Moved|46.7||2|2|1|1|F|Black||16|Yes|Mother|28208|One Parent: Female|$20,000 to $24,999|Y|No||Service Organization|General Community|Amachi|Match Support|F|Black||41|28216|||Finance: Accountant||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500003657|500541089|31|0|2|500866129|31|0|2|500181618|2||500003586||4|1|500000294|500000294|-2||-2|0|11|||2238|7|||1|81898||4|0|45
500544934|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-17|2011-03-23|Followup|2010-06-17|2010-07-07|Complete|Done|4|3|4|2|3|2|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2|||||||||Yellow||Volunteer: Infraction of match rules/agency policies|33.1||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|$15,000 to $19,999|Y|No||Neighbor/Friend|General Community||Match Support|F|Black||67|28215||Married|Education: Teacher||0|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500010765|500545186|31|0|2|501213248|31|0|2|500269480|2||-2||4|2|||-2||-2|0|8|||2230|7|||1|81899||4|3|45
500545326|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2016-09-02|Followup|2010-10-29|2011-01-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|118.1|Y|1|1|1|1|M|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|Black||55|28214||Married|Clergy||12|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|1|500697845|31|0|1|500134545|2||-2||4|3|||-2||-2|0|10|||2238|7|||1|81900||4|0|45
500545328|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-02|2016-09-30|Followup|2010-07-02|2010-07-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|99||3|3|1|1|F|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|F|Black||43|28208|Masters Degree|Single|Business: Sales|28078|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|2|501033808|31|0|2|500274449|2||-2||4|1|||-2||-2|0|10|||46|2|||1|81901||4|1|45
500546821|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-21|2015-09-15|Followup|2011-02-21|2011-05-08|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|102.8||1|1|3|3|M|Black||20|No|Mother|28083|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||52|28025||Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500012459|500547073|31|0|1|500790181|31|0|1|500159910|2||-2||4|1|||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|81902||4|0|45
500566159|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-23|2012-03-12|Followup|2011-01-23|2011-04-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|49.6||2|2|1|1|F|Black||16||Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Enrollment|F|White||35|28207|||Business: Clerical||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|500565754|31|0|2|500966678|1|0|2|500230690|2||-2||4|2|||-2||-2|34|2|||46|2|||1|81904||4|0|45
500575861|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-22|2011-06-17|Followup|2010-07-22|2010-10-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|34.8||2|2|1|1|F|Black||23||Mother|28208|One Parent: Female|$10,000 to $14,999|Y|No||Neighbor/Friend|General Community||Match Support|F|White||37|28209|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008062|500576113|31|0|2|501202981|1|0|2|500274108|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|81912||4|0|45
500577339|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-16|2011-07-08|Followup|2011-04-16|2011-07-01|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|26.7||1|1|1|1|M|Black||20|No|Mother|28083|Two Parent|Unknown||No||Self|General Community||Match Support|M|White||37|28075|Some College|Married|Military||11|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500002335|500577557|31|0|1|501634485|1|0|1|500353354|2||-2||4|1|||-2||-2|0|10|||7446|3|||1|81913||4|0|45
500636603|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-21|2011-06-17|Followup|2011-03-21|2011-06-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|50.9||2|4|1|1|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|White||38|28226|Bachelors Degree|Married|Homemaker||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008062|500636863|31|0|2|500842825|1|0|2|500168014|2||-2||4|3|||-2||-2|0|8|||7671|13|||1|81915||4|0|45
500636617|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-10|2013-08-20|Followup|2011-01-10|2011-02-08|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|79.3||2|2|1|1|M|Black||17||Mother|28269|One Parent: Female|$20,000 to $24,999|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28262||Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500636863|31|0|1|500756919|31|0|1|500151137|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|81916||4|1|45
500705925|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-23|2011-03-22|Followup|2010-07-23|2010-09-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Moved|44||1|1|2|2|M|Black||23||Relative: Other|28269|Other Relative|$60,000 to $74,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|Black||48|28269||Divorced|Tech: Engineer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|500706192|31|0|1|500908500|31|0|1|500182939|2||-2||4|2|||-2||-2|34|2|||7496|10|||1|81923||4|1|45
500713145|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-30|2010-12-30|Followup|2010-08-30|2010-11-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|40||1|1|1|1|M|Black||21|Yes|GrandMother|28227|One Parent: Female|Less than $10,000|Y|No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||48|28227||Married|Military||21|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500713412|31|0|1|500932892|31|0|1|500187379|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|81926||4|0|45
500713817|BBBS of Greater Charlotte|Main Office|C|Active|2009-10-30|NaT|Followup|2010-10-30|2010-11-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||88.5||2|2|1|1|M|Black||16||Mother|28216|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28078|||Medical: Pharmacist|28210|10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|500714084|31|0|1|501834795|1|0|1|500396466|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|81927||4|1|45
500717519|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-08|2013-08-29|Followup|2010-12-08|2010-12-09|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|4|4|4|4|3|3.67|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2|||||||||Yellow||Child: Lost interest|80.7||1|1|2|2|M|Black||20||Mother|28205|One Parent: Female|$20,000 to $24,999|Y|No||School|General Community||Match Support|M|Black||37|28269|Bachelors Degree|Married|Education: Admin||0|0|Yahoo!|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|500717786|31|0|1|500188838|31|0|1|500145722|2||-2||4|2|||-2||-2|0|4|||32|2|||1|81928||4|3|45
500722500|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-20|2011-10-26|Followup|2010-06-20|2010-09-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|52.2||2|2|1|1|F|White||20||Mother|28027||Unknown||No||Service Organization|General Community||Match Support|F|White||34|28083|Bachelors Degree|Single|Education: Teacher Asst/Aid|28147|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|500722767|1|0|2|500830633|1|0|2|500180184|2||-2||4|1|||-2||-2|0|11|||7464|9|||1|81929||4|0|45
500724632|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-07|NaT|Followup|2011-03-07|2011-05-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||120.3||1|1|1|1|F|Black||17||Mother|28213|One Parent: Female|Less than $10,000|Y|No||School|General Community||Match Support|F|Black||32|28214|Bachelors Degree|Married|Architect|28270|0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|500724899|31|0|2|500803551|31|0|2|500164708|2||-2||2|1|||-2||-2|0|4|||46|2|||1|81930||4|0|45
500726828|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-14|2011-09-12|Followup|2011-05-14|2011-07-29|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Feels incompatible with child/family|52||1|1|3|3|M|Black||22||Mother|28027|One Parent: Female|$40,000 to $44,999||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||49|28027|Bachelors Degree|Married|Transport: Driver|28208|6|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|277|60|598|500000170|500002335|500187529|31|0|1|500863980|31|0|1|500173102|2||-2||4|1|||-2|500014505, 500014506|-1|34|2|||7671|13|||1|81931||4|0|45
500727291|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-17|2016-07-29|Followup|2011-05-17|2011-05-12|Complete|Done|3|2|3|2|3|3|2.67|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|110.4||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|Black||46|28269|||Human Services: Non-Profit||0|0|BBBS National Site|Web Link|Big|General Community|VOL - Adjudicated, VOL - Cultural Comp, VOL - PreMatch|Match Support|277|60|598|500000170|500008321|500727558|31|0|1|500857838|31|0|1|500176403|2||-2||4|1|||-2|500007913, 500007920, 500011311|-2|0|10|||46|2|||1|81932||4|3|45
500728622|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-16|2012-05-23|Followup|2010-08-16|2010-10-01|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|57.2||1|2|1|2|M|Black||18|No|Mother|28205|One Parent: Female|Unknown||No||School|General Site||Match Support|M|Black||78|28216||Married|Retired||20|0|Other|BBBS Board/Staff|Big|General Site||Match Support|277|60|598|500000170|500008629|500730811|31|0|1|500546003|31|0|1|500188249|2||-2||4|2|||-1||-1|0|4|||7671|13|||1|81933||4|1|45
500730385|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-15|2011-06-17|Followup|2011-03-15|2011-05-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|51.1||1|1|1|1|F|Black||18||Mother|28217|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|F|Black||38|28217|Bachelors Degree|Single|Finance: Banking|29715|5|0|Recruitment Event|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008062|500730652|31|0|2|500761242|31|0|2|500166676|2||-2||4|3|||-2||-2|0|10|||7460|12|||1|81934||4|0|45
500730544|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-21|2011-04-08|Followup|2010-06-21|2010-09-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|45.6||1|2|1|2|F|Black||21|No|Mother|28205|One Parent: Female|$25,000 to $29,999||Yes||School|General Site||Match Support|F|American Indian or Alaska Native||65|28270|Bachelors Degree|Married|Business: Mgt, Admin||5|0|Coworker|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500008629|500730811|31|0|2|500569158|6|0|2|500181810|2||-2||4|1|||-1||-1|0|4|||7447|3|||1|81935||4|0|45
500732462|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-18|2012-02-28|Followup|2010-07-18|2010-07-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|55.4||1|1|1|1|F|Black||22||Mother|28205|One Parent: Female|$30,000 to $34,999|Y|No||School|General Community||Match Support|F|Black||40|28269|Masters Degree|Single|Education: Admin|28223|1|9|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500732729|31|0|2|500878773|31|0|2|500184327|2||-2||4|1|||-2||-2|0|4|||7458|9|||1|81936||4|1|45
500732858|BBBS of Greater Charlotte|Main Office|C|Completed|2006-11-28|2011-04-29|Followup|2010-11-28|2011-02-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|53||1|1|1|1|M|Black||18|No|Mother|28203|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28212|Bachelors Degree|Single|Business: Marketing|28202|1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500733125|31|0|1|500344509|1|0|1|500142645|2||-2||4|1||500005291|-2||-2|0|10|||7464|9|||1|81937||4|0|45
500733695|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-26|2015-03-03|Followup|2010-12-26|2011-02-08|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.2||1|1|1|1|F|Black||19|Yes|GrandMother|28217|Grandparents|Less than $10,000|Y|No|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||34|28210|Bachelors Degree|Married|Finance: Accountant|28202|0|2|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500733962|31|0|2|500307108|1|0|2|500150172|2||500003586||4|3|500000294|500000294|-2||-2|7294|13|||2238|7|||1|81938||4|1|45
500740293|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2010-06-12|2010-06-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Lost interest|85||1|1|1|1|M|Black||19||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|Black||39|28216||Single|Transport: Pilot||3|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500876177|31|0|1|500179697|2||-2||4|2|||-2||-2|0|5|||6450|12|||1|81941||4|1|45
500740295|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2010-06-12|2010-06-30|Complete|Done|3|4|4|2|4|4|3.5|||||||||4|3|4|4|4|4|3.83|||||||||4|4|3|3.67||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Yellow||Volunteer: Feels incompatible with child/family|85||1|1|1|1|M|Black||18||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|White||55|28216|Bachelors Degree|Divorced|Tech: Engineer||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500794907|1|0|1|500179696|2||-2||4|2|||-2||-2|0|5|||46|2|||1|81942||4|3|45
500740296|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-25|2011-09-21|Followup|2010-06-25|2010-06-30|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|1|4|4|4|4|3.5|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Yellow||Volunteer: Lost contact with child/agency|50.9||2|2|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Therapist/Counselor|General Community||Match Support|F|Black||33|28269|Bachelors Degree|Single|Human Services: Non-Profit||0|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|2|500928282|31|0|2|500181834|2||-2||4|2|||-2||-2|0|5|||7671|13|||1|81943||4|3|45
500741571|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-15|2012-01-10|Followup|2010-08-15|2010-10-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|52.9||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Some Other Race||31|28262|||Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500002335|500724899|31|0|1|500938541|41|0|1|500187546|2||-2||4|1|||-2||-2|0|10|||46|2|||1|81944||4|0|45
500747371|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-31|2011-06-17|Followup|2010-12-31|2011-03-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|29.5||3|3|1|1|F|Black||20|No|Mother|28213|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||34|28025|Some College|Married|Business: Marketing|28262|11|0|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008062|500747638|31|0|2|501279505|1|0|2|500329319|2||-2||4|2|||-2|500000294|-2|0|4|||7464|9|||1|81945||4|0|45
500752612|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-17|2011-06-17|Followup|2010-08-17|2010-11-01|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|46||1|1|1|1|F|Black||20||Mother|28205|Foster Home|Unknown||No||Self|General Community||Match Support|F|White||33|28207||Divorced|Consultant||5|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500008062|500752880|31|0|2|500915297|1|0|2|500186913|2||-2||4|1|||-2||-2|0|10|||130|1|||1|81946||4|0|45
500764136|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-10|2012-08-23|Followup|2011-02-10|2011-03-31|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|30.4||3|3|1|1|M|Black||22|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community|Amachi|Match Support|M|White||32|28210|Some College|Single|Business: Mgt, Admin|28206|8|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500764404|31|0|1|501915488|1|0|1|500428501|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|81950||4|1|45
500764138|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-07|2013-02-21|Followup|2011-02-07|2011-03-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|72.5||2|2|1|1|M|Black||17|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community|Amachi|Match Support|M|Black||33|28214||Single|Tech: Research/Design||1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500764404|31|0|1|500696779|31|0|1|500154924|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81951||4|1|45
500764773|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-06|2011-06-17|Followup|2011-01-06|2011-03-23|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|41.3||2|2|1|1|F|Black||22||Mother|28212|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||36|28205|Bachelors Degree|Single|Medical: Nurse||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008062|500765039|31|0|2|501091276|1|0|2|500235607|2||-2||4|3|||-2||-2|0|10|||46|2|||1|81952||4|0|45
500765381|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-26|2015-10-20|Followup|2011-02-26|2011-03-11|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|1|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Moved|79.7||1|1|1|1|M|Black||16|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|10019|Bachelors Degree|Single|Business: Marketing|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500739190|31|0|1|501579025|1|0|1|500342803|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81953||4|3|45
500767208|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-03-24|Followup|2010-07-10|2010-07-16|Complete|Done|4|3|3|3|4|4|3.5|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green|Project Big|Child: Graduated|68.4||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|Black||32|28216|Masters Degree|Single|Human Services|28215|0|7|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Enrollment|277|60|598|500000170|500017732|500767473|31|0|2|501341042|31|0|2|500276669|2||500004641||4|1|500004640||-2|500014506|-1|0|10|||7671|13|||1|81954||4|3|45
500771298|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-02|2011-10-26|Followup|2010-11-02|2010-10-29|Complete|Done|4|3|3|2|2|4|3|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Time constraint|47.8||1|1|1|1|M|Black||19||Mother|28105|One Parent: Female|$35,000 to $39,999||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28110|||Finance: Banking||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|500771566|31|0|1|500953236|31|0|1|500206613|2||-2||4|2|||-2||-2|34|2|||46|2|||1|81956||4|3|45
500771746|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2016-06-15|Followup|2010-05-29|2010-08-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Child: Graduated|84.6||3|4|1|2|F|Black||19||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||37|28012|Some College|Married|Finance: Banking|28208|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500772014|31|0|2|500996153|1|0|2|500366437|2||500004641||4|1|500004640||-2||-2|0|4|||7464|9|||1|81957||4|0|45
500781988|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-16|2013-09-04|Followup|2011-02-16|2011-05-03|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|78.6||1|1|1|1|M|White||21||Mother|28027||Unknown||No||Self|General Community||Match Support|M|White||71|28083|Some College|Married|Business: Mgt, Admin|28027|13|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500002335|500782256|1|0|1|500773716|1|0|1|500160560|2||-2||4|1|||-2||-2|0|10|||46|2|||1|81960||4|0|45
500783100|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-08-29|Followup|2011-04-30|2011-05-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|112||1|1|1|1|M|Black||16||Mother|28206|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||36|28203|||Retail: Sales|28226|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|500783368|31|0|1|500777047|1|0|1|500174449|2||-2||4|2|||-2||-2|0|10|||46|2|||1|81961||4|1|45
500791567|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-31|2013-04-11|Followup|2011-01-31|2011-04-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|74.3||1|1|2|2|M|Multi-Race (None of the above)||18|No|Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|M|Black||32|28215||Married|Finance: Banking||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|500187654|7|0|1|500578720|31|0|1|500155823|2||-2||4|2|||-2||-2|0|10|||7447|3|||1|81964||4|0|45
500795704|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-30|2011-06-01|Followup|2011-01-30|2011-04-16|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Lost interest|52||1|1|1|1|F|Multi-Race (None of the above)||23|Yes|Mother|28081|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||42|28075||Single|Medical: Pharmacist|28025|7|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|500766037|7|0|2|500723270|31|0|2|500154833|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81966||4|0|45
500796255|BBBS of Greater Charlotte|Main Office|C|Active|2010-01-20|NaT|Followup|2011-01-20|2011-02-16|Complete|Done|2|1|2|1|4|2|2|||||||||2|2|3|4|2|4|2.83|||||||||4|4|4|4||||||3|2|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|||85.8||3|3|1|1|M|White||18|No|Mother|28031|One Parent: Male|$20,000 to $24,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||60|28269|||Medical: Admin|28207|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500796529|1|0|1|501846438|1|0|1|500424314|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|81967||4|3|45
500799303|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-27|2016-08-19|Followup|2011-03-27|2011-06-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|112.8||1|1|1|1|M|White||19|No|Mother|28081|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||46|28202||Single|Business: Sales||0|4|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500799571|1|0|1|500798390|1|0|1|500167062|2||-2||4|3||500016374|-2|500016374|-2|34|2|||7464|9|||1|81969||4|0|45
500801567|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-26|2013-12-12|Followup|2010-10-26|2010-12-01|Complete|Done|4|4|4|3|3|3|3.5|||||||||3|4|4|2|3|3|3.17|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|49.5||2|2|1|1|M|Black||20||Mother|28213|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||62|28078|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500801835|31|0|1|501834907|1|0|1|500391790|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81970||4|3|45
500806676|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-25|2010-10-26|Followup|2010-06-25|2010-07-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|40||1|1|1|1|M|Black||24||Mother|28269|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|Black||39|28213|Some College|Single|Military|28213|13|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500009007|500806944|31|0|1|500878893|31|0|1|500181682|2||-2||4|2|||-2||-2|0|10|||131|1|||1|81971||4|1|45
500809082|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-01|2012-03-13|Followup|2010-06-01|2010-07-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|57.4||1|1|1|1|M|Black||23||Mother|28210|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|White||34|28203|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||RTBM|277|60|598|500000170|500011746|500809351|31|0|1|500878459|1|0|1|500178590|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|81972||4|1|45
500814240|BBBS of Greater Charlotte|Main Office|C|Active|2008-04-24|NaT|Followup|2011-04-24|2011-06-30|Complete|Late|3|2|3|2|3|3|2.67|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|3|3|3|3|3.43||||||||||3|4|3|3.33||||||3|3|3|||||2|2|||||||||Green|Amachi||106.7||1|1|1|1|M|Black||18|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||46|28215|Bachelors Degree|Single|Business: Mgt, Admin|28226|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500814509|31|0|1|500981509|31|0|1|500248568|2||500003586||2|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|81974||4|3|45
500824037|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-15|NaT|Followup|2011-03-15|2011-05-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||120||1|1|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|F|White||34|28210|Bachelors Degree|Single|Education: Teacher|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500824306|31|0|2|500789337|1|0|2|500165956|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|81975||4|0|45
500826592|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-08|2016-10-18|Followup|2010-10-08|2010-11-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|84.3||3|3|1|1|F|Black||20|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|F|White||33|28277|Bachelors Degree|Living w/ Significant Other|Unknown|28209|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|2|501314246|1|0|2|500382768|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|81978||4|1|45
500826594|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-21|2016-06-15|Followup|2010-08-21|2010-10-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|105.8||1|1|1|1|M|Black||18|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Some Other Race||36|28209|||Business: Sales||0|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|1|500920342|41|0|1|500185735|2||-2||4|1|||-2||-2|0|5|||6450|12|||1|81979||4|1|45
500826596|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-07|2011-04-06|Followup|2010-08-07|2010-09-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|19.9||3|3|1|1|M|Black||17|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Black||35|28226|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500826861|31|0|1|501799403|31|0|1|500375650|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|81980||4|1|45
500835156|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2016-11-10|Followup|2010-07-10|2010-07-27|Complete|Done|2|3|4|3|4|4|3.33|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child/Family: Lost contact with volunteer/agency|100||1|2|1|2|M|Black||17||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Multi-Race (None of the above)||38|29710|Bachelors Degree|Single|Architect||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500835425|31|0|1|500466903|7|0|1|500277232|2||-2||4|1|||-2||-2|0|4|||46|2|||1|81982||4|3|45
500838847|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-15|2011-06-09|Followup|2010-06-15|2010-08-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|23.8||2|2|1|1|M|Black||19|No|Mother|28278|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community||Match Support|M|Black||37|28226|||Finance: Accountant|28110|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500839116|31|0|1|501647679|31|0|1|500364921|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81983||4|0|45
500843860|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-14|2011-03-31|Followup|2010-12-14|2011-02-28|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Moved|27.5||2|2|1|1|M|Black||22|Yes|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|No|TV|Media|General Community||Match Support|M|White||33|28202|Bachelors Degree|Single|Finance: Banking|28255|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500003657|500844129|31|0|1|501340550|1|0|1|500320896|2||500003586||4|1|500000294||-2||-2|56|1|||46|2|||1|81984||4|0|45
500843863|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-21|2016-06-17|Followup|2011-02-21|2011-03-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Changed workplace/school partnership|99.8||2|2|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|No|TV|Media|General Community|Amachi|Match Support|F|Black||32|28269|Bachelors Degree|Single|Business: Marketing|28273|0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500844129|31|0|2|501078655|31|0|2|500241388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|56|1|||2238|7|||1|81985||4|1|45
500847570|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-07|2011-08-16|Followup|2011-05-07|2011-06-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|51.3||2|2|1|1|F|Black||16|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||53|28216||Married|Business: Clerical||4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188056|31|0|2|500848661|31|0|2|500174103|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81986||4|1|45
500849042|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-14|2010-12-21|Followup|2010-11-14|2010-12-10|Complete|Done|4|1|4|2|4|4|3.17|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||1|1|1|||||2|2|||||||||Green||Child/Family: Moved|25.2||2|3|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||No||Service Organization|General Community||Match Support|F|Black||33|28202|Bachelors Degree|Divorced|Finance: Accountant||0|4|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500001281|500849311|31|0|2|501379402|31|0|2|500314655|2||-2||4|1|||-2||-2|0|11|||7446|3|||1|81987||4|3|45
500850236|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-04|2013-09-16|Followup|2011-04-04|2011-04-05|Complete|Done|4|2|4|1|4|4|3.17|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green||Child: Graduated|77.4||1|1|2|2|M|Black||21|No|Mother|28205|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|Black||37|28262|Bachelors Degree|Single|Real Estate: Realtor||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500850505|31|0|1|500189198|31|0|1|500169235|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81988||4|3|45
500853690|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-07|2011-07-22|Followup|2011-05-07|2011-06-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Moved|50.5||1|1|1|1|F|Multi-Race (None of the above)||18|No|Mother|28214|One Parent: Female|$15,000 to $19,999|Y|No||BBBS Board/Staff|General Community||Match Support|F|White||38|28226||Living w/ Significant Other|Child/Day Care Worker||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|500853959|7|0|2|500846213|1|0|2|500173015|2||-2||4|2|||-2||-2|0|13|||46|2|||1|81990||4|1|45
500859789|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-29|2013-02-28|Followup|2011-03-29|2011-03-30|Complete|Done|4|1|1|1|1|4|2|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|71.1||1|1|1|1|F|Black||18|Yes|Mother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||65|28078|||Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500860058|31|0|2|500856753|31|0|2|500169338|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|81992||4|3|45
500863413|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-31|2011-06-17|Followup|2010-08-31|2010-09-02|Complete|Done|2|2|2|2|2|2|2|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Time constraint|33.5||2|2|1|1|M|White||18|No|Mother|28227|One Parent: Female|$25,000 to $29,999||No||School|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Finance: Economist||0|6|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500001281|500863682|1|0|1|501292217|1|0|1|500281316|2||-2||4|1|||-2||-2|0|4|||7447|3|||1|81993||4|3|45
500867579|BBBS of Greater Charlotte|Main Office|C|Completed|2007-09-22|2013-04-02|Followup|2010-09-22|2010-11-10|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|66.3||1|1|1|1|M|Black||23|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|No||Faith Organization|General Community|Amachi|Match Support|M|Black||42|28269||Single|Finance: Banking||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|500867843|31|0|1|500577903|31|0|1|500195387|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|81994||4|1|45
500867581|BBBS of Greater Charlotte|Main Office|C|Completed|2007-09-28|2014-02-06|Followup|2010-09-28|2010-11-12|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|76.3||1|1|2|2|M|Black||21|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999||No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||40|28269|Masters Degree|Single|Finance: Accountant|28255|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|500867843|31|0|1|500708515|1|0|1|500195388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|81995||4|1|45
500870686|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-26|2011-06-17|Followup|2011-02-26|2011-05-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|39.7||1|1|1|1|M|Black||16|No|Mother|28078|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|M|White||38|28031|Bachelors Degree|Single|Business: Mgt, Admin||0|7|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008062|500870955|31|0|1|501101027|1|0|1|500248098|2||||4|3|||-2||-2|0|10|||46|2|||1|81996||4|0|45
500870948|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-22|2011-03-31|Followup|2010-05-22|2010-08-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|22.3||3|3|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||38|28204|Bachelors Degree|Single|Consultant|28036|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500003657|501616314|31|0|2|501559777|1|0|2|500358785|2||500003586||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|81997||4|0|45
500870996|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-16|2011-09-21|Followup|2011-05-16|2011-06-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|52.2||1|1|1|1|M|Black||23|No|Mother|28208|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community||Match Support|M|White||41|28209|Bachelors Degree|Divorced|Business: Sales|28202|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500871265|31|0|1|500869085|1|0|1|500176243|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81998||4|1|45
500871269|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-23|2011-02-09|Followup|2010-05-23|2010-08-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|44.6||1|1|1|1|F|Black||17|No|Mother|28205|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|F|Black||35|28227|Bachelors Degree|Single|Education: Teacher|28227|1|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500418342|31|0|2|500798511|31|0|2|500177506|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|81999||4|0|45
500871683|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-01|2016-02-22|Followup|2010-10-01|2010-11-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|100.7||1|1|1|1|M|Black||19|Yes|Aunt|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|M|White||46|28209|Masters Degree|Single|Self-Employed, Entrepreneur|28209|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500871952|31|0|1|500933829|1|0|1|500199601|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|82000||4|1|45
500872449|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-30|2013-02-28|Followup|2010-05-30|2010-06-16|Comprehension|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|69||1|1|2|2|M|Black||22|No|Mother|28211|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|White||37|28209|Masters Degree|Single|Business: Marketing|28208|1|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500872718|31|0|1|500846955|1|0|1|500178294|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|82001||4|2|45
500876141|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-27|2011-04-06|Followup|2010-07-27|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|44.3||1|1|1|1|M|Black||20|Yes|Mother|28216|One Parent: Female|$10,000 to $14,999|Y|No||Faith Organization|General Community|Amachi|Match Support|M|Black||62|28216||Married|Clergy||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|500876410|31|0|1|500899158|31|0|1|500183024|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|82003||4|1|45
500881634|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-14|NaT|Followup|2010-07-14|2010-07-23|Complete|Done|3|4|2|2|2|3|2.67|||||||||3|3|4|3|3|3|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|||104||1|2|1|2|M|Black||18||Mother|28213|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||38|28213||Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500881903|31|0|1|500816190|31|0|2|500277615|2||-2||2|1|||-2||-2|0|4|||46|2|||1|82005||4|3|45
500882189|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-22|2011-03-31|Followup|2010-05-22|2010-08-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Moved|22.3||2|2|1|1|F|Black||18|Yes|Mother|28216|One Parent: Female|$20,000 to $24,999||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Multi-race (Hispanic & White)||34|28211|Bachelors Degree|Single|Business: Human Resources|28280|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500003657|501616314|31|0|2|501535504|35|0|2|500360654|2||500003586||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|82007||4|0|45
500887773|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-25|2010-12-30|Followup|2010-05-25|2010-08-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|43.2||1|1|1|1|F|Black||17|Yes|Mother|28206|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Enrollment|F|Black||59|28205||Single|Business: Mgt, Admin|28277|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500888043|31|0|2|500847506|31|0|2|500177121|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|82008||4|0|45
500892903|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-29|2012-12-23|Followup|2010-05-29|2010-08-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Graduated|54.8||1|1|1|1|F|Black||22|Yes|Mother|28216|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||36|28273|Juris Doctorate (JD)|Single|Law: Lawyer|28052|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500893173|31|0|2|501189856|31|0|2|500268753|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|82009||4|0|45
500892907|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-29|2012-09-11|Followup|2010-05-29|2010-08-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Graduated|51.4||1|1|3|3|F|Black||22|No|Mother|28216|One Parent: Female|Unknown||No||Faith Organization|General Community|Amachi|Match Support|F|Hispanic||37|28203|Some College|Single|Education: Teacher|28217|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500893173|31|0|2|500188541|3|0|2|500268211|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|82010||4|0|45
500892914|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-16|2014-09-11|Followup|2011-02-16|2011-03-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Graduated|54.8||2|2|1|1|M|Black||20|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Sales|28269|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500893173|31|0|1|501964388|1|0|1|500429157|2||500003586||4|3|500000294|500000294|-2||-2|0|5|||7464|9|||1|82011||4|1|45
500896018|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-03|2014-08-14|Followup|2010-07-03|2010-09-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|73.4||1|1|1|1|F|Black||20|Yes|Mother|28027|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||40|28027|Bachelors Degree|Separated|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500896288|31|0|2|501225232|31|0|2|500269506|2||-2||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|82012||4|0|45
500896361|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-14|2014-02-27|Followup|2011-01-14|2011-03-31|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|61.4||2|2|1|1|F|Black||20|Yes|Mother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28075||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500012459|500896631|31|0|2|501276501|31|0|2|500291021|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|82014||4|0|45
500896588|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2016-06-15|Followup|2010-07-20|2010-07-22|Complete|Done|3|3|4|3|3|3|3.17|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|106.9||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28273|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||36|28269|Masters Degree|Married|Education|28205|6|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|500896858|3|15|2|500924445|1|0|2|500183434|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|82015||4|3|45
500897065|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-17|2012-05-23|Followup|2010-09-17|2010-12-02|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|32.2||3|4|2|3|F|Black||18|Yes|Mother|28269|Other/Unknown|Unknown||No||Service Organization|General Community||Match Support|F|Black||34|28105|Bachelors Degree|Married|Education: Admin|28202|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500897335|31|0|2|501454753|31|0|2|500384418|2||-2||4|1|||-2||-2|0|11|||7464|9|||1|82016||4|0|45
500897083|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-13|2012-11-19|Followup|2010-11-13|2011-01-17|Declined|Late||||||||4|1|4|1|3|4|2.83|||||||||3|3|3|4|4|4|3.5||||||4|4|4|4|||||||3|3|4|3|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Red|Amachi|Child/Family: Infraction of match rules/agency policies|36.2||1|1|1|1|M|Black||21|Yes|Mother|28269|One Parent: Female|Unknown|Y|No||Service Organization|General Community|Amachi|Match Support|M|White||54|28210||Married|Self-Employed, Entrepreneur||0|0|Holy Comforter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|500897335|31|0|1|501862348|1|0|1|500407273|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|11|||9216|7|||1|82017|268|4|1|45
500897406|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-26|2010-10-26|Followup|2010-06-26|2010-09-10|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Moved|40||1|1|1|1|F|Black||20|Yes|Mother|28270|Two Parent|$20,000 to $24,999|Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||37|28262|Masters Degree||Human Services: Social Worker||2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|501224558|31|0|2|500843337|31|0|2|500181575|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|9|||7464|9|||1|82018||4|0|45
500903951|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-04|2013-02-26|Followup|2011-04-04|2011-05-24|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Lost interest|58.8||1|1|1|1|M|Black||21|Yes|Mother|28203|One Parent: Female|Less than $10,000|Y|No||Faith Organization|General Community|Amachi|Match Support|M|White||34|28202|Bachelors Degree|Single|Finance: Banking||3|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|500904221|31|0|1|501167853|1|0|1|500252953|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|82022||4|1|45
500905603|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2010-10-20|Followup|2010-07-20|2010-10-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|39||2|3|2|2|F|Hispanic|Puerto Rican|20|No|Mother|28025|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||35|28081|Some College|Single|Law: Police Officer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|500905873|3|11|2|500783324|1|0|2|500185515|2||-2||4|1|||-2|500000294|-2|0|10|||2238|7|||1|82023||4|0|45
500905608|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-31|2010-10-20|Followup|2010-05-31|2010-06-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|40.7||1|1|1|1|M|Hispanic|Puerto Rican|22|No|Mother|28025|Two Parent|Unknown||No||Self|General Community||Match Support|M|White||42|28036|Associate Degree|Divorced|Business: Clerical|28078|9|5|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500002335|500905873|3|11|1|500772804|1|0|1|500178425|2||-2||4|1|||-2||-2|0|10|||7459|10|||1|82025||4|1|45
500910037|BBBS of Greater Charlotte|Main Office|C|Active|2009-06-22|NaT|Followup|2010-06-22|2010-08-02|Complete|Done|3|3|1|1|2|3|2.17|||||||||2|4|3|3|3|4|3.17|||||||||4|4|4|4||||||5|2|5|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||2|2|2|2||||||4|1|2.5|||||2|2|||||||||Green|||92.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||46|28277||Married|Business: Mgt, Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|500910307|31|0|1|500856100|1|0|1|500368834|2||-2||2|1|||-2||-2|0|10|||46|2|||1|82026||4|3|45
500910040|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2014-05-08|Followup|2010-05-29|2010-08-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|59.3||1|1|1|1|M|White||21|No|Mother|28270|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||31|28209|||Human Services: Non-Profit|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500910310|1|0|1|501600417|1|0|1|500363806|2||||4|3|||-2||-2|0|10|||7464|9|||1|82027||4|0|45
500914579|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-16|2014-12-04|Followup|2010-12-16|2010-12-27|Complete|Done|3|3|2|1|4|4|2.83|||||||||2|3|3|2|1|3|2.33|||||||||4|3|3|3.33||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|2|2|||||2|2|||||||||Yellow||Child: Severity of challenges|71.6||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|M|White||32|28277|Bachelors Degree|Single|Tech: Engineer|28117|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500914849|31|0|1|501345550|1|0|1|500323102|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|82030||4|3|45
500915359|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-10|2011-11-09|Followup|2010-11-10|2010-12-10|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Green||Volunteer: Time constraint|35.9||3|3|1|1|F|Black||19|No|Mother|28227|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|F|White||38|28105|PHD|Married|Human Services: Non-Profit|28110|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500915629|31|0|2|501189280|1|0|2|500311316|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|82031||4|3|45
500916976|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-08|2010-12-30|Followup|2010-09-08|2010-11-23|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|27.7||1|1|1|1|M|Black||21|Yes|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||35|28269|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500003657|500917246|31|0|1|501262371|31|0|1|500273621|2||500003586||4|1|500000294|500000294|-2||-2|0|8|||7496|10|||1|82032||4|0|45
500918264|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-13|2012-02-28|Followup|2011-02-13|2011-02-22|Blank|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Severity of challenges|48.5||1|1|1|1|M|Multi-Race (None of the above)||16|No|Mother|28227|Two Mothers|$45,000 to $49,999||No||Self|General Community||Match Support|M|Black||33|28269|Some College|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|500918534|7|0|1|501074231|31|0|1|500236477|2||-2||4|2|||-2||-2|0|10|||46|2|||1|82033||4|3|45
500930976|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-13|2013-04-26|Followup|2010-08-13|2010-10-28|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|56.4||1|1|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|Y|No||Service Organization|General Community||Match Support|F|Black||66|28205|Masters Degree|Single|Self-Employed, Entrepreneur||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500931243|31|0|2|501176751|31|0|2|500280106|2||-2||4|1|||-2||-2|0|11|||46|2|||1|82034||4|0|45
500931662|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-07|NaT|Followup|2010-09-07|2010-11-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||114.3||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$60,000 to $74,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||58|28270|Bachelors Degree|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500931932|31|0|1|500894084|1|0|1|500193824|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|82035||4|0|45
500934359|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-08|2010-12-21|Followup|2010-11-08|2010-12-01|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Time constraint|37.4||2|2|1|1|F|Black||20|Yes|Mother|28212|One Parent: Female|$10,000 to $14,999|Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||35|28215|Bachelors Degree|Single|Business: Human Resources||3|0|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|500934629|31|0|2|500991215|31|0|2|500209165|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|9|||7671|13|||1|82036||4|1|45
500934906|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-31|2013-02-12|Followup|2010-07-31|2010-08-04|Complete|Done|3||4|1|3|4||||||||||1|4|3|4|4|3|3.17|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|3|3.5|||||2|2|||||||||Red|Amachi|Volunteer: Lost contact with child/agency|66.5||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||52|28216|Bachelors Degree|Married|Tech: Engineer||13|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500935173|31|0|2|500859806|31|0|2|500186448|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|82037||4|3|45
500936718|BBBS of Greater Charlotte|Main Office|C|Completed|2007-12-20|2016-06-16|Followup|2010-12-20|2011-02-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Agency: Challenges with program/partnership|101.9||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28210|Bachelors Degree|Married|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500017732|500915629|31|0|1|501027885|1|0|1|500224574|2||-2||4|1|||-2|500014505, 500015184|-1|34|2|||46|2|||1|82038||4|1|45
500938154|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-12|NaT|Followup|2011-01-12|2011-03-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||98.1||2|2|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||32|28208|Associate Degree|Single|Service: Restaurant|28211|4|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500938424|31|0|1|501446421|1|0|1|500323753|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|82039||4|1|45
500948129|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-18|2016-06-30|Followup|2011-03-18|2011-05-19|Complete|Late|4|3|2|2|3|3|2.83|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Green|Amachi|Child: Graduated|75.4||2|2|1|1|F|Black||18|No|Mother|28217|One Parent: Female|$25,000 to $29,999|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||40|28203|Some College|Living w/ Significant Other|Finance: Banking|28281|1|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501891556|1|0|2|500438403|2||500003586||4|1|500000294|500000294|-2||-2|34|2|||7464|9|||1|82042||4|3|45
500948379|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-30|2011-04-21|Followup|2010-08-30|2010-10-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Lost interest|43.7||1|1|1|1|M|Black||23|No|Mother|28214|One Parent: Female|$30,000 to $34,999||Yes||Neighbor/Friend|General Community||Match Support|M|Black||48|28273||Married|Tech: Research/Design||0|0|General|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500011639|500948655|31|0|1|500952605|31|0|1|500192958|2||-2||4|2|||-2||-2|0|8|||6450|12|||1|82043||4|1|45
500948385|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-28|2013-01-09|Followup|2010-08-28|2010-10-04|Complete|Done|1|4|4|4|4|4|3.5|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|4|5|2|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Yellow||Child/Family: Lost contact with volunteer/agency|64.4||1|1|1|1|F|Black||17|No|Mother|28214|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Asian|Chinese|32|28216|||Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|500948655|31|0|2|500885771|4|16|2|500187434|2||-2||4|2|||-2||-2|34|2|||46|2|||1|82044||4|3|45
500954724|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-21|2011-06-17|Followup|2010-08-21|2010-11-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|45.9||1|1|1|1|F|Black||21|No|GrandMother|28273|One Parent: Female|Less than $10,000|Y|No||Service Organization|General Community||Match Support|F|Black||38|28273|||Finance: Accountant||0|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008062|500954994|31|0|2|500922418|31|0|2|500187226|2||-2||4|2|||-2||-2|0|11|||46|2|||1|82045||4|0|45
500956242|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-14|2013-02-28|Followup|2011-04-14|2011-06-18|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Moved|58.5||1|1|2|2|M|Multi-Race (None of the above)||19|No|Mother|28210|One Parent: Female|$20,000 to $24,999||Yes||Therapist/Counselor|General Community||Match Support|M|White||38|28210|||Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500956512|7|0|1|500189847|1|0|1|500259433|2||-2||4|3|||-2||-2|0|5|||7464|9|||1|82046||4|1|45
500958307|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-19|NaT|Followup|2010-09-19|2010-12-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi, Cabarrus County||113.9|Y|1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$40,000 to $44,999|Y|No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|Black||62|28213||Married|Finance: Economist||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500958577|31|0|1|500876132|31|0|1|500193868|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|82048||4|0|45
500961015|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-11|2014-10-02|Followup|2011-04-11|2011-06-26|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|77.7||1|1|1|1|M|Black||20|Yes|Mother|28227|Two Parent|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||43|28104||Married|Tech: Computer/Programmer|29607|10|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500013781|500934638|31|0|1|501210561|31|0|1|500257073|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||17161|11|||1|82049||4|0|45
500968246|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-29|2015-04-30|Followup|2011-04-29|2011-04-27|Complete|Done|4|3|4|1|4|1|2.83|||||||||1|3|3|2|2|4|2.5|||||||||3|3|3|3||||||3|2|3|3|2.75|||||||4|4|4|4|4|3|4|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child/Family: Lost contact with volunteer/agency|84||1|1|1|1|M|Black||19|No|Aunt|28269|One Parent: Female|$10,000 to $14,999|Y|No||Therapist/Counselor|General Community||Match Support|M|Black||35|28213|Bachelors Degree|Single|Business: Sales||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500968516|31|0|1|501179573|31|0|1|500251681|2||-2||4|1|||-2||-2|0|5|||46|2|||1|82051||4|3|45
500969481|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-22|2011-10-13|Followup|2010-07-22|2010-07-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Project Big|Child/Family: Lost contact with volunteer/agency|38.7||1|1|2|2|F|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|No||Therapist/Counselor|General Community||Match Support|F|Black||41|28209|Bachelors Degree|Single|Finance: Banking|28255|0|6|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500011639|500969749|31|0|2|501202092|31|0|2|500274109|2||-2||4|2|500004640||-2||-2|0|5|||130|1|||1|82052||4|1|45
500970181|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-31|2012-08-29|Followup|2010-10-31|2010-12-01|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Severity of challenges|58||1|1|1|1|M|Black|Other African|20|No|Mother|28208|One Parent: Female|$15,000 to $19,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||37|28210|Bachelors Degree|Single|Finance: Accountant||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|500970452|31|31|1|500969057|1|0|1|500203109|2||-2||4|3|||-2||-2|34|2|||46|2|||1|82053||4|1|45
500970495|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-10|2017-03-09|Followup|2010-09-10|2010-10-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|101.9||3|3|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$35,000 to $39,999||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black|Other African|44|28212||Single|Consultant||1|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500970766|31|0|2|500965698|31|31|2|500285645|2||-2||4|2|||-2||-2|7294|13|||46|2|||1|82054||4|1|45
500981435|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-24|2010-12-30|Followup|2010-07-24|2010-07-26|Complete|Done|4|4|4|4|3|4|3.83|||||||||2|4|4|3|1|4|3|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|2|1.5|||||2|2|||||||||Red||Volunteer: Time constraint|17.2||2|2|1|1|F|Multi-Race (None of the above)||21|No|Mother|28205|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||42|28203|||Business: Mgt, Admin|28210|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500981706|7|0|2|501623866|1|0|2|500374604|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|82055||4|3|45
500997812|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-12|2012-11-16|Followup|2011-01-12|2011-01-13|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|46.1||1|1|1|1|M|Black||20|No|Mother|28266|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community||Match Support|M|White||40|28203|Bachelors Degree|Single|Transport: Pilot||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|500998085|31|0|1|501429055|1|0|1|500329285|2||-2||4|1|||-2|500000294|-2|0|10|||7496|10|||1|82056||4|1|45
500997880|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-19|2016-07-29|Followup|2011-02-19|2011-04-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|101.3||1|1|1|1|M|Black||18|No|Mother|28204|Two Parent|$40,000 to $44,999||Yes||Self|General Community||Match Support|M|White||33|28202|Bachelors Degree|Married|Business: Marketing||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500998153|31|0|1|500990660|1|0|1|500237316|2||-2||4|1|||-2||-2|0|10|||46|2|||1|82057||4|1|45
501015201|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-13|2011-04-21|Followup|2010-11-13|2011-01-28|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|41.2||1|1|1|1|F|Black||19|No|Mother|28227|One Parent: Female|Less than $10,000||No|AARTF|Neighbor/Friend|General Community||Enrollment|F|White||36|28211|Bachelors Degree|Single|Finance: Auditor||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011639|501015474|31|0|2|500953684|1|0|2|500208541|2||-2||4|2|||-2||-2|6855|8|||46|2|||1|82059||4|0|45
501015962|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-12|2012-05-31|Followup|2011-02-12|2011-03-12|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|3|4|2|4|3.17|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||1|1|1|||||2|2|||||||||Yellow|Amachi|Volunteer: Time constraint|51.6||1|1|1|1|F|Black||18|Yes|GrandMother|28208|One Parent: Female|Less than $10,000||Yes||Self|General Community|Amachi|Enrollment|F|White||33|28202|Bachelors Degree|Single|Education: Teacher|28025|1|4|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|501065096|1|0|2|500241396|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||2238|7|||1|82060||4|3|45
501015965|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-29|2013-10-09|Followup|2011-04-29|2011-04-27|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|5|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2|||||||||Yellow|Amachi|Child: Lost interest|41.4||2|2|2|2|F|Black||17|Yes|Mother|28208|One Parent: Female|Less than $10,000||Yes||Self|General Community|Amachi|Match Support|F|Black||60|28269|Bachelors Degree|Married|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|500189376|31|0|2|500447721|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|82061||4|3|45
501023408|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-05|NaT|Followup|2010-11-05|2010-11-01|Complete|Done|3|1|4|2|3|3|2.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green|||100.3||1|1|1|1|M|Hispanic|Other South American|17|No|Mother|28273|One Parent: Female|Less than $10,000||Yes||Self|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501023677|3|15|1|501356600|1|0|1|500296545|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|82062||4|3|45
501045211|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-23|2011-09-12|Followup|2011-01-23|2011-04-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|43.6||1|1|1|1|M|Black||21|No|GrandMother|28269|Grandparents|$20,000 to $24,999||Yes||BBBS Board/Staff|General Community||Match Support|M|Black||47|28226|Bachelors Degree|Married|Business: Marketing||1|2|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500002335|501045484|31|0|1|501132288|31|0|1|500239114|2||-2||4|1|||-2||-2|0|13|||7671|13|||1|82066||4|0|45
501045214|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-30|2015-12-16|Followup|2010-11-30|2011-02-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|96.5||1|1|2|2|F|Black||20|No|Relative: Other|28269|Grandparents|$20,000 to $24,999||Yes||BBBS Board/Staff|General Community||Match Support|F|Black||35|28213|Masters Degree|Single|Business||4|0|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|277|60|598|500000170|500002335|501045484|31|0|2|500953330|31|0|2|500217682|2||-2||4|1|||-2|500014505, 500016394|-1|0|13|||46|2|||1|82067||4|0|45
501060196|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-26|2015-08-03|Followup|2010-11-26|2011-01-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|92.2||1|1|1|1|M|Black||19|No|Mother|28205|One Parent: Female|$15,000 to $19,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28226|Masters Degree|Single|Finance: Accountant||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501060469|31|0|1|501036081|1|0|1|500223215|2||-2||4|1|||-2||-2|34|2|||46|2|||1|82069||4|1|45
501068953|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-06|2012-03-31|Followup|2010-10-06|2010-11-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|29.8||2|2|2|2|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||40|28262|Bachelors Degree|Married|Law: Paralegal|28280|4|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008629|501060469|31|0|2|500874318|31|0|2|500380111|2||-2||4|1|||-2||-2|34|2|||46|2|||1|82074||4|1|45
501070152|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-29|2012-04-17|Followup|2010-11-29|2011-02-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|52.6||1|1|2|2|M|Black||20|Yes|Mother|28212|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community|Amachi|Match Support|M|Black||45|28079|Bachelors Degree|Married|Business||13|6|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501070425|31|0|1|501052547|31|0|1|500224306|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||7671|13|||1|82076||4|1|45
501072636|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-25|2013-06-19|Followup|2010-06-25|2010-07-02|Complete|Done|3|2|2|3|3|3|2.67|||||||||2|3|3|2|2|4|2.67|||||||||3|3|3|3||||||5|3|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2|||||||||Red||Child/Family: Lost contact with volunteer/agency|47.8||2|2|1|1|M|White||18||Mother|28134|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||50|28277|Bachelors Degree|Married|Tech: Management||10|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500004169|500965396|1|0|1|501637727|1|0|1|500368653|2||-2||4|3|||-2|500000294|-2|0|10|||7462|13|||1|82077||4|3|45
501074345|BBBS of Greater Charlotte|Main Office|C|Active|2008-03-31|NaT|Followup|2011-03-31|2011-06-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi, Cabarrus County||107.5||1|1|1|1|M|White||16|Yes|GrandMother|28025|Grandparents|Unknown||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|White||46|28027|Bachelors Degree|Divorced|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501074618|1|0|1|501158523|1|0|1|500250038|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|5635|9|||46|2|||1|82080||4|0|45
501078559|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-04|2012-06-21|Followup|2010-08-04|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|46.6||1|1|1|1|M|Black||22|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||37|28269|Bachelors Degree|Single|Medical: Admin|19380|0|9||Relative|Big|General Community||Match Support|277|60|598|500000170|500013781|501078832|31|0|1|501262050|1|0|1|500279449|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||0|11|||1|82082||4|1|45
501086649|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-20|2013-01-09|Followup|2010-11-20|2010-12-01|Complete|Done|4|3|3|3|4|4|3.5|4|3|4|2|3|4|3.33|5.11|3|3|3|3|3|3|3|4|4|4|4|3|3|3.67|-18.26|4|4|4|4|4|3|3|3.33|20.12|4|4|4|5|4.25|5|4|4|5|4.5|-5.56|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|3|4|3|3.33|20.12|2|2|2|4|4|4|-50|2|2|2|2|0||||||Red||Volunteer: Feels incompatible with child/family|37.7||1|1|1|1|M|Black||21|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Relative|General Community||Match Support|M|White||39|28205|Bachelors Degree|Single|Transport: Pilot|30320|2|0|Other Church Partner|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500004169|501086923|31|0|1|501833794|1|0|1|500399391|2||-2||4|3|||-2||-2|0|3|||7453|7|||1|82083|385|4|3|45
501092911|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-01|2015-08-18|Followup|2011-05-01|2011-05-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|87.6||1|1|1|1|M|Black||19||Mother|28226|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|M|White||37|28210|Some College|Single|Business: Mgt, Admin||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|501064244|31|0|1|501176101|1|0|1|500261235|2||-2||4|3|||-2||-2|0|4|||46|2|||1|82084||4|1|45
501098842|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-25|2012-03-31|Followup|2011-02-25|2011-02-16|Complete|Done|3|4|4|1|4|3|3.17|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||2|5|3|4|3.5|||||||4|4|4|4|3|3|3|3.57||||||||||3|4|3|3.33||||||2|1|1.5|||||2|2|||||||||Green||Child: Graduated|49.1||1|1|2|2|M|Black||23|No|Mother|28216|One Parent: Female|$25,000 to $29,999||No||Neighbor/Friend|General Community||Match Support|M|Black||60|28269|Bachelors Degree|Married|Business: Sales|28079|9|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008629|501099116|31|0|1|500967139|31|0|1|500247572|2||-2||4|1|||-2||-2|0|8|||4748|14|||1|82087||4|3|45
501099294|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-28|2011-06-17|Followup|2011-02-28|2011-05-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Unrealistic expectations|39.6||1|1|1|1|F|Black||22|No|Mother|28206|One Parent: Female|$15,000 to $19,999||Yes||Neighbor/Friend|General Community||Match Support|F|White||40|28205|Bachelors Degree|Single|Business: Sales|28277|0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008062|501099568|31|0|2|500897787|1|0|2|500244827|2||-2||4|2|||-2||-2|0|8|||46|2|||1|82089||4|0|45
501101149|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-01|NaT|Followup|2010-07-01|2010-09-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|||104.5||1|2|1|2|F|White||16||Mother|28270|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||55|28277|Masters Degree|Widowed|Consultant||5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|501101423|1|0|2|500834694|1|0|2|500276073|2||-2||2|2|||-2||-2|0|4|||7671|13|||1|82091||4|0|45
501101153|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-30|2013-08-30|Followup|2010-09-30|2010-11-08|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Severity of challenges|59||1|2|2|3|M|Black||19||Mother|28205|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||62|28214|Bachelors Degree|Married|Human Services: Non-Profit|28214|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501101427|31|0|1|500789916|1|0|1|500293277|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|82092||4|1|45
501114434|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-23|2014-06-12|Followup|2010-12-23|2011-02-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|65.6||1|1|1|1|M|Black||20|No|Uncle|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||33|28207|Masters Degree|Single|Finance: Accountant|28244|0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501114708|31|0|1|501315131|1|0|1|500324423|2||-2||4|3|500000294|500000294|-2||-2|0|10|||130|1|11|3|1|82093||4|1|45
501114443|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-08|2013-07-25|Followup|2010-10-08|2010-11-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|57.5||1|1|2|2|M|Black||22|No|Uncle|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||34|28205|Juris Doctorate (JD)|Married|Law: Lawyer||0|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501114708|31|0|1|501180846|1|0|1|500290376|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||46|2|||1|82094||4|1|45
501130354|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-15|2012-11-29|Followup|2011-02-15|2011-03-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|57.5||1|1|1|1|M|Black||21|Yes|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||BBBS Board/Staff|General Community|Amachi|Match Support|M|White||43|28205|Bachelors Degree|Married|Finance: Banking||7|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501130628|31|0|1|501124346|1|0|1|500245525|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|13|||46|2|||1|82100||4|1|45
501160894|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-07|2011-08-24|Followup|2010-11-07|2010-11-09|Complete|Done|4|2|3|3|4|4|3.33|||||||||3|3|3|3|3|3|3|||||||||3|3|3|3||||||3|3|3|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Yellow||Child/Family: Moved|33.5||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|$10,000 to $14,999||Yes||Self|General Community||Match Support|M|White||33|28204||Single|Real Estate: Realtor|28204|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501161168|31|0|1|501442606|1|0|1|500309909|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|82110||4|3|45
501164779|BBBS of Greater Charlotte|Main Office|C|Completed|2008-03-27|2011-06-17|Followup|2011-03-27|2011-04-01|Complete|Done|3|3|3|3|3|3|3|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|2|2|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2|||||||||Green||Volunteer: Moved|38.7||1|1|1|1|M|White||20|No|Mother|28210|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|White||40|22314|Bachelors Degree|Single|Business: Sales||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|501165053|1|0|1|501159259|1|0|1|500251850|2||-2||4|1|||-2||-2|0|10|||46|2|||1|82112||4|3|45
501165117|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-03|2011-06-09|Followup|2010-07-03|2010-09-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|35.2||2|3|1|2|F|Black||16||Mother|28205|Other/Unknown|Unknown||Yes||Self|General Community||Enrollment|F|White||34|28031||Single|Business: Clerical||0|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008629|501165391|31|0|2|501159184|1|0|2|500276436|2||-2||4|1|||-2||-2|0|10|||131|1|||1|82113||4|0|45
501174643|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-06|2012-11-08|Followup|2011-05-06|2011-06-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|42.1||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|Black||34|28214||Married|Business: Sales|28210|0|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011349|501174917|31|0|1|501687908|31|0|1|500358149|2||-2||4|3|||-2||-2|0|10|||7446|3|||1|82114||4|1|45
501176569|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-08|2012-02-29|Followup|2011-01-08|2011-01-04|Complete|Done|4|3|3|4|4|4|3.67|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green||Child/Family: Moved|37.7||1|1|1|1|M|Multi-race (Black & White)||18||Mother|28031|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28078|Bachelors Degree|Living w/ Significant Other|Education: Admin|28035|2|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501176843|36|0|1|501457533|1|0|1|500327489|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|82118||4|3|45
501184645|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-22|2011-08-05|Followup|2011-02-22|2011-05-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|41.4||1|1|2|2|M|Multi-race (Black & White)||19|No|Mother|28081|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||37|28027|Bachelors Degree|Married|Business: Sales|27263|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|501184919|36|0|1|500781896|1|0|1|500245777|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82120||4|0|45
501185594|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-29|2016-06-15|Followup|2011-03-01|2011-02-16|Complete|Done|3|4|4|3|3|4|3.5|||||||||3|4|3|2|4|4|3.33|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||4|2|3|||||2|2|||||||||Green||Child: Graduated|99.5||1|1|1|1|M|Multi-race (Black & White)||19|No|Mother|28227|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Consultant|28226|0|8|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501153366|1|0|1|500248756|2||-2||4|1|||-2||-2|0|4|||7452|6|||1|82121||4|3|45
501188642|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-28|2011-07-29|Followup|2011-04-28|2011-06-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|27||1|1|1|1|M|Black||18|No|Mother|28105|One Parent: Female|$45,000 to $49,999||No||Neighbor/Friend|General Community||Match Support|M|White||56|28270|Bachelors Degree|Married|Real Estate: Realtor|28277|11|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|501188916|31|0|1|501507244|1|0|1|500359356|2||-2||4|3|||-2||-2|0|8|||7496|10|||1|82122||4|1|45
501190094|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-20|2011-04-21|Followup|2010-11-20|2010-12-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|29||1|1|1|1|F|Black||21||Aunt|28215|Two Mothers|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|F|Black||42|28215||Single|Business: Clerical||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500009007|501190365|31|0|2|500721829|31|0|2|500314463|2||-2||4|3|||-2||-2|34|2|||46|2|||1|82123||4|1|45
501194364|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-27|2011-10-12|Followup|2010-05-27|2010-06-15|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Moved|40.5||1|1|1|1|F|Multi-Race (None of the above)||18|No|Mother|28216|Two Parent|$15,000 to $19,999||Yes||Self|General Community||Enrollment|F|Black||48|28214|Masters Degree|Single|Medical: Doctor, Provider|28207|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501194638|7|0|2|501143598|31|0|2|500265628|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|82124||4|1|45
501194563|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-21|2012-04-26|Followup|2011-04-21|2011-05-25|Complete|Done|3|2|4|1|4|4|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Time constraint|36.2||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$40,000 to $44,999||Yes||Self|General Community||Match Support|M|White||37|28269|Masters Degree|Single|Tech: Management|28262|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501194837|31|0|1|501486345|1|0|1|500357443|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82125||4|3|45
501195410|BBBS of Greater Charlotte|Main Office|C|Active|2008-08-15|NaT|Followup|2010-08-15|2010-10-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||103||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Asian||35|28210|Bachelors Degree|Married|Business: Sales|28217|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501195684|31|0|1|501277677|4|0|1|500278978|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|82126||4|0|45
501197292|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-06|2012-03-31|Followup|2010-06-06|2010-08-21|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|45.8||1|1|1|1|M|White||18|No|Mother|28110|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||50|28112|High School Graduate|Married|Business: Marketing|28105|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501197566|1|0|1|501240286|1|0|1|500269444|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82127||4|0|45
501201068|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2012-08-29|Followup|2010-10-30|2010-10-29|Complete|Done|3|2|2|1|4|4|2.67|3|2|3|2|4|4|3|-11|2|3|3|2|2|3|2.5|2|4|4|2|2|4|3|-16.67|4|4|4|4|4|4|4|4|0|4|4|4|3|3.75|4|4|5|3|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|2|2.5|2|2|2|25|2|2|1|1|100||||||Green||Child/Family: Lost contact with volunteer/agency|34||1|1|1|1|M|Black||21|No|Mother|28215|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||60|28262|Masters Degree|Single|Tech: Engineer||5|0|AA Task Force|Service Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501201342|31|0|1|501771844|31|0|1|500396764|2||-2||4|1|||-2|500000294|-2|6854|8|||9226|6|||1|82129|5730|4|3|45
501201092|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-26|2012-04-30|Followup|2010-08-26|2010-10-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Moved|44.1||1|1|1|1|M|White||20|No|Mother|28105|One Parent: Female|Unknown||No||Relative|General Community||Match Support|M|White||35|28270|Bachelors Degree|Single|Tech: Engineer|48121|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501201366|1|0|1|501285276|1|0|1|500280817|2||-2||4|3|||-2||-2|0|3|||7464|9|||1|82130||4|1|45
501201377|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-31|2016-08-26|Followup|2011-01-31|2011-01-24|Complete|Done|3|3|4|4|4|4|3.67|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Red||Child: Graduated|90.8||1|1|1|1|F|Hispanic||18|No|Mother|28212|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community||Match Support|F|Hispanic||65|28269|Masters Degree|Single|Medical: Admin|28262|8|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500017777|501201651|3|0|2|501497622|3|0|2|500331903|2||-2||4|3|||-2||-2|7016|11|||7446|3|||1|82131||4|3|45
501212047|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-07|NaT|Followup|2011-05-07|2011-05-31|Complete|Done|3|4|4|2|4|4|3.5|||||||||3|4|4|2|4|3|3.33|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|2|2|||||2|2|||||||||Green|||106.3||1|1|1|1|F|White||18|No|Father|28207|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||33|28226||Single|Human Services: Non-Profit|28205|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501212321|1|0|2|501242250|1|0|2|500264889|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|82133||4|3|45
501212662|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-23|2013-04-22|Followup|2010-06-23|2010-09-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|58||1|1|1|1|M|Multi-Race (None of the above)||16|Yes|Mother|28211|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Multi-Race (None of the above)||34|28205|Bachelors Degree|Single|Business: Sales|28210|0|10|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501212937|7|0|1|501252394|7|0|1|500269647|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|82134||4|0|45
501224287|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-30|2014-01-23|Followup|2010-10-30|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|62.8||1|1|1|1|M|Black||19|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||43|28262|Bachelors Degree|Married|Customer Service|28211|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501224558|31|0|1|501343190|31|0|1|500298289|2||-2||4|3|500000294|500000294|-2|500000294|-2|5635|9|||2230|7|||1|82137||4|1|45
501224288|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-17|2011-12-21|Followup|2010-11-17|2011-01-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Moved|37.1|Y|1|1|2|2|M|Black||17|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Enrollment|M|Black||49|28213|Bachelors Degree|Married|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500003657|501224558|31|0|1|500856618|31|0|1|500311410|2||500003586||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|82138||4|1|45
501226826|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-07|2011-09-29|Followup|2010-11-07|2010-12-28|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Lost contact with child/agency|34.7||1|1|1|1|M|Black||19|Yes|Mother|28215|One Parent: Female|Unknown||Yes||Relative|General Community|Amachi|Match Support|M|White||33|28202|Masters Degree|Single|Finance: Economist||0|8|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008629|501227093|31|0|1|501293480|1|0|1|500310244|2||-2||4|3|500000294|500000294|-2||-2|0|3|||7447|3|||1|82140||4|1|45
501226882|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-21|2013-06-07|Followup|2011-04-21|2011-07-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|61.5||1|1|2|2|M|Black||18|Yes|GrandMother|28027|Grandparents|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||52|28027|Bachelors Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500002335|501227158|31|0|1|500914929|31|0|1|500259581|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||2238|7|||1|82141||4|0|45
501227649|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-12|2011-11-08|Followup|2011-02-12|2011-04-29|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|32.8||2|2|1|1|M|White||16|Yes|GrandMother|28083|Grandparents|Unknown|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||37|28083|Masters Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|501227925|1|0|1|501485340|1|0|1|500340341|2||500003586||4|1|500000294|500000294, 500016374|-2||-2|0|10|||7464|9|||1|82146||4|0|45
501228176|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-05|2013-08-13|Followup|2010-08-05|2010-08-11|Complete|Done|3|4|4|3|4|4|3.67|||||||||3|3|3|4|3|4|3.33|||||||||4|4|4|4||||||5|3|4|2|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red||Volunteer: Lost contact with child/agency|60.3||1|1|1|1|M|Black||20|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|28078|Masters Degree|Married|Finance: Auditor|28202|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|501228452|31|0|1|501279790|1|0|1|500279399|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|82147||4|3|45
501228477|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-11|2011-06-17|Followup|2010-09-11|2010-11-26|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|33.1||1|1|1|1|M|Black||19|No|Mother|28105|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|M|White||59|28227|Some College|Married|Insurance|28211|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008062|501228753|31|0|1|501317923|1|0|1|500286344|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|82148||4|0|45
501234601|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-24|2012-08-29|Followup|2010-06-24|2010-09-08|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|50.2||1|1|2|2|F|Black||23|No|Mother|28215|Grandparents|Unknown||No|TV|Media|General Community||Match Support|F|Black||48|28211|Bachelors Degree|Single|Consultant|28278|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500008629|501234877|31|0|2|501223094|31|0|2|500271822|2||-2||4|2|||-2|500014505, 500015184|-1|56|1|||7462|13|||1|82150||4|0|45
501234604|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-23|2012-09-06|Followup|2010-07-23|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Severity of challenges|49.5||1|1|1|1|F|Black||19|No|Mother|28215|Grandparents|Unknown||No||Self|General Community||Match Support|F|Black||38|28213|Masters Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008629|501234880|31|0|2|501165150|31|0|2|500278984|2||-2||4|2|||-2||-2|0|10|||46|2|||1|82151||4|1|45
501234606|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-16|NaT|Followup|2010-09-16|2010-11-01|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||101.9||1|1|1|1|F|Black||16|No|Mother|28216|Grandparents|Unknown||No|TV|Media|General Community||Match Support|F|Black||42|28212|Bachelors Degree|Single|Unknown|28202|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501234882|31|0|2|501233675|31|0|2|500287478|2||-2||2|1|||-2||-2|56|1|||7464|9|||1|82152||4|1|45
501240369|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-10-09|Followup|2010-07-10|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|75||1|1|1|1|M|Black||20|Yes|Mother|28214|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||43|28269|Masters Degree|Single|Business: Mgt, Admin|28202|3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501240645|31|0|1|501240602|1|0|1|500272039|2||500003586||4|1|500000294|500000294|-2||-2|0|3|||131|1|||1|82154||4|1|45
501249455|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-03|2012-08-30|Followup|2010-12-03|2011-01-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|44.9||1|1|1|1|M|Black||22|No|Mother|28269|One Parent: Female|Unknown||Yes|Brochure|Media|General Community||Match Support|M|Black||36|28262|Masters Degree|Single|Finance: Banking||6|6|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|501249731|31|0|1|501488627|31|0|1|500317964|2||-2||4|3|||-2||-2|51|1|||7464|9|||1|82156||4|1|45
501250109|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-11|2013-02-27|Followup|2010-09-11|2010-08-20|Complete|Early|4|1|4|2|4|4|3.17|3|1|3|1|3|3|2.33|36.05|2|4|4|4|2|4|3.33|3|3|3|3|4|3|3.17|5.05|4|4|4|4|3|3|3|3|33.33|4|4|4|4|4|3|3|3|3|3|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|3|4|3.5|3|3|3|16.67|2|2|2|2|0||||||Red||Volunteer: Lost contact with child/agency|41.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28227|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501250385|31|0|1|501790515|31|0|1|500381167|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|82157|13945|4|3|45
501253904|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-17|2011-10-26|Followup|2011-02-17|2011-05-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|32.2|Y|1|1|1|1|M|White||18|No|Mother|28083|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||38|28115|High School Graduate|Married|Self-Employed, Entrepreneur||6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|501254180|1|0|1|501227814|1|0|1|500336488|2||-2||4|1||500000294|-2||-2|0|10|||7464|9|||1|82159||4|0|45
501257717|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-20|2012-10-30|Followup|2010-06-20|2010-09-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|52.3||2|2|2|2|F|Black||17|No|GrandMother|28203|Grandparents|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|White||31|28204|Bachelors Degree|Single|Finance: Banking||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|501257994|31|0|2|500839705|1|0|2|500271936|2||-2||4|1|||-2||-2|0|10|||46|2|||1|82161||4|0|45
501288021|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-27|2016-02-01|Followup|2010-08-27|2010-11-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|89.2||1|1|1|1|F|Black||16|No|Mother|28211|Two Parent|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28027|PHD|Single|Education: College Professor|27411|1|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501288299|31|0|2|501249338|31|0|2|500281778|2||-2||4|1|||-2||-2|0|10|||46|2|||1|82163||4|0|45
501292079|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-11|2013-07-18|Followup|2010-12-11|2011-02-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Lost interest|55.2||1|1|1|1|F|Black||17|Yes|GrandMother|28214|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||31|28203|Bachelors Degree|Single|Consultant|28204|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501292357|31|0|2|501519897|1|0|2|500323243|2||500003586||4|1|500000294|500000294|-2||-2|7294|13|||7464|9|||1|82164||4|1|45
501296349|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-01|2014-02-27|Followup|2010-12-01|2011-02-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|62.9||1|1|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||42|28214|Bachelors Degree|Single|Business: Mgt, Admin|28205|3|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501296627|31|0|2|501471640|31|0|2|500318555|2||||4|2|||-2|500000294|-2|0|4|||7464|9|||1|82165||4|1|45
501299223|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-26|2010-10-26|Followup|2010-06-26|2010-07-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Unrealistic expectations|28||1|1|1|1|F|White||23|No|Father|28214|One Parent: Male|Unknown||No||Therapist/Counselor|General Community||Match Support|F|White||35|28207|Associate Degree|Single|Business: Mgt, Admin|28217|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500009007|501299501|1|0|2|501158791|1|0|2|500273953|2||-2||4|3|||-2||-2|0|5|||7464|9|||1|82166||4|1|45
501300013|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-14|2012-05-01|Followup|2010-08-14|2010-10-29|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Agency: Challenges with program/partnership|44.6||2|2|2|2|F|Black||17|Yes|GrandMother|28273|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||40|28277|Associate Degree|Single|Unknown||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500003657|500561354|31|0|2|500188952|31|0|2|500281427|2||-2||4|1|500000294|500000294|-2||-2|7294|13|||7464|9|||1|82167||4|0|45
501300101|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-14|2015-05-11|Followup|2010-08-14|2010-10-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|80.9||1|1|4|4|F|Black||19|Yes|GrandMother|28273|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501300379|31|0|2|500346193|31|0|2|500281421|2||500003586||4|2|500000294|500000294|-2||-2|7294|13|||46|2|||1|82168||4|1|45
501309092|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-24|2011-12-21|Followup|2010-10-24|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|37.9||1|1|1|1|M|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Black||35|28269|Masters Degree|Single|Tech: Computer/Programmer|28110|3|0|Other|Service Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|501309370|31|0|1|501322778|31|0|1|500300356|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7452|6|||1|82170||4|1|45
501309634|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-12|NaT|Followup|2010-09-12|2010-10-29|Complete|Late|3|2|3|3|3|3|2.83|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Amachi||102.1||1|1|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||46|27704|Associate Degree|Divorced|Medical: Admin||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501309912|31|0|2|501046221|31|0|2|500281317|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7462|13|||1|82171||4|3|45
501313839|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-11|2013-06-18|Followup|2010-11-11|2011-01-18|Declined|Late||||||||3|2|3|3|4|4|3.17|||||||||2|3|4|4|2|4|3.17||||||3|4|4|3.67|||||||4|5|5|5|4.75||||||||||4|4|4|3|2|2|1|2.86||||||3|4|3|3.33|||||3|3|3||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|43.2||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||36|28204|Bachelors Degree|Single|Consultant||4|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501314117|31|0|1|501788563|1|0|1|500396680|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|82173|590|4|1|45
501330620|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-29|2011-03-17|Followup|2010-09-29|2010-12-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|29.5||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||43|28078|Masters Degree|Married|Self-Employed, Entrepreneur||1|6|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011184|501330898|31|0|2|501236896|31|0|2|500290146|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82175||4|0|45
501330628|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-29|2011-03-31|Followup|2010-09-29|2010-11-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|30||1|1|2|2|F|Black||19|Yes|Mother|28208|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||33|28215|Bachelors Degree|Single|Tech: Support, Writing|28204|6|0|Other|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|277|60|598|500000170|500003657|501330906|31|0|2|501245666|31|0|2|500287591|2||500003586||4|1|500000294|500000294|-2|500014506|-2|34|2|||7671|13|||1|82176||4|1|45
501340097|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-23|2016-09-19|Followup|2011-03-23|2011-05-19|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|77.9||2|2|1|1|M|Multi-race (Black & Hispanic)||17|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Hispanic||28|28277|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340376|38|0|1|501934966|3|0|1|500440292|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|82177||4|1|45
501340102|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-03|2013-04-25|Followup|2010-10-03|2010-11-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Time constraints|54.7||1|1|1|1|M|Multi-race (Black & Hispanic)||18|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||50|28269|Masters Degree|Married|Customer Service|28269|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340381|38|0|1|501316292|1|0|1|500287888|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|82178||4|1|45
501340105|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2013-06-27|Followup|2010-12-12|2011-02-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Graduated|54.5||1|1|1|1|F|Multi-race (Black & Hispanic)||21|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||53|28269||Married|Medical: Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340376|38|0|2|501514453|1|0|2|500322778|2||-2||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|82179||4|1|45
501342393|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-22|2014-06-06|Followup|2010-10-22|2010-10-29|Complete|Done|3|2|2|2|2|3|2.33|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||||||||||||Green||Child: Lost interest|67.4||1|1|1|1|F|White||19|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Business: Sales||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501342672|1|0|2|501210017|1|0|2|500293459|2||-2||4|1|||-2||-2|0|10|||46|2|||1|82180||4|3|45
501347056|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2015-10-12|Followup|2010-12-12|2010-12-09|Complete|Done|4|1|4|1|4|4|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|5|2|1|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Yellow||Child: Graduated|82||1|1|1|1|M|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28226|Bachelors Degree|Married|Tech: Engineer|28202|2|8|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|501347335|31|0|1|501217000|1|0|1|500322327|2||-2||4|2|||-2||-2|34|2|||7446|3|||1|82182||4|3|45
501347097|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-30|2014-10-16|Followup|2010-07-30|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|74.5||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||35|28078|Bachelors Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501347376|31|0|2|501099568|1|0|2|500278256|2||-2||4|2|||-2||-2|0|10|||46|2|||1|82183||4|1|45
501353940|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2011-05-11|Followup|2010-05-29|2010-06-20|Complete|Done|4|2|1|1|4|4|2.67|||||||||2|3|3|2|3|3|2.67|||||||||3|3|3|3||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2|||||||||Yellow|Amachi|Volunteer: Time constraint|23.4||3|3|1|1|M|Black||16|No|Relative: Other|28205|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||35|28211||Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010355|501354219|31|0|1|501587399|1|0|1|500360226|2||500003586||4|2|500000294|500000294, 500005291|-2||-2|34|2|||7464|9|||1|82185||4|3|45
501356328|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-21|2012-09-06|Followup|2010-11-21|2011-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|45.5||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||33|28269|Masters Degree|Single|Finance: Banking|28255|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501356607|31|0|2|501371070|31|0|2|500315101|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|82186||4|1|45
501361902|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-23|NaT|Followup|2011-01-23|2011-04-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||97.7||1|1|1|1|M|White||17|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28227|Bachelors Degree|Divorced|Business: Sales|28273|9|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501249611|1|0|1|501307192|1|0|1|500328424|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|82187||4|0|45
501363890|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-21|2012-08-29|Followup|2010-11-21|2010-12-09|Complete|Done|3|1|3|3|4|3|2.83|||||||||4|3|4|4|4|4|3.83|||||||||3|3|3|3||||||2|3|4|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Yellow||Volunteer: Lost contact with child/agency|45.2||1|1|2|2|M|Black||21|No|Mother|28216|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||37|28213|Masters Degree|Single|Medical: Healthcare Worker||2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501356607|31|0|1|500189279|31|0|1|500315105|2||-2||4|2|||-2|500000294|-2|0|8|||7464|9|||1|82188||4|3|45
501376745|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-01|2016-01-11|Followup|2011-04-01|2011-03-15|Complete|Early|3|4|4|4|4|4|3.83|||||||||2|4|3|4|2|3|3|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2|||||||||Green||Volunteer: Time constraint|81.3||1|1|3|4|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28269|||Business: Marketing||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|501377024|31|0|2|500725077|31|0|2|500350905|2||-2||4|1|||-2||-2|6854|8|||46|2|||1|82190||4|3|45
501378357|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-13|NaT|Followup|2011-02-13|2011-03-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||97||1|1|2|2|M|Multi-race (Black & White)||18|No|Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Mgt, Admin|28215|10|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501378636|36|0|1|501174997|31|0|1|500339619|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|82191||4|1|45
501379296|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-15|2011-08-24|Followup|2010-10-15|2010-11-05|Complete|Done|4|4|1|1|4|4|3|||||||||2|3|3|2|3|3|2.67|||||||||4|4|4|4||||||3|3|3|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||2|2|||||||||Green||Child/Family: Moved|34.3||1|1|1|1|M|Black||17||Mother|28227|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||33|28211|Bachelors Degree|Single|Unemployed||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|501161168|31|0|1|501296492|1|0|1|500297204|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|82192||4|3|45
501386394|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2011-03-25|Followup|2010-09-30|2010-09-30|Complete|Done|3|2|3|1|3|3|2.5|2|3|2|3|4|3|2.83|-11.66|3|3|3|3|3|3|3|1|4|4|2|2|4|2.83|6.01|4|4|4|4|4|4|4|4|0|4|5|4|4|4.25|2|4|4|4|3.5|21.43|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|3|4|3|3.33|3|4|3|3.33|0|4|2|3|2|1|1.5|100|2|2|1|1|100||||||Yellow||Volunteer: Time constraint|17.8||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||RTBM|M|Black||45|28215||Married|Tech: Research/Design||0|0|Mayfield Memorial|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500001281|501386675|31|0|1|501818567|31|0|1|500388796|2||-2||4|2|||-2||-2|34|2|||9212|7|||1|82193|3316|4|3|45
501388847|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-25|2011-09-23|Followup|2011-01-25|2011-02-24|Complete|Done|3|4|4|1|4|3|3.17|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|5|3|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|31.9||1|1|1|1|M|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||31|28202|Bachelors Degree|Single|Medical: Healthcare Worker|28207|1|5|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500001281|501389128|31|0|1|501452657|1|0|1|500334726|2||-2||4|1|||-2||-2|0|10|||7446|3|||1|82194||4|3|45
501389722|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-06|2014-04-24|Followup|2011-02-06|2011-04-23|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|62.5||1|1|1|1|F|White||21|No|Mother|28027|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||56|28027||Divorced|Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500012459|501390003|1|0|2|500787778|1|0|2|500337267|2||-2||4|1|||-2||-2|0|10|||46|2|||1|82195||4|0|45
501394276|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-19|2011-11-11|Followup|2010-11-19|2010-12-01|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Health|35.7||1|1|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community||Enrollment|F|White||33|28202|Bachelors Degree|Single|Arts, Entertainment, Sports||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501394557|31|0|2|501358317|1|0|2|500311375|2||-2||4|2|||-2||-2|7016|11|||7464|9|||1|82198||4|1|45
501394968|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-21|2011-03-30|Followup|2010-11-21|2010-12-09|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|28.2||1|1|1|1|M|Black||19|No|Mother|28278|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||44|28277|Masters Degree|Single|Business: Mgt, Admin|28277|0|2|BFKS|Special Event|Big|General Community||Match Support|277|60|598|500000170|500010765|501395249|31|0|1|501322428|1|0|1|500310512|2||-2||4|1|||-2||-2|0|10|||7454|8|||1|82199||4|1|45
501402710|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-19|2015-06-17|Followup|2010-06-19|2010-07-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|71.9||1|1|1|1|M|Black||18|No|Mother|30058|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28215||Married|Consultant|28285|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501402995|31|0|1|501728845|1|0|1|500368860|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82201||4|1|45
501409296|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-06|2011-11-11|Followup|2011-05-06|2011-06-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|30.2||1|1|1|1|M|Black||20|No|Mother|28278|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||54|28278|High School Graduate|Married|Tech: Management||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500001281|501409581|31|0|1|501632500|31|0|1|500357952|2||-2||4|2|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|82202||4|1|45
501428294|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-25|2011-10-25|Followup|2010-11-25|2011-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|35||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|M|Black||40|28209|Associate Degree|Married|Unknown|28208|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008629|501428579|31|0|1|501517334|31|0|1|500317955|2||-2||4|1|||-2||-2|6854|8|||7671|13|||1|82204||4|1|45
501428903|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-21|2015-02-25|Followup|2011-01-21|2011-01-04|Complete|Early|3|3|4|1|4|4|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2|||||||||Green||Child/Family: Lost contact with volunteer/agency|73.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|White||53|15001|Masters Degree|Single|Consultant|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501429188|31|0|1|501441245|1|0|1|500331206|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82205||4|3|45
501431901|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-22|2011-07-08|Followup|2010-09-22|2010-12-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|21.5||1|1|1|1|M|Black||22|No|Mother|28083|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||48|28081||Single|Medical: Healthcare Worker||0|0|AA Task Force|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500002335|501432186|31|0|1|501780241|31|0|1|500384909|2||-2||4|1|||-2||-2|0|8|||9226|6|||1|82207||4|0|45
501434147|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2011-03-31|2011-03-18|Complete|Done|2|1|1|4|1|4|2.17|3|1|4|3|1|3|2.5|-13.2|1|4|4|4|4|4|3.5|2|4|4|4|4|4|3.67|-4.63|4|4|4|4|4|4|4|4|0|4|3|4|5|4|4|5|2|5|4|0|4|4|4|4|4|4|1|3.57|4|4|4|4|4|4|4|4|-10.75|4|4|4|4|4|4|4|4|0|4|2|3|4|4|4|-25|2|2|2|2|0||||||Green|||83.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||26|28215|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501434432|31|0|1|501926474|31|0|1|500441566|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|82208|29966|4|3|45
501457406|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-20|2013-07-16|Followup|2010-08-20|2010-08-20|Complete|Done|4|4|4|4|4|3|3.83|||||||||4|4|3|2|4|4|3.5|||||||||4|4|4|4||||||2|3|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|46.9||1|1|1|1|M|Black||21|No|Mother|28269|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28205|||Finance: Banking|28217|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|501457691|31|0|1|501720969|1|0|1|500375964|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|82212||4|3|45
501457664|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-17|2010-09-29|Followup|2010-06-17|2010-09-01|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|15.4||1|1|1|1|M|Black||22|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||36|28203||Single|Business: Marketing||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501457949|31|0|1|501728924|1|0|1|500368257|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|82213||4|0|45
501506214|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-28|2016-06-23|Followup|2011-03-28|2011-03-18|Complete|Done|3|3|3|3|4|4|3.33|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|86.9||1|1|1|1|M|Black||19|No|Mother|28105|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||55|28173|||Unknown|28203|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501506506|31|0|1|501588885|31|0|1|500351462|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|82221||4|3|45
501516900|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-28|2015-08-27|Followup|2011-01-28|2011-01-04|Complete|Early|3|2|2|2|2|2|2.17|||||||||3|4|4|4|4|4|3.83|||||||||4|3|4|3.67||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|4|3.5|||||2|2|||||||||Green||Child: Graduated|78.9||1|1|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||39|28212|Bachelors Degree|Single|Medical: Healthcare Worker|28210|1|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500018987|501517192|31|0|2|501438601|31|0|2|500332399|2||-2||4|1|||-2||-2|6854|8|||7462|13|||1|82224||4|3|45
501522348|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-17|2013-02-28|Followup|2011-03-17|2011-03-14|Complete|Done|3|4|4|1|4|4|3.33|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||1|4|2.5|||||1|1|||||||||Red||Volunteer: Lost contact with child/agency|47.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28031|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Single|Retail: Sales|28117|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|501522640|36|0|1|501223351|1|0|1|500349995|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|82225||4|3|45
501525308|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-16|2015-06-18|Followup|2011-02-16|2011-03-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|76||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28205|Some College|Married|Retail: Sales|28206|1|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|501525600|31|0|1|501536144|1|0|1|500335230|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|82226||4|1|45
501526673|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-25|2013-10-09|Followup|2011-02-25|2011-05-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Lost interest|55.4||1|1|1|1|F|White||18|Yes||28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||34|28213|Bachelors Degree|Single|Real Estate: Realtor|28215|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500012459|501526965|1|0|2|501361484|1|0|2|500332705|2||500003586||4|2|500000294||-2||-2|0|10|||7496|10|||1|82227||4|0|45
501529921|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-06|2011-07-28|Followup|2011-02-06|2011-02-11|Complete|Done|3|4|1|4|4|4|3.33|||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|29.6||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||39|28209|Masters Degree|Married|Finance: Banking|28202|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501530213|31|0|2|501571404|1|0|2|500337752|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|82229||4|3|45
501535013|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-26|2011-07-22|Followup|2011-03-26|2011-03-18|Complete|Done|3|2|4|3|4|4|3.33|||||||||3|4|4|4|3|4|3.67|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Moved|27.9||1|1|1|1|M|Black||21|No|Mother|28273|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||36|28277|Bachelors Degree|Single|Retail: Mgt|28105|3|3|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501535305|31|0|1|501609664|31|0|1|500351430|2||-2||4|2|||-2|500000294|-2|0|10|||7496|10|||1|82231||4|3|45
501535016|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-12|2011-09-21|Followup|2011-01-12|2010-12-29|Complete|Done|3|4|4|3|4|4|3.67|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||5|3|4|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|4|4||||||4|3|3.5|||||2|2|||||||||Yellow||Volunteer: Time constraint|32.3||1|1|1|1|F|Black||18|No|Mother|28273|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||36|28277|Masters Degree|Single|Finance: Banking||0|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501535308|31|0|2|501438980|31|0|2|500331054|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|82232||4|3|45
501543766|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2010-10-26|Followup|2010-09-29|2010-10-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Moved|12.9||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28078|Masters Degree|Single|Business: Mgt, Admin|28115|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500009007|501544058|31|0|1|501422869|1|0|1|500383624|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|82233||4|1|45
501560189|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-11|2012-05-25|Followup|2011-03-11|2011-03-18|Complete|Done|3|2|3|2|3|3|2.67|||||||||3|4|4|4|3|3|3.5|||||||||4|4|4|4||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|26.5||2|2|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||39|28273||Single|Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501560485|31|0|2|501621478|31|0|2|500439156|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82235||4|3|45
501574315|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-11|2011-08-16|Followup|2011-02-11|2011-03-31|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|30.1||1|1|1|1|M|Black||15|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Relative|General Community|Amachi|Enrollment|M|White||33|28269|Bachelors Degree|Single|Finance: Banking|28202|4|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|501574611|31|0|1|501567524|1|0|1|500338128|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|3|||7464|9|||1|82239||4|1|45
501575246|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-20|2011-08-24|Followup|2011-02-20|2011-03-11|Complete|Done|4|2|4|2|4|4|3.33|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|3|4|4|3.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||2|4|3|||||2|2|||||||||Yellow||Volunteer: Time constraint|30.1||1|1|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||41|28212|Bachelors Degree|Married|Education: Teacher|28202|1|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500001281|501575542|31|0|1|501546450|31|0|1|500341366|2||-2||4|2|||-2||-2|0|10|||7671|13|||1|82240||4|3|45
501582592|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-20|2010-08-26|Followup|2010-08-20|2010-07-22|Declined|Early||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|12.2||1|1|1|1|M|Multi-Race (None of the above)||17|No|Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Hispanic||34|28227|||Insurance||2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500009007|501582912|7|0|1|501783333|3|0|1|500373122|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|82243||4|1|45
501588819|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-29|2011-06-09|Followup|2010-07-29|2010-07-26|Complete|Done|4|1|4|4|4|4|3.5|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1|||||||||Green||Volunteer: Time constraint|22.3||2|2|1|1|F|Black||18||Mother|28208|Two Parent|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28273|Masters Degree|Single|Govt: Mgmt/Admin|28216|1|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500008629|501589139|31|0|2|501454413|31|0|2|500373948|2||-2||4|1||500004640, 500005291|-2||-2|0|10|||129|1|||1|82244||4|3|45
501588821|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-10|2012-05-23|Followup|2011-02-10|2011-04-01|Declined|Late||||||||4|1|2|1|3|3|2.33|||||||||1|4|3|1|1|4|2.33||||||4|4|4|4|||||||5|1|1|2|2.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|4|3||||2|2|||||||Green||Volunteer: Lost contact with child/agency|27.4||1|1|2|2|F|Black||16||Mother|28208|Two Mothers|Unknown||Yes||Self|General Community||Match Support|F|Black||34|28273|Masters Degree|Living w/ Significant Other|Consultant|28273|1|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501589141|31|0|2|501359582|31|0|2|500429105|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|82245|28524|4|1|45
501597228|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-04|NaT|Followup|2010-09-04|2010-10-05|Complete|Done|3|4|4|4|3|2|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|Amachi||90.3||1|1|1|1|F|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||40|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28204|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501597548|31|0|2|501397328|31|0|2|500379964|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|82246||4|3|45
501604440|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-23|2014-11-19|Followup|2010-07-23|2010-06-10|Complete|Early|3|4|4|4|3|3|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|1|2.5|||||2|2|||||||||Green||Child: Graduated|63.9||1|1|1|1|M|Black||20|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||38|28269||Married|Govt||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501758365|3|0|1|500373108|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|82247||4|3|45
501604443|BBBS of Greater Charlotte|Main Office|C|Active|2009-07-10|NaT|Followup|2010-07-10|2010-06-11|Complete|Early|3|3|3|3|2|3|2.83|||||||||2|3|3|2|3|3|2.67|||||||||3|3|3|3||||||3|3|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|2|1.5|||||2|2|||||||||Green|||92.2||1|1|1|1|M|Black||18|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||35|28209|Bachelors Degree|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501729878|1|0|1|500371104|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|82248||4|3|45
501609876|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-13|2016-04-29|Followup|2010-07-13|2010-07-06|Complete|Done|3|3|3|3|3|3|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|Project Big|Child: Graduated|81.5||1|2|1|2|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Black||38|28269|Masters Degree|Single|Medical: Nurse|28262|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501610196|31|0|2|501425392|31|0|2|500373716|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7464|9|||1|82250||4|3|45
501614040|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-11|2013-02-28|Followup|2010-11-11|2010-11-12|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|39.6||1|1|1|1|M|Hispanic||16|No|Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||29|28273|||Facilities/Maintenance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|501614360|3|0|1|501864748|1|0|1|500404360|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|82254||4|1|45
501614044|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-06|2011-07-22|Followup|2011-04-06|2011-04-08|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|3|5|4|||||||4|4|4|4|4|4|4|4||||||||||2|2|3|2.33||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Lost contact with child/agency|27.5||1|1|1|1|F|Hispanic||19|No|Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||41|28273|Bachelors Degree|Single|Tech: Research/Design|28217|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501614360|3|0|2|501315493|1|0|2|500349169|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|82255||4|3|45
501614157|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-29|2013-04-04|Followup|2010-07-29|2010-07-29|Complete|Done|1||||3|3||||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||4|3|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2|||||||||Green||Volunteer: Moved|44.2||1|1|1|1|F|Black||21|No|Mother|28202|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28273|||Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|501614477|31|0|2|501596246|31|0|2|500374258|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82256||4|3|45
501614902|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-02|2011-03-31|Followup|2010-07-02|2010-09-16|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child/Family: Moved|20.9||1|1|1|1|M|Black||18|Yes|Mother|28105|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Black||39|28205|Bachelors Degree|Single|Business: Engineer||2|5|AA Task Force|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500003657|501615222|31|0|1|501745988|31|0|1|500370268|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||9226|6|||1|82257||4|0|45
501619710|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-16|2011-06-09|Followup|2011-03-16|2011-05-31|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|26.8||1|1|1|1|M|Black||20|No|Mother|28208|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|M|Black||38|28211|Masters Degree|Single|Finance: Banking|28202|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501620030|31|0|1|501380737|31|0|1|500344198|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|82259||4|0|45
501621811|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-16|2017-03-09|Followup|2011-03-16|2011-03-16|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|3|3|3|3|3|2.83|||||||||3|3|3|3||||||2|1|2|5|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|1|2.5|||||2|2|||||||||Yellow|Project Big|Child/Family: Lost contact with volunteer/agency|95.8||1|1|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||36|28269||Married|Self-Employed, Entrepreneur|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501622131|31|0|2|501621016|31|0|2|500344465|2||-2||4|2|500004640||-2||-2|0|10|||7464|9|||1|82260||4|3|45
501622497|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-31|2012-01-27|Followup|2011-03-31|2011-03-18|Complete|Done|3|2|3|3|3|3|2.83|||||||||2|4|3|4|3|3|3.17|||||||||4|4|4|4||||||4|5|5|3|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child/Family: Unrealistic expectations|33.9||1|1|1|1|M|Black||21|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||43|28227||Married|Business: Engineer|28227|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|501622817|31|0|1|501446203|31|0|1|500350734|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|82261||4|3|45
501626199|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-26|2013-09-30|Followup|2011-03-26|2011-03-18|Complete|Done|3|2|2|2|2|2|2.17|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|54.2||1|1|1|1|F|Black||21|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||33|28203|Masters Degree|Single|Finance: Accountant|28211|1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|501622822|31|0|2|501293622|1|0|2|500351814|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|82262||4|3|45
501626218|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-24|2014-12-18|Followup|2011-03-24|2011-03-18|Complete|Done|4|4|4|1|4|4|3.5|||||||||3|4|3|3|2|4|3.17|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|68.8||1|1|1|1|F|Black||20|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||30|11215|Bachelors Degree|Single|Consultant|11215|0|5|other|College Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501622822|31|0|2|501587214|31|0|2|500350222|2||-2||4|1|||-2|500000294|-2|0|10|||7670|5|||1|82263||4|3|45
501628854|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-15|2010-12-01|Followup|2010-06-15|2010-07-29|Complete|Done|4|2|3|2|2|3|2.67|||||||||3|3|3|3|3|3|3|||||||||3|3|3|3||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3||3|||||||3|3|3|||||1|1|||||||||Green|Amachi|Volunteer: Time constraint|17.5||3|3|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||34|28217|||Business: Engineer|28134|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010355|501629177|31|0|2|501595632|31|0|2|500368527|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|82264||4|3|45
501631059|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-26|2012-09-10|Followup|2010-05-26|2010-08-10|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|39.5||1|1|1|1|F|Black||18|No|Mother|28202|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||29|28216|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501631382|31|0|2|501589359|31|0|2|500364875|2||-2||4|2|||-2|500000294|-2|34|2|||7464|9|||1|82266||4|0|45
501631140|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-17|2016-03-03|Followup|2010-06-17|2010-07-02|Complete|Done|3|2|2|2|2|2|2.17|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|80.5||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Service: Hotel|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501631463|31|0|1|501628976|1|0|1|500367187|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82267||4|3|45
501631547|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2010-12-21|Followup|2010-09-30|2010-10-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Project Big|Volunteer: Lost contact with child/agency|14.7||2|2|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||32|28202|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501631870|31|0|1|501645587|1|0|1|500388261|2||500004641||4|2|500004640|500004640, 500005291|-2||-2|0|10|||7464|9|||1|82268||4|1|45
501639256|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-04|2011-12-21|Followup|2011-05-04|2011-06-30|Complete|Late|2|2|2|2|3|2|2.17|||||||||2|2|2|2|3|2|2.17|||||||||3|3|3|3||||||3|4|3|3|3.25|||||||4|4|4|3|3|3|3|3.43||||||||||3|4|3|3.33||||||3|2|2.5|||||2|2|||||||||Green|Amachi|Volunteer: Time constraint|31.6||2|2|1|1|M|Multi-Race (None of the above)||18|No|Mother|28211|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Black||35|28212||Single|Human Services: Non-Profit||2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|501639579|7|0|1|501721160|31|0|1|500360117|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|82269||4|3|45
501641337|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-07|2015-03-13|Followup|2010-08-07|2010-09-21|Complete|Done|3|4|4|3|4|4|3.67|||||||||3|3|3|4|3|4|3.33|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Moved|67.2||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||31|28269|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|2|500835981|31|0|2|500373972|2||-2||4|1||500000294|-2|500000294|-2|0|10|||46|2|||1|82270||4|3|45
501645192|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-21|2016-08-19|Followup|2010-07-21|2010-10-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|85||1|1|2|2|M|Hispanic||19|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501645515|3|0|1|501519306|1|0|1|500374818|2||-2||4|3||500016374|-2|500016374|-2|0|10|||7464|9|||1|82271||4|0|45
501669649|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-26|2012-03-31|Followup|2010-10-26|2010-10-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|29.1||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Enrollment|M|Black||67|28262||Married|Business: Mgt, Admin||32|0|Mayfield Memorial|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013709|501669987|31|0|1|501818546|31|0|1|500388262|2||-2||4|3|||-2||-2|6854|8|||9212|7|||1|82272||4|1|45
501670169|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2012-04-04|Followup|2010-09-30|2010-10-14|Declined|Done||||||||4|4|4|4|4|4|4|||||||||2||4|||4|||||||4|4|3|3.67|||||||4|2|4|5|3.75||||||||||4|4|4|4|4|4|4|4||||||4|3|4|3.67|||||4|2|3||||1|1|||||||Green||Volunteer: Time constraint|30.1||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|F|Black||32|28269||Single|Consultant|28209|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501670507|31|0|2|501466072|31|0|2|500379969|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|82273|2678|4|1|45
501686310|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2013-03-13|Followup|2010-10-30|2011-01-14|Expired|Late||||||||3|4|4|4|3|4|3.67|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||4|5|5|5|4.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|4|4||||1|1|||||||Red||Child/Family: Lost contact with volunteer/agency|40.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28211|One Parent: Female|Unknown||No|Radio|Media|General Community||Match Support|M|Black||34|28202|Juris Doctorate (JD)|Single|Law: Lawyer||1|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501686648|36|0|1|501818631|31|0|1|500392214|2||-2||4|3|||-2||-2|55|1|||7446|3|||1|82275|14832|4|0|45
501687515|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-21|2010-11-30|Followup|2010-05-21|2010-06-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|18.3||1|1|1|1|M|White||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||36|28078|Bachelors Degree|Single|Tech: Support, Writing|28204|2|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500001281|501687853|1|0|1|501284245|1|0|1|500361402|2||-2||4|1|||-2||-2|0|10|||6450|12|||1|82276||4|1|45
501714939|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-03|2012-12-23|Followup|2010-06-03|2010-06-29|Complete|Done|4|2|3|1|3|||||||||||2|3|3|2|3|4|2.83|||||||||3|3|3|3||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|42.7||1|1|1|1|M|Black||19|Yes|Mother|28105|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||34|28277||Single|Business: Sales|28206|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501715277|31|0|1|501584958|1|0|1|500365824|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|82279||4|3|45
501716763|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-07|2016-11-11|Followup|2011-05-07|2011-07-22|Expired|Late||||||||1|1|1|1|1|1|1|||||||||2|1|2|2|3|2|2||||||3|3|3|3|||||||2|3|2|2|2.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||1|1|||||||Red||Child/Family: Lost contact with volunteer/agency|78.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Amachi, Cabarrus County|Match Support|F|Black||39|28269||Single|Self-Employed, Entrepreneur|28027|7|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501716992|31|0|2|502112513|31|0|2|500449029|2||-2||4|3||500000294, 500016374|-2|500016374|-2|6854|8|||7458|9|||1|82280|30228|4|0|45
501721760|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-22|2016-11-01|Followup|2010-06-22|2010-09-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Infraction of match rules/agency policies|88.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||59|28269|Masters Degree|Married|Clergy||0|0|Coca Cola|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|501722098|31|0|1|501755476|1|0|1|500368545|2||-2||4|1|||-2|500000294|-2|0|10|||9610|3|||1|82281||4|0|45
501724170|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-06|2011-04-06|Followup|2010-07-06|2010-09-20|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Feels incompatible with child/family|21||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|Asian||41|28210|Bachelors Degree|Married|Tech: Management|28255|8|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008629|501724510|31|0|1|501681407|4|0|1|500370969|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|82282||4|0|45
501724491|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2011-03-30|Followup|2010-10-29|2010-12-06|Declined|Done||||||||4|2|4|1|1|4|2.67|||||||||1|1|3|1|1|2|1.5||||||4|4|4|4|||||||2|3|5|2|3||||||||||4|4|4|4|4|4|3|3.86||||||4|3|4|3.67|||||4|3|3.5||||1|1|||||||Green||Volunteer: Moved|17||1|1|1|1|M|Multi-race (Black & Asian)||19|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|M|White||42|28216||Divorced|Medical|28078|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501724831|39|0|1|501852487|1|0|1|500397005|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82283|7914|4|1|45
501725162|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2016-10-14|Followup|2010-10-29|2010-12-06|Blank|Done||||||||4|1|2|1|4|4|2.67|||||||||3|4|2|3|3|3|3||||||1|4|4|3|||||||5|1|5|5|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|2|3.33|||||4|3|3.5||||2|2|||||||Green||Agency: Challenges with program/partnership|83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501724831|39|0|1|501833178|1|0|1|500394157|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82284|16143|4|3|45
501725168|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-31|2013-12-18|Followup|2010-08-31|2010-08-18|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|51.6||2|2|1|1|F|Multi-Race (None of the above)||15|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28269|Bachelors Degree|Married|Human Services: Non-Profit||2|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017777|501724831|7|0|2|501824761|1|0|2|500381463|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|82285||4|3|45
501726201|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2015-01-30|Followup|2010-07-08|2010-08-06|Complete|Done|4|1|2|2|3|3|2.5|||||||||3|3|3|3|3|3|3|||||||||3|3|3|3||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|3|3|3.33||||||2|2|2|||||2|2|||||||||Red|Amachi|Child/Family: Moved|66.8||1|1|1|1|F|Black||17|Yes|Mother|28212|One Parent: Female|Unknown||Yes|YeaGod|Faith Organization|General Community|Amachi|Match Support|F|Black||51|28262|PHD|Married|Real Estate: Realtor||0|0|Weeping Willow|Faith Organization|Big|General Community||Enrollment|277|60|598|500000170|500008321|501726541|31|0|2|501734664|31|0|2|500371036|2||-2||4|3|500000294|500000294|-2||-2|5634|9|||9218|7|||1|82286||4|3|45
501731841|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-05|2013-08-30|Followup|2010-06-05|2010-08-20|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|50.8||1|1|1|1|F|Black||18|Yes|Father|28210|One Parent: Male|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||49|28277|Bachelors Degree|Single|Business: Mgt, Admin||4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|501732181|31|0|2|501182066|31|0|2|500367022|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||46|2|||1|82290||4|0|45
501735420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2015-08-13|Followup|2011-01-26|2011-01-04|Complete|Early|3|4|4|3|1|3|3|||||||||2|2|2|2|1|2|1.83|||||||||3|3|3|3||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2|||||||||Green||Child: Lost interest|66.5||2|2|2|2|F|Black||16||GrandMother|28215|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||41|28277|Bachelors Degree|Single|Business: Mgt, Admin||9|0|General|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500017732|501735760|31|0|2|500956022|1|0|2|500428818|2||-2||4|1|||-2||-2|6854|8|||6450|12|||1|82291||4|3|45
501744683|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-06|2012-11-28|Followup|2010-11-06|2011-01-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|36.7||1|1|1|1|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||56|28270|Some College|Separated|Unknown|28277|7|7|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500013781|501745023|31|0|1|501863268|31|0|1|500405317|2||-2||4|1|||-2||-2|0|10|||46|2|||1|82292||4|1|45
501750507|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-29|2011-02-09|Followup|2010-07-29|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|18.4||2|2|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||42|28262||Single|Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501750847|31|0|2|501582859|1|0|2|500374145|2||-2||4|1||500005291|-2||-2|0|10|||7464|9|||1|82293||4|1|45
501765404|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-20|2013-08-29|Followup|2011-04-20|2011-04-19|Complete|Done|4|2|3|2|4|4|3.17|3|3|3|1|4|3|2.83|12.01|3|3|3|4|2|3|3|2|3|3|2|3|3|2.67|12.36|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|5|5|4|4.25|-5.88|4|4|4|4|4|4|3|3.86|4|4|4|3|2|3|1|3|28.67|4|4|4|4|4|3|4|3.67|8.99|4|4|4|4|3|3.5|14.29|2|2|1|1|100||||||Yellow||Volunteer: Lost contact with child/agency|40.3||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Multi-race (Black & White)||28|28262||Single|Student: College|28262|3|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501765751|31|0|1|501958658|36|0|1|500443642|2||-2||4|2|||-2||-2|0|10|||9221|5|||1|82294|36416|4|3|45
501771253|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2011-04-21|Followup|2010-09-29|2010-12-14|Expired|Late||||||||4|1|4|1|4|4|3|||||||||2|4|4|3|3|4|3.33||||||4|4|4|4|||||||3|5|5|5|4.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|4|3||||||||||||Yellow||Volunteer: Feels incompatible with child/family|18.7||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||34|28269|Bachelors Degree|Single|Medical: Nurse|28054|3|6|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500009007|501741899|31|0|2|501322818|31|0|2|500383563|2||500003586||4|2|||-2|500000294|-2|0|10|||7462|13|||1|82296|13780|4|0|45
501776333|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-08|2013-07-25|Followup|2010-09-08|2010-09-02|Complete|Done|4|1|1|1|1|4|2|3|2|3|2|4|4|3|-33.33|4|4|4|2|2|4|3.33|3|3|3|2|3|3|2.83|17.67|4|4|4|4|3|3|3|3|33.33|4|4|4|3|3.75|4|4|4|4|4|-6.25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|2|2|0||||||Green||Volunteer: Moved|46.5||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28210|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|501776688|31|0|1|501832599|31|0|1|500381636|2||-2||4|1|||-2|500000294|-2|34|2|||7464|9|||1|82297|9814|4|3|45
501777213|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-15|2011-01-19|Followup|2010-12-15|2011-01-06|Declined|Done||||||||4|1|3|1|2|4|2.5|||||||||2|4|3|3|3|3|3||||||4|4|4|4|||||||5|1|2|4|3||||||||||4|4|4|4|4|4|4|4||||||4|4|2|3.33|||||2|2|2||||2|2|||||||Green||Volunteer: Moved|13.1||2|2|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||37|28217|Bachelors Degree|Single|Unemployed||0|0|Yahoo!|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500011639|501777568|31|0|1|501897253|31|0|1|500417596|2||-2||4|1||500005291|-2||-2|0|10|||32|2|||1|82298|21893|4|1|45
501788773|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-27|2012-06-28|Followup|2010-10-27|2010-12-14|Declined|Late||||||||3|2|2|1|4|4|2.67|||||||||2|4|3|4|4|3|3.33||||||4|4|3|3.67|||||||3|4|4|5|4||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||2|2|2||||2|2|||||||Green|Amachi|Volunteer: Moved|32||1|1|1|1|M|Black||18|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|RTBM|M|White||33|28202|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501789128|31|0|1|501845020|1|0|1|500393644|2||-2||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|82301|7735|4|1|45
501791428|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-29|2012-09-06|Followup|2010-07-29|2010-09-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|37.3||1|1|1|1|M|Black||19|No|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Multi-Race (None of the above)||33|28273|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501163776|31|0|1|501726049|7|0|1|500374912|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82304||4|1|45
501792675|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2011-09-21|Followup|2010-09-30|2010-09-14|Complete|Early|4|4|4|4|4|4|4|4|4|4|1|3|4|3.33|20.12|2|3|3|2|2|3|2.5|2|4|3|2|4|3|3|-16.67|4|4|4|4|4|4|4|4|0|4|3|3|3|3.25|3|3|2|3|2.75|18.18|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|4|3.5|4|3|3.5|0|2|2|2|2|0||||||Green||Volunteer: Moved|23.7||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|19085|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501793030|31|0|1|501664548|1|0|1|500386328|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|82305|12540|4|3|45
501796006|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-03|2011-12-20|Followup|2010-11-03|2010-12-09|Complete|Done|4|2|4|4|3|4|3.5|3|4|4|2|3|4|3.33|5.11|4|3|3|4|4|4|3.67|2|4|4|4|2|4|3.33|10.21|4|4|4|4|4|4|4|4|0|5|5|5|5|5||3|3|5|||4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|3|4|3.5|4|2|3|16.67|2|2|2|2|0||||||Green||Volunteer: Time constraint|25.5||3|3|1|1|F|Black||17|No|Mother|28031|Two Parent|Unknown|Y|Yes||School|General Community||Match Support|F|White||37|28078|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501489205|31|0|2|501621517|1|0|2|500396069|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|82306|6008|4|3|45
501811375|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-27|2013-08-28|Followup|2010-07-27|2010-10-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|49.1||1|1|3|3|F|Black||21|No|Mother|28027|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||41|28027|PHD|Single|Medical: Doctor, Provider|28075|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|501811730|31|0|2|501391123|31|0|2|500374230|2||-2||4|2|||-2|500016374|-2|0|8|||7464|9|||1|82307||4|0|45
501811385|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-27|2011-03-08|Followup|2010-07-27|2010-10-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|19.4||2|2|2|2|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||40|28075|Masters Degree|Married|Finance: Banking||8|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|501811730|31|0|2|500981458|31|0|2|500374643|2||-2||4|1||500016374|-2|500000294|-2|6854|8|||2238|7|||1|82308||4|0|45
501820715|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-23|2010-11-30|Followup|2010-10-23|2010-11-15|Declined|Done||||||||4|1|1|2|3|3|2.33|||||||||3|4|1|4|4|3|3.17||||||4|3|4|3.67|||||||4|3|3|1|2.75||||||||||4|4|4|4|2|4|4|3.71||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Green||Volunteer: Health|13.2||1|1|2|2|M|Black||22|No|Mother|28227|One Parent: Female|Unknown|Y|Yes||Relative|General Community||Match Support|M|Black||68|28212|Associate Degree|Married|Craftsman||25|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501821070|31|0|1|501049119|31|0|1|500387870|2||-2||4|1|||-2|500000294|-2|0|3|||2238|7|||1|82310|7575|4|1|45
501825910|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-24|2016-09-23|Followup|2010-08-24|2010-10-04|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Lost contact with child/agency|85||1|1|1|1|M|Black||16|Yes|Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|White||51|28214|Masters Degree|Married|Business: Sales|94108|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|501196986|1|0|1|500380446|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||7496|10|||1|82311||4|1|45
501829369|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-03|2012-01-10|Followup|2010-08-03|2010-10-18|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|29.2|Y|1|1|1|1|M|White||16|No|Mother|28027|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||61|28025||Married|Medical: Doctor, Provider||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|501829737|1|0|1|501687434|1|0|1|500376549|2||500003586||4|1|||-2||-2|0|10|||7464|9|||1|82312||4|0|45
501853848|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-30|2014-08-29|Followup|2010-11-30|2011-01-12|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Time constraint|56.9||1|1|1|1|M|Black||15|Yes|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|M|Black||33|28273|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501854219|31|0|1|501839466|31|0|1|500405366|2||-2||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|82316||4|1|45
501860404|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-21|2012-07-31|Followup|2011-01-21|2011-02-08|Declined|Done||||||||3|1|4|2|4|4|3|||||||||2|4|2||4|3|||||||4|4|4|4|||||||5|3|2|4|3.5||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||4|1|2.5||||2|2|||||||Green||Volunteer: Moved|30.3||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Enrollment|M|White||30|28202||Single|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501860777|31|31|1|501893096|1|0|1|500425993|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|82317|26821|4|1|45
501868921|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2010-12-21|Followup|2010-10-30|2010-10-29|Complete|Done|3|2|2|2|3|3|2.5|3|1|1|1|1|2|1.5|66.67|2|3|3|3|3|3|2.83|3|2|4|4|4|4|3.5|-19.14|3|3|3|3|4|3|3|3.33|-9.91|3|5|3|5|4|4|5|5|4|4.5|-11.11|4|4|4|4|3|4|3|3.71|4|4|4|4|3|3|3|3.57|3.92|3|3|3|3|2|4|3|3|0|3|3|3|2|1|1.5|100|2|2|1|1|100||||||Yellow||Volunteer: Lost contact with child/agency|13.7||2|2|1|1|F|Black||19|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||34|28217|Juris Doctorate (JD)|Married|Law: Lawyer|28204|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501869291|31|0|2|501220647|31|0|2|500398441|2||-2||4|2||500005291|-2||-2|0|10|||7464|9|||1|82319|4527|4|3|45
501877268|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2011-10-13|Followup|2011-01-26|2011-02-02|Comprehension|Done||||||||4|3|4|4|3|4|3.67|||||||||2|3|2|2|1|3|2.17||||||4|4|4|4|||||||4|5|3|4|4||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||4|4|4||||2|2|||||||Red||Child/Family: Lost contact with volunteer/agency|20.5||1|1|1|1|M|Black||19|No|Mother|28213|One Parent: Female|Unknown|Y|Yes|Radio|Media|General Community||Match Support|M|White||33|28269|||Construction||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011639|501877641|31|0|1|501942543|1|0|1|500429020|2||-2||4|3|||-2||-2|55|1|||7447|3|||1|82323|28469|4|2|45
501904094|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-15|2013-06-19|Followup|2011-01-15|2011-01-04|Complete|Done|4|2|3|2|4|4|3.17|4|1|4|2|4|4|3.17|0|4|3|3|4|4|4|3.67|2|4|4|3|4|4|3.5|4.86|4|4|4|4|4|4|4|4|0|5|4|4|4|4.25|3|4|2|5|3.5|21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0||||||Red||Volunteer: Lost contact with child/agency|41.1||1|1|1|1|F|Black||16|No|Mother|28214|One Parent: Female|Unknown|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||56|28208|Some College|Single|Finance: Accountant|28203|19|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500004169|501904482|31|0|2|501342148|31|0|2|500420809|2||-2||4|3|||-2|500000294|-2|34|2|||7446|3|||1|82324|23717|4|3|45
501919423|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-24|NaT|Followup|2011-03-24|2011-05-11|Declined|Late||||||||4|4|4|4|4|4|4|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||4|5|4|3|4||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|3|3.5||||1|1|||||||Green|Project Big||83.7||1|1|1|1|M|Multi-race (Black & Hispanic)||17|No|Mother|28214|One Parent: Female|Unknown||No|TV|Media|General Community|Project Big|Match Support|M|White||34|28164|Masters Degree||Finance|28210|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501919819|38|0|1|502034798|1|0|1|500442066|2||500004641||2|1|500004640|500004640|-2||-2|56|1|||7464|9|||1|82325|36152|4|1|45
501936316|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-28|2016-08-29|Followup|2011-01-28|2011-01-28|Declined|Done||||||||3|3|3|2|2|2|2.5|||||||||3|3||3|3|3|||||||3|3|3|3|||||||4|5|4|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Child/Family: Lost contact with volunteer/agency|79||1|1|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||54|28203|||Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|501936714|31|0|1|501872326|1|0|1|500428557|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|82326|28181|4|1|45
501938887|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2011-10-26|Followup|2011-04-30|2011-06-14|Declined|Done||||||||4|3|4|3|4|4|3.67|||||||||2|3|3|3|3|3|2.83||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||1|1|||||||Red||Child/Family: Lost contact with volunteer/agency|17.9||1|1|1|1|M|Black||18|No|Mother|28205|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|M|White||34|28205|||Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|501939285|31|0|1|502014005|1|0|1|500447313|2||-2||4|3|||-2||-2|0|8|||7496|10|||1|82328|38283|4|1|45
501955313|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-29|2011-08-16|Followup|2011-01-29|2011-02-01|Declined|Done||||||||4|2|3|2|4|4|3.17|||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||1|3|3|3|2.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Volunteer: Moved|18.5||2|2|1|1|F|Black||16||Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28270||Single|Business: Clerical||10|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500010765|501955711|31|0|2|500915390|1|0|2|500427542|2||-2||4|1||500005291|-2||-2|0|10|||130|1|||1|82331|27768|4|1|45
501957505|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-25|2012-03-31|Followup|2011-02-25|2011-04-18|Declined|Late||||||||4|1|1|1|3|4|2.33|||||||||2|3|4|3|3|3|3||||||4|3|4|3.67|||||||5|2|5|5|4.25||||||||||4|4|4|4|4|4|4|4||||||4|3|4|3.67|||||3|3|3||||1|1|||||||Green|Amachi|Volunteer: Moved|25.1||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||55|28078|||Business: Marketing|28070|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501957903|31|0|1|501718938|1|0|1|500432245|2||-2||4|1|500000294||-2||-2|0|10|||7464|9|||1|82333|30477|4|1|45
501990745|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-14|2012-08-29|Followup|2011-05-14|2011-05-18|Complete|Done|3|3|4|3|4|4|3.5|2|2|3|1|1|2|1.83|91.26|3|3|3|4|4|4|3.5|3|3|3|3|4|3|3.17|10.41|4|4|4|4|3|3|3|3|33.33|4|3|3|5|3.75|5|4|3|5|4.25|-11.76|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|3|4|3|3.33|20.12|4|3|3.5|4|4|4|-12.5|2|2|1|1|100||||||Red||Child: Severity of challenges|27.5||1|1|1|1|M|Black||16||Mother|28269|One Parent: Female|Unknown||Yes||BBBS Board/Staff|General Community||Match Support|M|Black||35|28213||Married|Human Services: Youth Worker||0|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500011746|501991144|31|0|1|502098002|31|0|1|500447817|2||-2||4|3|||-2||-2|0|13|||4748|14|||1|82336|38490|4|3|45
502076679|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2012-09-06|Followup|2011-04-30|2011-06-17|Declined|Late||||||||4|2|3|2|3|4|3|||||||||3|3||3|3|3|||||||3|3|3|3|||||||2|4|4|4|3.5||||||||||4|4|4|4||4|4|||||||4|4|4|4|||||3|3|3||||2|2|||||||Red||Volunteer: Time constraint|28.3||1|1|1|1|M|Black||17|No|Mother|28273|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||37|28278|||Finance: Banking||0|0|AA Task Force|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502077103|31|0|1|502003579|1|0|1|500446859|2||-2||4|3|||-2||-2|0|4|||9228|10|||1|82347|38100|4|1|45
502083450|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-20|2011-08-26|Followup|2011-05-20|2011-08-04|Expired|Late||||||||4|4|4|4|3|4|3.83|||||||||4|2|3|2|4|3|3||||||4|4|4|4|||||||3|4|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green|Amachi|Volunteer: Time constraint|15.2||2|2|1|1|M|Black||16|No|Mother|28027|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||44|28262||Divorced|Service: Restaurant|28027|0|10|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|502083874|31|0|1|502104415|31|0|1|500453680|2||500003586||4|1|500000294|500005291|-2||-2|7016|11|||7464|9|12|3|1|82348|39542|4|0|45
501868918|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-27|2014-05-22|Baseline|2010-05-24|2010-05-27|Complete|Done|3|3|3|4|3|3|3.17|||||||||3|4|4|2|3|3|3.17|||||||||4|4|3|3.67||||||3|3|5|5|4|||||||3|4|3|3|4|3|2|3.14||||||||||3|4|3|3.33||||||2|3|2.5|||||1|1|||||||||Green||Child: Graduated|47.8||1|1|1|1|M|Black||20|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||35|27612|Juris Doctorate (JD)|Living w/ Significant Other|Law|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|501869291|31|0|1|501921115|1|0|1|500454496|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|128915|-1|4|3|44
501365520|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-28|2011-07-29|Baseline|2010-05-24|2010-05-28|Complete|Done|3|3|4|3|3|3|3.17|||||||||3|4|3|3|3|3|3.17|||||||||4|3|3|3.33||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Green||Child/Family: Lost contact with volunteer/agency|14||1|1|4|4|F|Black||19||Mother|28203|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||38|28214|Bachelors Degree|Single|Business: Clerical|28273|2|3|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008629|501365799|31|0|2|500868727|31|0|2|500454745|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|129441|-1|4|3|44
502083504|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-26|2011-10-20|Baseline|2010-05-26|2010-05-26|Complete|Done|4|4|4|1|4|4|3.5|||||||||3|3|3|3|4|3|3.17|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red|Amachi|Volunteer: Lost contact with child/agency|16.8||1|1|2|2|M|Asian||18|Yes|Mother|28025|One Parent: Female|Unknown||Yes||Service Organization|General Community|Amachi|Match Support|M|Black||52|28027||Married|Business: Human Resources|28273|0|0|Big Champions|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|502083919|4|0|1|502089653|31|0|1|500454472|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|11|||7461|12|||1|131834|-1|4|3|44
502124485|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-28|2011-08-30|Baseline|2010-05-26|2010-05-28|Complete|Done|4|1|2|1|2|4|2.33|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green||Volunteer: Time constraint|15.1||2|2|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|White||32|28206||Single|Medical: Nurse||0|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500008629|502142970|31|0|2|502066586|1|0|2|500454581|2||-2||4|1|||-2||-2|0|4|||7438|1|||1|132622|-1|4|3|44
502180719|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-04|2014-03-20|Baseline|2010-05-28|2010-06-04|Complete|Done|4|2|4|4|4|4|3.67|||||||||2|4|4|4|4|4|3.67|||||||||3|4|4|3.67||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|45.5||2|2|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|Black||42|28273|Masters Degree|Divorced|Business: Marketing||1|6|Michael Baisden|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502181148|31|0|2|502184470|31|0|2|500454904|2||500004772||4|1|500000294, 500004640, 500004901|500000294|-2|500000294|-2|7016|11|||11146|1|||1|134611|-1|4|3|44
502045254|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-08|2015-10-09|Baseline|2010-05-28|2010-06-08|Complete|Done|2|4|4|4|3|4|3.5|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||2|4|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|3|2|3||||||3|3|3|||||1|1|||||||||Yellow||Child: Graduated|64||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502171015|31|0|2|500454926|2||-2||4|2|||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1|134736|-1|4|3|44
501224282|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-16|2012-06-14|Followup|2010-10-16|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Feels incompatible with child/family|43.9||2|2|1|1|F|Black||15|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||35|28215|Bachelors Degree|Single|Finance: Banking|28262|2|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501224558|31|0|2|501389463|31|0|2|500296679|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||7453|7|||1|134997||4|1|45
502034622|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-23|2010-07-22|Baseline|2010-06-01|2010-06-23|Complete|Done|3|1|4|1|3|4|2.67|||||||||3|4|4|2|4|4|3.5|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child/Family: Infraction of match rules/agency policies|1||1|1|2|2|M|Black||18|No|Mother|28214|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500009007|502035021|31|0|1|502127058|1|0|1|500456536|2||-2||4|1|||-2||-2|0|4|||130|1|||1|135405|-1|4|3|44
501965241|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-29|2012-07-31|Baseline|2010-06-02|2010-06-29|Complete|Done|4|1|4|1|1|1|2|||||||||1|1|4|4|4|4|3|||||||||4|4|4|4||||||4|3|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Green||Child/Family: Lost contact with volunteer/agency|25.1||1|1|1|1|M|Black||19||Mother|28208|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|M|Black||37|28210||Single|Law||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501578929|31|0|1|502081691|31|0|1|500457757|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|137801|-1|4|3|44
501994951|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2014-09-18|Baseline|2010-06-03|2010-06-15|Complete|Done|3|3|3|1|4|4|3|||||||||4|4|3|4|4|4|3.83|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|3|3|3|3|3.43||||||||||3|3|3|3||||||3|1|2|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|51.1||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|Unknown||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||36|28078||Single|Customer Service||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501843047|31|0|2|502048623|31|0|2|500455478|2||-2||4|2|||-2||-2|7294|13|||7464|9|||1|139614|-1|4|3|44
502053779|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2012-09-05|Baseline|2010-06-04|2010-06-15|Complete|Done|3|3|3|2|3|4|3|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||3|3|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Red||Child/Family: Feels incompatible with volunteer|26.7||2|2|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community||Match Support|F|Black||39|28216|||Education: College Professor||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|502054203|31|0|2|501912080|31|0|2|500455628|2||-2||4|3|||-2||-2|7295|11|||7464|9|||1|140517|-1|4|3|44
502142541|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-18|2015-07-23|Baseline|2010-06-07|2010-06-18|Complete|Done|3|4|4|3|4|4|3.67|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|5|3|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|61.1||1|1|2|2|F|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502142970|31|0|2|501905673|31|0|2|500455759|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|141478|-1|4|3|44
502045254|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-08|2015-10-09|Followup|2011-05-28|2011-05-18|Complete|Done|3|3|4|3|4|4|3.5|2|4|4|4|3|4|3.5|0|2|4|3|2|3|3|2.83|2|4|3|2|2|3|2.67|5.99|4|4|4|4|4|4|4|4|0|4|3|2|4|3.25|2|4|3|3|3|8.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|4|3|2|3|0|3|2|2.5|3|3|3|-16.67|2|2|1|1|100||||||Yellow||Child: Graduated|64||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502171015|31|0|2|500454926|2||-2||4|2|||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1|142235|134736|4|3|45
501987736|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-29|2014-06-18|Baseline|2010-06-08|2010-06-29|Complete|Done|4|4|4|2|4|4|3.67|||||||||2|4|4|2|4|4|3.33|||||||||4|2|2|2.67||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|1|1.5|||||1|1|||||||||Green||Child: Graduated|47.6||1|1|1|1|F|White||20|No|Father|28217|One Parent: Male|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||40|28203|Masters Degree|Single|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501988135|1|0|2|502109789|1|0|2|500456045|2||-2||4|1|||-2||-2|6855|8|||7464|9|||1|142908|-1|4|3|44
501604440|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-23|2014-11-19|Followup|2011-07-23|2011-07-12|Complete|Done|3|3|3|3|4|4|3.33|||||||||2|3|3|2|3|3|2.67|||||||||3|3|3|3||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Child: Graduated|63.9||1|1|1|1|M|Black||20|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||38|28269||Married|Govt||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501758365|3|0|1|500373108|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|144352||4|3|45
502072733|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2010-09-02|Baseline|2010-06-10|2010-06-15|Complete|Done|3|3|3|4|4|4|3.5|||||||||2|2|3|3|1|4|2.5|||||||||4|4|4|4||||||3|4|5|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|1|2|||||2|2|||||||||Green||Child: Lost interest|2.6||1|1|2|2|F|Black||19|No|GrandMother|28216|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|White||33|28078|High School Graduate|Single|Self-Employed, Entrepreneur|28269|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010765|502073157|31|0|2|502080569|1|0|2|500456384|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|144779|-1|4|3|44
501938310|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-25|2010-08-24|Baseline|2010-06-11|2010-06-25|Complete|Done|3|3|3|2|2|3|2.67|||||||||1|2|2|2|1|2|1.67|||||||||4|3|3|3.33||||||3|4|2|4|3.25|||||||2|3|3|3|2|2|2|2.43||||||||||2|2|2|2||||||3|3|3|||||1|1|||||||||Green||Child: Lost interest|2||1|1|4|5|F|White||20|Yes|Father|28081|Two Parent|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|277|60|598|500000170|500002335|501938708|1|0|2|501306527|1|0|2|500456460|2||500003586||4|1||500000294|-2|500014681, 500016374|-2|0|10|||7464|9|||1|145202|-1|4|3|44
501604443|BBBS of Greater Charlotte|Main Office|C|Active|2009-07-10|NaT|Followup|2011-07-10|2011-07-18|Complete|Done|1|4|4|4|3|3|3.17|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|||92.2||1|1|1|1|M|Black||18|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||35|28209|Bachelors Degree|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501729878|1|0|1|500371104|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|145261||4|3|45
501868918|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-27|2014-05-22|Followup|2011-05-27|2011-04-20|Complete|Early|3|4|3|3|4|4|3.5|3|3|3|4|3|3|3.17|10.41|2|3|3|2|2|3|2.5|3|4|4|2|3|3|3.17|-21.14|4|4|4|4|4|4|3|3.67|8.99|2|4|4|2|3|3|3|5|5|4|-25|4|4|4|4|4|4|3|3.86|3|4|3|3|4|3|2|3.14|22.93|3|3|3|3|3|4|3|3.33|-9.91|3|2|2.5|2|3|2.5|0|2|2|1|1|100||||||Green||Child: Graduated|47.8||1|1|1|1|M|Black||20|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||35|27612|Juris Doctorate (JD)|Living w/ Significant Other|Law|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|501869291|31|0|1|501921115|1|0|1|500454496|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|146415|128915|4|3|45
502106926|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-25|2012-06-28|Followup|2011-05-25|2011-04-20|Complete|Early|3|1|4|1|2|4|2.5|4|4|4|1|2|4|3.17|-21.14|1|4|4|4|1|4|3|1|2|4|3|3|3|2.67|12.36|4|4|4|4|4|4|4|4|0|5|4|3|3|3.75|5|1|5|1|3|25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|4|4|4|4|-8.25|2|2|2|4|4|4|-50|2|2|2|2|0||||||Red||Volunteer: Time constraint|25.1||2|2|1|1|M|Black||17|No|Mother|28031|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28031||Single|Govt||0|0|AA Task Force|Special Event|Big|General Community||Match Support|277|60|598|500000170|500011746|502107353|31|0|1|502072628|1|0|1|500453665|2||-2||4|3|||-2||-2|0|10|||11098|8|||1|146416|40460|4|3|45
502083495|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-26|2011-10-20|Followup|2011-05-26|2011-08-10|Expired|Late||||||||4|4|4|1|4|4|3.5|||||||||3|4|3|3|3|3|3.17||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|3|4|4|3.86||||||4|4|4|4|||||3|3|3||||2|2|||||||Red|Amachi|Volunteer: Lost contact with child/agency|16.8||1|1|2|2|M|Black||18|Yes|Mother|28025|One Parent: Female|Unknown||Yes||Service Organization|General Community|Amachi|Match Support|M|Black||52|28027||Married|Business: Human Resources|28273|0|0|Big Champions|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|502083919|31|0|1|502089653|31|0|1|500453681|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|11|||7461|12|||1|146417|40468|4|0|45
501312033|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-04|2013-02-27|Followup|2011-06-04|2011-07-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Lost interest|32.8||2|2|1|1|F|Black||17|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||35|28226|||Customer Service||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500015820|501312311|31|0|2|502053746|31|0|2|500452835|2||-2||4|3||500000294|-2||-2|0|10|||7464|9|||1|146418||4|1|45
502083504|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-26|2011-10-20|Followup|2011-05-26|2011-08-10|Expired|Late||||||||4|4|4|1|4|4|3.5|||||||||3|3|3|3|4|3|3.17||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Red|Amachi|Volunteer: Lost contact with child/agency|16.8||1|1|2|2|M|Asian||18|Yes|Mother|28025|One Parent: Female|Unknown||Yes||Service Organization|General Community|Amachi|Match Support|M|Black||52|28027||Married|Business: Human Resources|28273|0|0|Big Champions|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|502083919|4|0|1|502089653|31|0|1|500454472|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|11|||7461|12|||1|146419|131834|4|0|45
502180719|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-04|2014-03-20|Followup|2011-06-04|2011-06-30|Complete|Done|4|3|4|2|4|4|3.5|4|2|4|4|4|4|3.67|-4.63|4|4|4|3|4|4|3.83|2|4|4|4|4|4|3.67|4.36|4|4|4|4|3|4|4|3.67|8.99|4|3|2|2|2.75|5|4|4|5|4.5|-38.89|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|2|2|2|2|2|0|2|2|2|2|0||||||Green|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|45.5||2|2|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|Black||42|28273|Masters Degree|Divorced|Business: Marketing||1|6|Michael Baisden|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502181148|31|0|2|502184470|31|0|2|500454904|2||500004772||4|1|500000294, 500004640, 500004901|500000294|-2|500000294|-2|7016|11|||11146|1|||1|146420|134611|4|3|45
502124485|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-28|2011-08-30|Followup|2011-05-28|2011-06-17|Complete|Done|3|1|4|2|4|4|3|4|1|2|1|2|4|2.33|28.76|4|4|4|4|4|4|4|3|4|4|4|4|4|3.83|4.44|4|4|4|4|4|4|4|4|0|5|4|5|5|4.75|5|5|5|5|5|-5|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|4|3|2|4|3|0|2|2|2|2|0||||||Green||Volunteer: Time constraint|15.1||2|2|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|White||32|28206||Single|Medical: Nurse||0|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500008629|502142970|31|0|2|502066586|1|0|2|500454581|2||-2||4|1|||-2||-2|0|4|||7438|1|||1|146421|132622|4|3|45
501622502|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-04|2012-01-31|Followup|2011-06-04|2011-06-13|Complete|Done|3|2|4|1|2|2|2.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Time constraint|19.9||2|2|1|1|M|Black||17|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||32|28210|Bachelors Degree|Single|Tech: Engineer||0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501622822|31|0|1|502162227|1|0|1|500454573|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|146423||4|3|45
500545470|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-01-25|Followup|2011-04-30|2011-06-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|104.9||1|1|1|1|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||34|29708|Bachelors Degree|Single|Self-Employed, Entrepreneur|29708|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501750989|31|0|1|500815012|1|0|1|500173957|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|3|||2238|7|||1|146424||4|1|45
501034365|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-06|2011-02-09|Followup|2010-07-06|2010-09-20|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Health|19.2||2|2|1|1|M|Black||15|Yes|Mother|28216|One Parent: Female|$30,000 to $34,999||No|BBBS National Site|Web Link|General Community|Amachi|Enrollment|M|Black||52|28262|Associate Degree|Married|Finance: Banking||7|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501034638|31|0|1|501580873|31|0|1|500370326|2||-2||4|1|500000294|500000294|-2|500000294|-2|34|2|||7453|7|||1|147497||4|0|45
501994951|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2014-09-18|Followup|2011-06-03|2011-08-02|Declined|Late||||||||3|3|3|1|4|4|3|||||||||4|4|3|4|4|4|3.83||||||4|4|4|4|||||||4|5|5|4|4.5||||||||||4|4|4|3|3|3|3|3.43||||||3|3|3|3|||||3|1|2||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|51.1||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|Unknown||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||36|28078||Single|Customer Service||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501843047|31|0|2|502048623|31|0|2|500455478|2||-2||4|2|||-2||-2|7294|13|||7464|9|||1|147518|139614|4|1|45
501194364|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-27|2011-10-12|Followup|2011-05-27|2011-06-28|Complete|Done|3|2|3|2|3|3|2.67|||||||||3|3|3|4|4|3|3.33|||||||||4|3|3|3.33||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Moved|40.5||1|1|1|1|F|Multi-Race (None of the above)||18|No|Mother|28216|Two Parent|$15,000 to $19,999||Yes||Self|General Community||Enrollment|F|Black||48|28214|Masters Degree|Single|Medical: Doctor, Provider|28207|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501194638|7|0|2|501143598|31|0|2|500265628|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|147738||4|3|45
502210299|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-16|2011-08-01|Baseline|2010-06-15|2010-06-16|Complete|Done|3|2|3|2|2|3|2.5|||||||||2|4|3|3|3|3|3|||||||||3|2|2|2.33||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||1|1|||||||||Green||Volunteer: Moved|13.5||1|1|1|1|M|Hispanic||16|No|Mother|28213|Two Parent: Not Married|Unknown|Y|Yes||School|General Community||RTBM|M|White||39|28209|||Transport: Pilot||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010765|502210728|3|0|1|501993351|1|0|1|500456811|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|147809|-1|4|3|44
502053779|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2012-09-05|Followup|2012-06-15|2012-08-30|Expired|Late||||||||3|3|3|2|3|4|3|||||||||2|3|3|1|2|3|2.33||||||4|4|4|4|||||||3|3|2|4|3||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Red||Child/Family: Feels incompatible with volunteer|26.7||2|2|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community||Match Support|F|Black||39|28216|||Education: College Professor||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|502054203|31|0|2|501912080|31|0|2|500455628|2||-2||4|3|||-2||-2|7295|11|||7464|9|||1|147833|140517|4|0|45
502045258|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-25|2016-08-29|Baseline|2010-06-15|2010-06-25|Complete|Done|4|2|4|1|4|4|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||4|3|3.5|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|74.2||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28262|Bachelors Degree|Single|Medical: Nurse|28262|4|9|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502190790|31|0|2|500457916|2||-2||4|1|||-2||-2|0|10|||6247|12|||1|148107|-1|4|3|44
500872449|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-30|2013-02-28|Followup|2011-05-30|2011-06-05|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|69||1|1|2|2|M|Black||22|No|Mother|28211|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|White||37|28209|Masters Degree|Single|Business: Marketing|28208|1|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500872718|31|0|1|500846955|1|0|1|500178294|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|148464||4|1|45
501994934|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-29|2011-07-29|Baseline|2010-06-16|2010-06-29|Complete|Done|3|3|3|2|3|3|2.83|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Green||Volunteer: Lost contact with child/agency|13||1|1|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||No||BBBS Board/Staff|General Community||Match Support|F|Black||29|28202|||Tech: Production Line||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501843047|31|0|2|501930790|31|0|2|500457779|2||-2||4|1|||-2||-2|0|13|||7464|9|||1|148512|-1|4|3|44
501967613|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2013-02-26|Baseline|2010-06-16|2010-12-31|Complete|Done|4|3|3|3|3|4|3.33|||||||||3|4|3|3|3|2|3|||||||||4|3|3|3.33||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Time constraint|25.9||1|1|1|1|F|Black||20|No|Mother|28273|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Finance: Accountant|28277|3|5|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500012459|501968011|31|0|2|502311344|1|0|2|500498762|2||-2||4|2|||-2|500000294, 500004640|-2|34|2|||7496|10|||1|148519|-1|4|3|44
502173821|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-16|2010-10-25|Baseline|2010-06-16|2010-06-16|Complete|Done|4|1|1|1|4|4|2.5|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1|||||||||Green|Amachi|Volunteer: Time constraint|4.3||2|2|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||30|28205||Married|Child/Day Care Worker||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500010355|502174240|31|0|2|502057248|1|0|2|500457033|2||500003586||4|1|500000294|500000294|-2|500000294|-2|7016|11|||7464|9|||1|148526|-1|4|3|44
502210299|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-16|2011-08-01|Followup|2011-06-15|2011-07-19|Complete|Done|2|4|4|1|4|4|3.17|3|2|3|2|2|3|2.5|26.8|1|4|4|1|1|3|2.33|2|4|3|3|3|3|3|-22.33|4|2|2|2.67|3|2|2|2.33|14.59|4|3|3|4|3.5|3|3|3|3|3|16.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|4|2|3|3|3|3|0|2|2|1|1|100||||||Green||Volunteer: Moved|13.5||1|1|1|1|M|Hispanic||16|No|Mother|28213|Two Parent: Not Married|Unknown|Y|Yes||School|General Community||RTBM|M|White||39|28209|||Transport: Pilot||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010765|502210728|3|0|1|501993351|1|0|1|500456811|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|148558|147809|4|3|45
502114924|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-24|2012-01-27|Baseline|2010-06-16|2010-06-24|Complete|Done|4|1|1|1|1|2|1.67|||||||||1|1|3|1|2|2|1.67|||||||||1|4|3|2.67||||||2|3|4|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|19.1||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||32|28207|Masters Degree|Single|Medical||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|502115351|31|0|2|502019135|1|0|2|500457063|2||-2||4|1|||-2||-2|34|2|||7496|10|||1|148581|-1|4|3|44
502114704|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-20|2012-01-10|Baseline|2010-06-17|2010-08-20|Complete|Done|1|4|2|1|3|3|2.33|||||||||4|4|2|4|4|4|3.67|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||1|1|||||||||Green||Volunteer: Moved|16.7||1|1|1|1|F|Black||18|No|Mother|28270|One Parent: Female|Unknown||Yes|Radio|Media|General Community||RTBM|F|White||32|28204|Masters Degree|Single|Business: Marketing||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502115131|31|0|2|502130736|1|0|2|500460157|2||-2||4|1|||-2||-2|55|1|||7496|10|||1|148929|-1|4|3|44
500934908|BBBS of Greater Charlotte|Main Office|C|Active|2010-06-18|NaT|Followup|2011-06-11|2011-08-02|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||80.9||2|2|1|1|M|Black||16|Yes|Aunt|28216|One Parent: Female|Less than $10,000|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||34|20175|Bachelors Degree|Single|Business: Sales|28211|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|500935173|31|0|1|502107314|1|0|1|500456443|2||500003586||2|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|149641||4|1|45
502142541|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-18|2015-07-23|Followup|2011-06-07|2011-06-17|Complete|Done|4|4|4|4|4|4|4|3|4|4|3|4|4|3.67|8.99|2|4|3|3|2|3|2.83|3|3|3|3|3|3|3|-5.67|4|4|4|4|4|4|4|4|0|4|5|5|4|4.5|4|4|5|3|4|12.5|4|4|4|4|3|4|3|3.71|4|4|4|4|3|4|3|3.71|0|3|4|4|3.67|4|4|4|4|-8.25|1|4|2.5|2|2|2|25|2|2|2|2|0||||||Green||Child: Graduated|61.1||1|1|2|2|F|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502142970|31|0|2|501905673|31|0|2|500455759|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|149723|141478|4|3|45
502070483|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-22|2010-08-24|Baseline|2010-06-18|2010-06-22|Complete|Done|3|4|2|3|2|3|2.83|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||5|1|3|4|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2|||||||||Green||Child/Family: Moved|2.1||1|1|3|3|M|Black||18|Yes|Mother|28269|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|M|Black||45|28262|Bachelors Degree|Married|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500010355|502070907|31|0|1|502087592|31|0|1|500457368|2||500003586||4|1||500000294|-2|500014505, 500015184|-1|34|2|||7462|13|||1|149783|-1|4|3|44
502030263|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2011-03-31|2011-03-10|Complete|Early|4|4|2|2|3|4|3.17|||||||||3|4|4|1|2|4|3|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|3|4|4|4|3.86||||||||||3|4|4|3.67||||||4|3|3.5|||||2|2|||||||||Green|||83.5||1|1|1|1|M|White||15|No|Mother|29710|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community||Match Support|M|White||38|28210|||Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502030662|1|0|1|501923553|1|0|1|500438867|2||-2||2|1|||-2||-2|6855|8|||7464|9|||1|150012||4|3|45
502212598|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2011-07-28|Baseline|2010-06-22|2010-07-22|Complete|Done|4|1|3|3|2|4|2.83|||||||||2|4|4|1|2|3|2.67|||||||||3|4|4|3.67||||||2|3|3|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|Amachi|Volunteer: Moved|12.2||2|2|1|1|F|Black||17|Yes|Mother|28215|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||29|28205|Bachelors Degree|Single|Education: Teacher|28208|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011184|502213028|31|0|2|502068243|1|0|2|500457783|2||-2||4|1|500000294|500000294|-2||-2|7016|11|||7464|9|||1|151061|-1|4|3|44
501955308|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-30|2011-12-15|Baseline|2010-06-22|2010-06-30|Complete|Done|4|2|3|2|3|3|2.83|||||||||2|3|4|3|2|3|2.83|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2|||||||||Red||Volunteer: Moved|17.5||1|1|1|1|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||Yes||School|General Community||RTBM|F|Black||47|28227||Single|Laborer||9|0|New Beginnings Comm.|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500011746|501955706|31|0|2|501734595|31|0|2|500458840|2||-2||4|3|||-2||-2|0|4|||9213|7|||1|151063|-1|4|3|44
502007951|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-28|2010-10-26|Baseline|2010-06-23|2010-06-28|Complete|Done|3|3|3|3|3|4|3.17|||||||||2|3|3|3|2|3|2.67|||||||||3|3|2|2.67||||||4|2|3|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||4|1|2.5|||||1|1|||||||||Red||Volunteer: Lost contact with child/agency|3.9||1|1|1|1|M|Black||20|No|Mother|28216|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|M|Black||27|28215|Some College|Single|Student: College||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500009007|502008350|31|0|1|502201951|31|0|1|500457933|2||-2||4|3|||-2||-2|0|8|||7464|9|||1|151391|-1|4|3|44
501536365|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-03|2014-07-17|Followup|2011-02-03|2011-03-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Time constraint|65.4||1|1|1|1|M|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Enrollment|M|Black||57|28105|Some College|Married|Retail: Sales|28105|10|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501536657|31|0|1|501443152|31|0|1|500336020|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|151770||4|1|45
502114924|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-24|2012-01-27|Followup|2011-06-16|2011-06-28|Declined|Done||||||||4|1|1|1|1|2|1.67|||||||||1|1|3|1|2|2|1.67||||||1|4|3|2.67|||||||2|3|4|3|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|4|3||||2|2|||||||Green||Volunteer: Lost contact with child/agency|19.1||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||32|28207|Masters Degree|Single|Medical||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|502115351|31|0|2|502019135|1|0|2|500457063|2||-2||4|1|||-2||-2|34|2|||7496|10|||1|151830|148581|4|1|45
502045258|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-25|2016-08-29|Followup|2011-06-23|2011-06-01|Complete|Early|2|4|4|4|4|4|3.67|4|2|4|1|4|4|3.17|15.77|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|5|5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|4|4|3.67|-9.26|4|4|4|4|3|3.5|14.29|2|2|2|2|0||||||Green||Volunteer: Lost contact with child/agency|74.2||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28262|Bachelors Degree|Single|Medical: Nurse|28262|4|9|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502190790|31|0|2|500457916|2||-2||4|1|||-2||-2|0|10|||6247|12|||1|152277|148107|4|3|45
501691220|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-02|2012-08-29|Followup|2010-07-02|2010-07-06|Complete|Done|2|3|2|2|2|2|2.17|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green||Child/Family: Moved|37.9||1|1|2|3|M|White||15|No|Mother|27949|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree||Business: Marketing|28031|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501691558|1|0|1|501721806|1|0|1|500367645|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|152475||4|3|45
501987736|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-29|2014-06-18|Followup|2011-06-08|2011-06-12|Complete|Done|3|4|4|4|3|3|3.5|4|4|4|2|4|4|3.67|-4.63|3|3|3|3|4|4|3.33|2|4|4|2|4|4|3.33|0|4|3|3|3.33|4|2|2|2.67|24.72|4|3|5|4|4|4|3|3|3|3.25|23.08|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|3|3.33|20.12|3|4|3.5|2|1|1.5|133.33|2|2|1|1|100||||||Green||Child: Graduated|47.6||1|1|1|1|F|White||20|No|Father|28217|One Parent: Male|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||40|28203|Masters Degree|Single|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501988135|1|0|2|502109789|1|0|2|500456045|2||-2||4|1|||-2||-2|6855|8|||7464|9|||1|153104|142908|4|3|45
501965241|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-29|2012-07-31|Followup|2011-06-22|2011-06-27|Complete|Done|2|4|4|4|4|4|3.67|4|1|4|1|1|1|2|83.5|4|3|4|2|2|4|3.17|1|1|4|4|4|4|3|5.67|4|4|4|4|4|4|4|4|0|5|4|4|5|4.5|4|3|2|3|3|50|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|1|4|2.5|3|3|3|-16.67|2|2|1|1|100||||||Green||Child/Family: Lost contact with volunteer/agency|25.1||1|1|1|1|M|Black||19||Mother|28208|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|M|Black||37|28210||Single|Law||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501578929|31|0|1|502081691|31|0|1|500457757|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|153110|137801|4|3|45
500187077|BBBS of Greater Charlotte|Main Office|C|Completed|2005-05-31|2013-04-02|Followup|2011-05-31|2011-07-11|Complete|Done|3|3|4|4|4|4|3.67|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|2|3|||||2|2|||||||||Green||Child: Graduated|94.1||2|2|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||41|28210|Bachelors Degree|Married|Medical: Pharmacist||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500188224|31|0|1|500189824|1|0|2|500037944|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|153366||4|3|45
500185624|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-28|2013-02-26|Followup|2011-06-28|2011-09-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Moved|68||1|1|1|1|M|Black||16|Yes|Mother|28213|Other/Unknown|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||61|28205||Married|Tech: Management||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|500187258|31|0|1|500923420|31|0|1|500182113|2||500003586||4|2|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|153373||4|0|45
500740293|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2011-06-12|2011-06-29|Complete|Done|3|2|4|2|3|3|2.83|||||||||4|4|4|4|2|3|3.5|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|3|4|4|4|4|4|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Yellow||Child: Lost interest|85||1|1|1|1|M|Black||19||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|Black||39|28216||Single|Transport: Pilot||3|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500876177|31|0|1|500179697|2||-2||4|2|||-2||-2|0|5|||6450|12|||1|153387||4|3|45
501714939|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-03|2012-12-23|Followup|2011-06-03|2011-06-06|Complete|Done|3|2|4|4|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||2|4|2|2.67||||||2|2|2|||||2|2|||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|42.7||1|1|1|1|M|Black||19|Yes|Mother|28105|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||34|28277||Single|Business: Sales|28206|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501715277|31|0|1|501584958|1|0|1|500365824|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|153441||4|3|45
501955308|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-30|2011-12-15|Followup|2011-06-28|2011-06-23|Complete|Done|3|3|3|3|3|3|3|4|2|3|2|3|3|2.83|6.01|4|4|4|3|3|4|3.67|2|3|4|3|2|3|2.83|29.68|4|3|3|3.33|4|4|4|4|-16.75|5|5|5|5|5|4|4|5|4|4.25|17.65|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|3|2.5|4|3|3.5|-28.57|2|2|2|2|0||||||Red||Volunteer: Moved|17.5||1|1|1|1|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||Yes||School|General Community||RTBM|F|Black||47|28227||Single|Laborer||9|0|New Beginnings Comm.|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500011746|501955706|31|0|2|501734595|31|0|2|500458840|2||-2||4|3|||-2||-2|0|4|||9213|7|||1|153977|151063|4|3|45
502221847|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-12|2011-08-23|Baseline|2010-06-30|2010-07-12|Complete|Done|3|1|2|1|4|2|2.17|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|4|3|||||2|2|||||||||Green|Amachi|Volunteer: Lost contact with child/agency|13.4||2|2|1|1|F|Black||16|Yes|GrandMother|28213|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28212|Bachelors Degree|Single|Law|29715|2|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502222278|31|0|2|502103416|31|0|2|500459547|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7496|10|||1|154081|-1|4|3|44
500186107|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-22|2012-10-17|Followup|2011-06-22|2011-07-06|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|5|||||||||4|4|4|4|4|3|3|3.71||||||||||4|4|4|4||||||4|1|2.5|||||2|2|||||||||Green||Child: Graduated|75.9||2|2|1|1|M|Black||22||Mother|28206|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|Black||52|28210|Masters Degree|Married|Business: Mgt, Admin||0|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500012459|500187654|31|0|1|500392161|31|0|1|500102003|2||-2||4|1|||-2||-2|0|10|||2230|7|||1|154140||4|3|45
500185778|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-17|2016-06-23|Followup|2011-06-17|2011-06-16|Complete|Done|3|1|2|2|3|3|2.33|||||||||2|3|3|3|2|3|2.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|4|3.33||||||2|2|2|||||2|2|||||||||Green||Child: Graduated|144.2||1|1|1|1|M|Black||18||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||42|27514||Married|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187368|31|0|1|500188776|1|0|1|500036776|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|154143||4|3|45
502067798|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-09|NaT|Baseline|2010-06-30|2010-07-09|Complete|Done|4|1|1|1|1|4|2|||||||||2|3|4|1|1|4|2.5|||||||||4|4|4|4||||||1|4|5|2|3|||||||3|4|4|4|2|4|3|3.43||||||||||2|2|3|2.33||||||2|4|3|||||2|2|||||||||Green|||80.2||1|1|1|1|M|Black||17|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||52|28270|Bachelors Degree|Married|Business: Mgt, Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|0|1|502062408|1|0|1|500459576|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|154145|-1|4|3|44
500740296|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-25|2011-09-21|Followup|2011-06-25|2011-06-16|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|50.9||2|2|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Therapist/Counselor|General Community||Match Support|F|Black||33|28269|Bachelors Degree|Single|Human Services: Non-Profit||0|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|2|500928282|31|0|2|500181834|2||-2||4|2|||-2||-2|0|5|||7671|13|||1|154182||4|3|45
500740295|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2011-06-12|2011-07-11|Complete|Done|4|4|4|2|3|4|3.5|||||||||4|3|4|4|2|4|3.5|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|2|3|3.57||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Yellow||Volunteer: Feels incompatible with child/family|85||1|1|1|1|M|Black||18||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|White||55|28216|Bachelors Degree|Divorced|Tech: Engineer||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500794907|1|0|1|500179696|2||-2||4|2|||-2||-2|0|5|||46|2|||1|154188||4|3|45
501626226|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-30|2017-03-14|Followup|2011-06-22|2011-06-13|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|2|2|4|2.67|||||||||4|4|4|4||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|80.5||2|2|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||33|28203|High School Graduate|Single|Retail: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501622822|31|0|2|502036832|1|0|2|500457771|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|154319||4|3|45
500545328|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-02|2016-09-30|Followup|2011-07-02|2011-07-07|Complete|Done|3|2|3|2|3|3|2.67|||||||||2|3|3|2|2|3|2.5|||||||||4|4|3|3.67||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Time constraint|99||3|3|1|1|F|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|F|Black||43|28208|Masters Degree|Single|Business: Sales|28078|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|2|501033808|31|0|2|500274449|2||-2||4|1|||-2||-2|0|10|||46|2|||1|154851||4|3|45
500186247|BBBS of Greater Charlotte|Main Office|C|Completed|2005-06-30|2012-09-26|Followup|2011-06-30|2011-07-01|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|3|3|2|3|3|2.83|||||||||3|3|3|3||||||3|2|3|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red||Child: Graduated|86.9||1|1|2|2|M|Black||21||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|M|Black||39|28269|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Site|mentor2.0 2014|RTBM|277|60|598|500000170|500008321|500187842|31|0|1|500189197|31|0|1|500037197|2||-2||4|3|||-2|500014506|-1|0|10|||7464|9|||1|154853||4|3|45
500186645|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-03|2016-01-06|Followup|2011-06-03|2011-06-17|Complete|Done|4|2|4|3|4|4|3.5|||||||||4|4|3|4|2|3|3.33|||||||||4|4|4|4||||||5|3|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2|||||||||Green|Amachi|Child: Graduated|139.1||1|1|1|1|M|Black||18|Yes|Mother|28208|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28256|High School Graduate|Married|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500018987|500188043|31|0|1|500189545|31|0|2|500037636|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|154915||4|3|45
501072636|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-25|2013-06-19|Followup|2011-06-25|2011-07-19|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|3|3|3|3|4|3.17|||||||||3|3|3|3||||||5|3|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Red||Child/Family: Lost contact with volunteer/agency|47.8||2|2|1|1|M|White||18||Mother|28134|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||50|28277|Bachelors Degree|Married|Tech: Management||10|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500004169|500965396|1|0|1|501637727|1|0|1|500368653|2||-2||4|3|||-2|500000294|-2|0|10|||7462|13|||1|154923||4|3|45
501631140|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-17|2016-03-03|Followup|2011-06-17|2011-06-14|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Moved|80.5||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Service: Hotel|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501631463|31|0|1|501628976|1|0|1|500367187|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|154924||4|3|45
501691220|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-02|2012-08-29|Followup|2011-07-02|2011-08-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|37.9||1|1|2|3|M|White||15|No|Mother|27949|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree||Business: Marketing|28031|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501691558|1|0|1|501721806|1|0|1|500367645|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|155093||4|1|45
501609876|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-13|2016-04-29|Followup|2011-07-13|2011-07-12|Complete|Done|2|3|3|4|3|3|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|Project Big|Child: Graduated|81.5||1|2|1|2|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Black||38|28269|Masters Degree|Single|Medical: Nurse|28262|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501610196|31|0|2|501425392|31|0|2|500373716|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7464|9|||1|155177||4|3|45
502165495|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-13|2012-02-28|Baseline|2010-07-07|2010-07-13|Complete|Done|3|4|4|3|3|4|3.5|||||||||3|3|4|4|2|3|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|19.5||1|1|1|1|F|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community||Enrollment|F|White||33|28203|Bachelors Degree|Single|Retail: Sales||2|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|502165924|31|0|2|502087652|1|0|2|500460127|2||-2||4|1|||-2||-2|5635|9|||7464|9|||1|155539|-1|4|3|44
502108064|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2014-02-06|Baseline|2010-07-07|2010-07-22|Complete|Done|3|4|4|4|4|4|3.83|||||||||1|4|3|1|1|3|2.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||1|1|||||||||Yellow||Child: Graduated|42.5||1|1|1|1|F|White||21|No|Father|28277|One Parent: Male|Unknown||No||Relative|General Community||Match Support|F|White||48|28277|High School Graduate|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502108491|1|0|2|502146885|1|0|2|500460150|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|155579|-1|4|3|44
501872144|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-30|NaT|Baseline|2010-07-07|2010-07-30|Complete|Done|4|4|3|1|3|3|3|||||||||2|3|2|1|2|2|2|||||||||2|3|2|2.33||||||2|2|1|2|1.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||1|1|1|||||2|2|||||||||Green|||79.5||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown|Y|Yes||Relative|General Community||Match Support|M|White||35|28205|Masters Degree|Married|Tech: Engineer|28115|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501872517|31|31|1|502063676|1|0|1|500460156|2||-2||2|1|||-2||-2|0|3|||46|2|||1|155585|-1|4|3|44
502173811|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-13|2011-09-02|Baseline|2010-07-08|2010-07-13|Complete|Done|4|2|4|3|4|4|3.5|||||||||2|4|4|4|2|4|3.33|||||||||4|3|3|3.33||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|4|3|||||2|2|||||||||Green|Amachi|Volunteer: Moved|13.7||1|1|2|2|M|Black||20|Yes|Mother|28269|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|RTBM|M|Black||32|28202|Bachelors Degree|Single|Finance: Banking||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011184|502174240|31|0|1|500776552|31|0|1|500460247|2||500003586||4|1|500000294|500000294|-2||-2|7016|11|||46|2|||1|155795|-1|4|3|44
502062624|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-30|2012-12-19|Baseline|2010-07-08|2010-08-30|Complete|Done|3|3|3|2|1|4|2.67|||||||||2|4|3|3|3|4|3.17|||||||||4|4|4|4||||||3|5|3|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Feels incompatible with child/family|27.7||1|1|1|1|F|Black||16|No|Mother|28081|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||32|28083|Bachelors Degree|Single|Tech: Computer/Programmer|28216|1|7|LPL Financial|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|502063048|31|0|2|502067861|31|0|2|500460279|2||-2||4|2|||-2||-2|0|10|||11247|3|||1|155833|-1|4|3|44
502234504|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-28|NaT|Baseline|2010-07-08|2010-07-28|Complete|Done|4|4|4|4|2|4|3.67|||||||||1|4|4|1|2|4|2.67|||||||||4|4|4|4||||||3|3|5|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||1|3|2|||||2|2|||||||||Yellow|Project Big||79.6||1|1|2|2|F|Black||16|No|GrandMother|28208|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|Project Big|Match Support|F|Black||37|28216|Bachelors Degree|Single|Customer Service||8|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500008321|502234935|31|0|2|502129464|31|0|2|500463451|2||500004641||2|2|500004640|500004640|-2||-1|0|4|||11247|3|1204|3|1|155881|-1|4|3|44
502067798|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-09|NaT|Followup|2011-06-30|2011-07-01|Complete|Done|3|3|3|3|3|3|3|4|1|1|1|1|4|2|50|3|3|3|3|3|3|3|2|3|4|1|1|4|2.5|20|3|3|3|3|4|4|4|4|-25|3|3|3|3|3|1|4|5|2|3|0|4|4|4|4|4|4|4|4|3|4|4|4|2|4|3|3.43|16.62|4|4|4|4|2|2|3|2.33|71.67|3|4|3.5|2|4|3|16.67|2|2|2|2|0||||||Green|||80.2||1|1|1|1|M|Black||17|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||52|28270|Bachelors Degree|Married|Business: Mgt, Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|0|1|502062408|1|0|1|500459576|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|156077|154145|4|3|45
502099440|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-23|2012-05-23|Baseline|2010-07-09|2010-07-23|Complete|Done|2|2|3|3|3|3|2.67|||||||||2|3|2|3|3|2|2.5|||||||||4|4|4|4||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||1|3|2|2||||||3|3|3|||||2|2|||||||||Green||Child/Family: Moved|22||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|F|Black||26|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500008629|502099867|31|0|2|502104508|31|0|2|500460403|2||-2||4|1|||-2||-2|0|3|||7496|10|||1|156098|-1|4|3|44
502221847|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-12|2011-08-23|Followup|2011-06-30|2011-06-20|Complete|Done|4|1|2|1|2|2|2|3|1|2|1|4|2|2.17|-7.83|3|4|4|3|4|4|3.67|4|4|4|2|4|4|3.67|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|4|5|5|4.75|5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|4|4|4|2|4|3|33.33|2|2|2|2|0||||||Green|Amachi|Volunteer: Lost contact with child/agency|13.4||2|2|1|1|F|Black||16|Yes|GrandMother|28213|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28212|Bachelors Degree|Single|Law|29715|2|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502222278|31|0|2|502103416|31|0|2|500459547|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7496|10|||1|156393|154081|4|3|45
502240205|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-15|2010-09-10|Baseline|2010-07-12|2010-07-15|Complete|Done|4|2|4|3|3|3|3.17|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|2|3|||||2|2|||||||||Yellow||Volunteer: Time constraint|1.9||3|3|1|1|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||35|28202|Bachelors Degree|Single|Retail: Sales||0|8|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500010355|502240634|31|0|2|502203053|1|0|2|500460610|2||500003586||4|2||500000294|-2|500000294|-2|0|10|||7464|9|||1|156483|-1|4|3|44
502171910|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2015-08-25|Baseline|2010-07-12|2010-07-30|Complete|Done|3|1|2|2|2|3|2.17|||||||||2|3|3|4|2|4|3|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red|Amachi|Volunteer: Time constraint|60.8||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28214|Some College|Married|Medical||3|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502172339|31|0|1|502141964|31|0|1|500460627|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|5|||7464|9|||1|156504|-1|4|3|44
502165495|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-13|2012-02-28|Followup|2011-07-07|2011-07-07|Complete|Done|3|2|3|2|3|3|2.67|3|4|4|3|3|4|3.5|-23.71|3|3|3|2|2|3|2.67|3|3|4|4|2|3|3.17|-15.77|4|3|3|3.33|4|4|4|4|-16.75|3|3|3|3|3|4|4|4|4|4|-25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|3|4|3.5|2|4|3|16.67|2|2|2|2|0||||||Green||Volunteer: Lost contact with child/agency|19.5||1|1|1|1|F|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community||Enrollment|F|White||33|28203|Bachelors Degree|Single|Retail: Sales||2|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|502165924|31|0|2|502087652|1|0|2|500460127|2||-2||4|1|||-2||-2|5635|9|||7464|9|||1|156696|155539|4|3|45
500280148|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-13|NaT|Followup|2011-07-13|2011-07-19|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|3|4|4|4|3.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow|Amachi||80.1||3|3|1|1|F|Black||16|Yes|Mother|28205|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|F|Black||30|28216|Bachelors Degree|Single|Human Services: Non-Profit|28216|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188151|31|0|2|502118494|31|0|2|500460767|2||500003586||2|2|500000294|500000294|-2||-2|0|3|||7464|9|||1|156731||4|3|45
502240203|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-23|2011-07-28|Baseline|2010-07-14|2010-07-23|Complete|Done|4|3|3|2|4|4|3.33|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||5|5|2|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||2|2|||||||||Green|Amachi|Volunteer: Moved|12.2||2|2|1|1|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|RTBM|F|Black||38|28262|Bachelors Degree|Single|Finance: Banking||5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011184|502240634|31|0|2|502110142|31|0|2|500460976|2||||4|1|500000294|500000294|-2|500000294|-2|0|10|||7496|10|||1|157089|-1|4|3|44
502241349|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2013-09-04|Baseline|2010-07-15|2010-07-22|Complete|Done|2|2|2|1|2|2|1.83|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child/Family: Moved|37.5||1|1|2|2|M|Black||19|No|Aunt|28081|Two Parent|Unknown||No|Other|Faith Organization|General Community||Match Support|M|Black||54|28025||Married|Clergy|28025|23|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500002335|502241780|31|0|1|502240986|31|0|1|500461089|2||-2||4|1|||-2|500016374|-2|5635|9|||7671|13|||1|157252|-1|4|3|44
502221899|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2012-06-28|Baseline|2010-07-15|2010-07-22|Complete|Done|3|2|2|2|4|4|2.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|4|2|3|3.5|||||||3|3|3|3|3|3|3|3||||||||||3|3|2|2.67||||||4|4|4|||||1|1|||||||||Green|Amachi|Child: Severity of challenges|23.2||1|1|1|1|F|Black||21|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Arby's|Workplace Partner/Business|General Community||Match Support|F|White||33|28262|Masters Degree|Single|Govt: Mgmt/Admin||5|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|502222330|31|0|2|502188288|1|0|2|500461229|2||-2||4|1|500000294||-2|500000294|-2|3394|14|||7464|9|||1|157469|-1|4|3|44
502222992|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-16|2013-12-12|Baseline|2010-07-16|2010-07-16|Complete|Done|3|3|3|1|2|3|2.5|||||||||2|4|3|2|2|4|2.83|||||||||4|4|3|3.67||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|40.9||1|1|1|1|F|Black||21|No|Aunt|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||32|28213|Bachelors Degree|Single|Education|28223|7|0|BBBS National Site|Web Link|Big|General Site||Enrollment|277|60|598|500000170|500017732|502223423|31|0|2|502085103|31|0|2|500461244|2||-2||4|1|||-2||-1|6854|8|||46|2|||1|157522|-1|4|3|44
502222992|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-16|2013-12-12|Followup|2011-07-16|2011-08-03|Complete|Done|3|2|3|1|4|3|2.67|3|3|3|1|2|3|2.5|6.8|3|3|4|3|4|4|3.5|2|4|3|2|2|4|2.83|23.67|4|4|4|4|4|4|3|3.67|8.99|4|4|3|4|3.75|3|4|4|4|3.75|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|2|2|2|2|0||||||Green||Child: Graduated|40.9||1|1|1|1|F|Black||21|No|Aunt|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||32|28213|Bachelors Degree|Single|Education|28223|7|0|BBBS National Site|Web Link|Big|General Site||Enrollment|277|60|598|500000170|500017732|502223423|31|0|2|502085103|31|0|2|500461244|2||-2||4|1|||-2||-1|6854|8|||46|2|||1|157529|157522|4|3|45
501833031|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2015-11-04|Baseline|2010-07-16|2011-02-28|Complete|Done|3|3|1|4|4|4|3.17|||||||||2|2|3|2|4|4|2.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Moved|56.2||1|1|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28205|Masters Degree|Single|Medical: Doctor, Provider|28277|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502427342|1|0|2|500518294|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|157600|-1|4|3|44
501833026|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-02|2016-09-30|Baseline|2010-07-16|2011-03-02|Complete|Done|2|4|4|3|1|3|2.83|||||||||2|1|3|2|3|2|2.17|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|2|3||||||2|4|3|||||1|1||||4|4||||Yellow|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|67||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28205|Masters Degree|Single|Education: Teacher|2122|1|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502451325|1|0|2|500518305|2||-2||4|2|500005291|500005291|-2|500000294|-2|0|10|||7464|9|||1|157601|-1|4|3|44
500767208|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-03-24|Followup|2011-07-10|2011-06-28|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Project Big|Child: Graduated|68.4||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|Black||32|28216|Masters Degree|Single|Human Services|28215|0|7|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Enrollment|277|60|598|500000170|500017732|500767473|31|0|2|501341042|31|0|2|500276669|2||500004641||4|1|500004640||-2|500014506|-1|0|10|||7671|13|||1|157634||4|3|45
502057402|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-28|2012-10-31|Baseline|2010-07-16|2010-07-27|Complete|Done|4|3|4|4|3|4|3.67|||||||||3|4|3|2|4|1|2.83|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||4|4|4|||||2|2|||||||||Red||Volunteer: Time constraint|27.1||1|1|1|1|M|White||17|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|White||38|28078|Some College|Married|Military||14|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502057826|1|0|1|502196301|1|0|1|500461316|2||-2||4|3|||-2|500000294|-2|0|4|||7496|10|||1|157640|-1|4|3|44
502218269|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2011-04-29|Baseline|2010-07-19|2010-07-30|Blank|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|9||1|1|1|1|F|Black||17|Yes|Mother|28203|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Enrollment|F|White||27|28262||Single|Service: Restaurant||1|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502218700|31|0|2|502083213|1|0|2|500461413|2||-2||4|1|500000294|500000294|-2||-2|7016|11|||7496|10|||1|157855|-1|4|3|44
502015842|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-21|2011-10-26|Baseline|2010-07-19|2010-07-21|Complete|Done|3|2|2|1|2|2|2|||||||||3|2|4|3|3|4|3.17|||||||||4|4|4|4||||||5|3|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2|||||||||Green|Amachi|Volunteer: Lost contact with child/agency|15.2||1|1|1|1|M|Black||17|Yes|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|RTBM|M|White||35|28211|Bachelors Degree|Single|Finance||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|502016241|31|0|1|502160380|1|0|1|500461467|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|157993|-1|4|3|44
502179379|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-25|2015-07-31|Baseline|2010-07-20|2010-07-25|Complete|Done|4|4|4|4|2|4|3.67|||||||||1|4|4|1|2|4|2.67|||||||||4|4|4|4||||||3|3|5|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||1|2|1.5|||||2|2|||||||||Red|Project Big|Volunteer: Lost contact with child/agency|60.2||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|Black||34|28269||Single|Student: College||0|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|502179808|31|0|2|502161458|31|0|2|500461681|2||-2||4|3|500004640|500004640|-2||-2|0|10|||9221|5|||1|158340|-1|4|3|44
502227959|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-23|2010-10-06|Baseline|2010-07-21|2010-07-23|Complete|Done|4|1|4|1|3|3|2.67|||||||||2|1|3|2|4|3|2.5|||||||||4|4|3|3.67||||||3|4|2|3|3|||||||4|4|4|4|3|4|2|3.57||||||||||3|4|3|3.33||||||3|3|3|||||1|1|||||||||Red||Volunteer: Unrealistic expectations|2.5||1|1|1|1|M|Black||18|No|GrandMother|28036|Grandparents|Unknown||Yes||Relative|General Community||Match Support|M|White||56|28031|High School Graduate|Married|Consultant|28031|25|0|BFKS|Special Event|Big|General Community||Match Support|277|60|598|500000170|500009007|502228390|31|0|1|502198861|1|0|1|500462034|2||-2||4|3|||-2||-2|0|3|||7454|8|||1|158674|-1|4|3|44
502015842|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-21|2011-10-26|Followup|2011-07-21|2011-10-05|Expired|Late||||||||3|2|2|1|2|2|2|||||||||3|2|4|3|3|4|3.17||||||4|4|4|4|||||||5|3|5|4|4.25||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||3|4|3.5||||2|2|||||||Green|Amachi|Volunteer: Lost contact with child/agency|15.2||1|1|1|1|M|Black||17|Yes|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|RTBM|M|White||35|28211|Bachelors Degree|Single|Finance||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|502016241|31|0|1|502160380|1|0|1|500461467|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|158722|157993|4|0|45
501253195|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-24|NaT|Followup|2010-10-24|2010-11-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||100.7||1|1|2|2|M|Black||15|Yes|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28203|Masters Degree|Single|Medical: Doctor, Provider|28211|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501253471|31|0|1|500395148|1|0|1|500282924|2||500003586||2|1|500000294||-2||-2|0|10|||7464|9|||1|158833||4|1|45
502241349|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2013-09-04|Followup|2011-07-22|2011-10-06|Expired|Late||||||||2|2|2|1|2|2|1.83|||||||||2|3|3|3|3|3|2.83||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Child/Family: Moved|37.5||1|1|2|2|M|Black||19|No|Aunt|28081|Two Parent|Unknown||No|Other|Faith Organization|General Community||Match Support|M|Black||54|28025||Married|Clergy|28025|23|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500002335|502241780|31|0|1|502240986|31|0|1|500461089|2||-2||4|1|||-2|500016374|-2|5635|9|||7671|13|||1|158866|157252|4|0|45
500969481|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-22|2011-10-13|Followup|2011-07-22|2011-08-03|Complete|Done|3|2|3|1|2|3|2.33|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2|||||||||Yellow|Project Big|Child/Family: Lost contact with volunteer/agency|38.7||1|1|2|2|F|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|No||Therapist/Counselor|General Community||Match Support|F|Black||41|28209|Bachelors Degree|Single|Finance: Banking|28255|0|6|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500011639|500969749|31|0|2|501202092|31|0|2|500274109|2||-2||4|2|500004640||-2||-2|0|5|||130|1|||1|158913||4|3|45
500732462|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-18|2012-02-28|Followup|2011-07-18|2011-08-01|Complete|Done|3|3|3|2|3|3|2.83|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|55.4||1|1|1|1|F|Black||22||Mother|28205|One Parent: Female|$30,000 to $34,999|Y|No||School|General Community||Match Support|F|Black||40|28269|Masters Degree|Single|Education: Admin|28223|1|9|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500732729|31|0|2|500878773|31|0|2|500184327|2||-2||4|1|||-2||-2|0|4|||7458|9|||1|158955||4|3|45
502108064|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2014-02-06|Followup|2011-07-22|2011-09-06|Declined|Late||||||||3|4|4|4|4|4|3.83|||||||||1|4|3|1|1|3|2.17||||||4|4|4|4|||||||5|5|5|5|5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||1|1|1||||1|1|||||||Yellow||Child: Graduated|42.5||1|1|1|1|F|White||21|No|Father|28277|One Parent: Male|Unknown||No||Relative|General Community||Match Support|F|White||48|28277|High School Graduate|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502108491|1|0|2|502146885|1|0|2|500460150|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|159085|155579|4|1|45
500896588|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2016-06-15|Followup|2011-07-20|2011-07-19|Complete|Done|3|3|4|3|4|4|3.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|3|3.33||||||3|1|2|||||2|2|||||||||Green||Child: Graduated|106.9||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28273|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||36|28269|Masters Degree|Married|Education|28205|6|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|500896858|3|15|2|500924445|1|0|2|500183434|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|159118||4|3|45
502221899|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2012-06-28|Followup|2011-07-22|2011-09-06|Declined|Late||||||||3|2|2|2|4|4|2.83|||||||||3|4|4|3|3|4|3.5||||||4|4|4|4|||||||5|4|2|3|3.5||||||||||3|3|3|3|3|3|3|3||||||3|3|2|2.67|||||4|4|4||||1|1|||||||Green|Amachi|Child: Severity of challenges|23.2||1|1|1|1|F|Black||21|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Arby's|Workplace Partner/Business|General Community||Match Support|F|White||33|28262|Masters Degree|Single|Govt: Mgmt/Admin||5|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|502222330|31|0|2|502188288|1|0|2|500461229|2||-2||4|1|500000294||-2|500000294|-2|3394|14|||7464|9|||1|159196|157469|4|1|45
500881634|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-14|NaT|Followup|2011-07-14|2011-09-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||104||1|2|1|2|M|Black||18||Mother|28213|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||38|28213||Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500881903|31|0|1|500816190|31|0|2|500277615|2||-2||2|1|||-2||-2|0|4|||46|2|||1|159252||4|1|45
502099440|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-23|2012-05-23|Followup|2011-07-23|2011-09-06|Declined|Done||||||||2|2|3|3|3|3|2.67|||||||||2|3|2|3|3|2|2.5||||||4|4|4|4|||||||3|2|4|4|3.25||||||||||4|4|4|4|4|4|4|4||||||1|3|2|2|||||3|3|3||||2|2|||||||Green||Child/Family: Moved|22||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|F|Black||26|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500008629|502099867|31|0|2|502104508|31|0|2|500460403|2||-2||4|1|||-2||-2|0|3|||7496|10|||1|159255|156098|4|1|45
500809082|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-01|2012-03-13|Followup|2011-06-01|2011-06-03|Complete|Done|2|1|4|4|4|4|3.17|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Yellow||Child: Graduated|57.4||1|1|1|1|M|Black||23||Mother|28210|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|White||34|28203|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||RTBM|277|60|598|500000170|500011746|500809351|31|0|1|500878459|1|0|1|500178590|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|159260||4|3|45
502157842|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-23|2011-10-13|Baseline|2010-07-23|2010-07-23|Complete|Done|4|1|1|1|4|2|2.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Time constraint|14.7||1|1|2|2|F|Black||16|No|Mother|28205|One Parent: Female|$15,000 to $19,999||Yes||Relative|General Community||Enrollment|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011639|502158281|31|0|2|502204211|31|0|2|500462416|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|159280|-1|4|3|44
502157842|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-23|2011-10-13|Followup|2011-07-23|2011-08-09|Complete|Done|4|2|4|2|4|4|3.33|4|1|1|1|4|2|2.17|53.46|3|3|3|2|3|3|2.83|4|4|4|4|4|4|4|-29.25|4|4|4|4|4|4|4|4|0|3|3|3|3|3|5|4|5|5|4.75|-36.84|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|2|2|0|4|4||||Green||Volunteer: Time constraint|14.7||1|1|2|2|F|Black||16|No|Mother|28205|One Parent: Female|$15,000 to $19,999||Yes||Relative|General Community||Enrollment|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011639|502158281|31|0|2|502204211|31|0|2|500462416|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|159329|159280|4|3|45
502137968|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-08|2013-01-08|Baseline|2010-07-23|2011-03-08|Complete|Done|3|4|3|1|3|4|3|||||||||3|3|4|3|2|4|3.17|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|22.1||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||41|28078|Bachelors Degree|Married|Govt|28262|7|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500011746|502138397|31|0|1|502417993|1|0|1|500521032|2||-2||4|3|500005291|500005291|-2|500000294, 500004640|-2|34|2|||7464|9|||1|159363|-1|4|3|44
502139829|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-12|2013-08-08|Baseline|2010-07-23|2010-08-12|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|3|2|4|3.17|||||||||4|3|4|3.67||||||5|4|4|4|4.25|||||||4|4|4|4|3|3|3|3.57||||||||||4|4|3|3.67||||||4|2|3|||||2|2|||||||||Red||Volunteer: Lost contact with child/agency|35.9||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||30|28226|Masters Degree|Single|Finance: Accountant||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502140258|31|0|1|502178005|1|0|1|500462499|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|159370|-1|4|3|44
502064627|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-20|NaT|Baseline|2010-07-23|2010-08-20|Complete|Done|2|2|4|2|3|4|2.83|||||||||3|3|4|3|2|4|3.17|||||||||4|3|2|3||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|2|3|2.67||||||2|3|2.5|||||1|1|||||||||Green|||78.9||1|1|2|2|M|Black||16|No|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|502065051|31|0|1|500773055|3|14|1|500462574|2||-2||2|1|||-2||-2|0|10|||46|2|||1|159373|-1|4|3|44
502179379|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-25|2015-07-31|Followup|2011-07-20|2011-07-27|Complete|Done|3|3|2|1|4|3|2.67|4|4|4|4|2|4|3.67|-27.25|3|4|4|1|3|4|3.17|1|4|4|1|2|4|2.67|18.73|4|4|4|4|4|4|4|4|0|5|3|5|5|4.5|3|3|5|5|4|12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|4|3.67|3|4|4|3.67|0|4|4|4|1|2|1.5|166.67|2|2|2|2|0||||||Red|Project Big|Volunteer: Lost contact with child/agency|60.2||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|Black||34|28269||Single|Student: College||0|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|502179808|31|0|2|502161458|31|0|2|500461681|2||-2||4|3|500004640|500004640|-2||-2|0|10|||9221|5|||1|159519|158340|4|3|45
500478936|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-14|2013-11-11|Followup|2011-07-14|2011-07-15|Complete|Done|3|4|4|3|3|3|3.33|||||||||3|4|3|2|3|3|3|||||||||4|3|4|3.67||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Green||Child: Graduated|63.9||1|1|3|3|M|Black||21|No|Mother|28078|One Parent: Female|$25,000 to $29,999||No||Neighbor/Friend|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|500479187|31|0|1|501284751|31|0|1|500275964|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|8|||132|8|||1|159573||4|3|45
502185074|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-16|2011-03-21|Baseline|2010-07-26|2010-08-13|Complete|Done|1|2|1|4|1|1|1.67|||||||||3|1|3|1|1|1|1.67|||||||||4|4|4|4||||||3|2|4|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||2|3|2|2.33||||||2|2|2|||||2|2|||||||||Yellow||Volunteer: Time constraint|7.1||2|2|1|1|F|Black||18|No|GrandMother|28208|Grandparents|Unknown||Yes|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28270|Bachelors Degree|Single|Medical: Nurse|28203|3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500011639|502185503|31|0|2|502189418|31|0|2|500462607|2||-2||4|2||500005291|-2||-2|5635|9|||131|1|||1|159621|-1|4|3|44
500186952|BBBS of Greater Charlotte|Main Office|C|Active|2004-07-15|NaT|Followup|2011-07-15|2011-07-06|Complete|Done|4|1|3|1|4|4|2.83|||||||||1|2|4|1|3|4|2.5|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|4|2.5|||||2|2|||||||||Green|Amachi||152||1|1|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||73|28203||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|500188132|31|0|2|500189723|1|0|2|500037836|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|159638||4|3|45
502145270|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2011-10-26|Baseline|2010-07-26|2010-07-30|Complete|Done|3|4|2|1|1|4|2.5|||||||||2|4|3|2|1|3|2.5|||||||||4|3|4|3.67||||||3|4|5|4|4|||||||4|2|4|4|4|4|3|3.57||||||||||4|4|3|3.67||||||1|1|1|||||1|1|||||||||Green||Child/Family: Lost contact with volunteer/agency|14.9||1|1|2|2|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|F|Black||39|28262|Masters Degree|Single|Human Services: Psychologist||3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502145699|31|0|2|500189131|31|0|2|500462648|2||-2||4|1|||-2||-2|0|8|||7496|10|||1|159664|-1|4|3|44
500835156|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2016-11-10|Followup|2011-07-10|2011-07-18|Complete|Done|4|2|4|4|4|4|3.67|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child/Family: Lost contact with volunteer/agency|100||1|2|1|2|M|Black||17||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Multi-Race (None of the above)||38|29710|Bachelors Degree|Single|Architect||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500835425|31|0|1|500466903|7|0|1|500277232|2||-2||4|1|||-2||-2|0|4|||46|2|||1|159993||4|3|45
502057402|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-28|2012-10-31|Followup|2011-07-16|2011-08-03|Complete|Done|3|2|3|2|3|2|2.5|4|3|4|4|3|4|3.67|-31.88|3|3|3|2|2|3|2.67|3|4|3|2|4|1|2.83|-5.65|4|3|3|3.33|4|4|4|4|-16.75|3|3|2|3|2.75|5|4|4|4|4.25|-35.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3.67|8.99|3|3|3|4|4|4|-25|2|2|2|2|0||||||Red||Volunteer: Time constraint|27.1||1|1|1|1|M|White||17|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|White||38|28078|Some College|Married|Military||14|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502057826|1|0|1|502196301|1|0|1|500461316|2||-2||4|3|||-2|500000294|-2|0|4|||7496|10|||1|160459|157640|4|3|45
502173588|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2012-08-30|Baseline|2010-07-28|2010-08-27|Complete|Done|3|1|2|1|3|3|2.17|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||2|2|2|1|1|2|1|1.57||||||||||4|4|4|4||||||2|1|1.5|||||1|1|||||||||Yellow|Amachi|Volunteer: Lost contact with child/agency|24.1||2|2|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||No|A Child's Place|Service Organization|General Community|Amachi|Enrollment|F|White||29|28217|Bachelors Degree|Single|Customer Service||5|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502174017|31|0|2|502085998|1|0|2|500463449|2||500003586||4|2|500000294|500000294|-2||-2|7016|11|||7496|10|||1|160541|-1|4|3|44
502234504|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-28|NaT|Followup|2011-07-28|2011-08-23|Complete|Done|4|1|4|1|4|4|3|4|4|4|4|2|4|3.67|-18.26|2|4|2|1|1|4|2.33|1|4|4|1|2|4|2.67|-12.73|4|4|4|4|4|4|4|4|0|2|3|2|2|2.25|3|3|5|5|4|-43.75|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|3|4|4|3.67|8.99|2|2|2|1|3|2|0|2|2|2|2|0|4|4||||Yellow|Project Big||79.6||1|1|2|2|F|Black||16|No|GrandMother|28208|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|Project Big|Match Support|F|Black||37|28216|Bachelors Degree|Single|Customer Service||8|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500008321|502234935|31|0|2|502129464|31|0|2|500463451|2||500004641||2|2|500004640|500004640|-2||-1|0|4|||11247|3|1204|3|1|160584|155881|4|3|45
501868351|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-16|2011-01-19|Baseline|2010-07-29|2010-08-16|Complete|Done|3|1|2|2|1|3|2|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|3|4|3.86||||||||||1|1|1|1||||||2|2|2|||||1|1|||||||||Green||Volunteer: Time constraint|5.1||2|2|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|F|Black||34|28205|Masters Degree|Single|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501868724|31|0|2|502163779|31|0|2|500463602|2||-2||4|1||500005291|-2||-2|0|10|||7464|9|||1|160870|-1|4|3|44
501614157|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-29|2013-04-04|Followup|2011-07-29|2011-09-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|44.2||1|1|1|1|F|Black||21|No|Mother|28202|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28273|||Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|501614477|31|0|2|501596246|31|0|2|500374258|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|160876||4|1|45
501444237|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-29|2011-10-13|Followup|2011-07-29|2011-08-09|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|14.5||3|3|1|1|M|Black||17||GrandMother|28215|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|Black||36|28213|Associate Degree|Single|Retail: Sales||3|6|Michael Baisden|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011639|501444522|31|0|1|502183206|31|0|1|500461448|2||-2||4|3|||-2|500000294|-2|0|10|||11146|1|||1|160965||4|1|45
502183055|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2012-06-30|Baseline|2010-07-30|2010-07-30|Complete|Done|3|3|3|2|2|2|2.5|||||||||3|4|3|3|3|4|3.33|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|3|3|||||1|1|||||||||Red||Volunteer: Lost contact with child/agency|23||1|1|2|2|F|Black||18|No|Mother|28226|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||35|28270|Bachelors Degree|Single|Human Services: Social Worker||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|502183484|31|0|2|501035952|31|0|2|500463671|2||-2||4|3|||-2||-2|0|10|||46|2|||1|161032|-1|4|3|44
502183055|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2012-06-30|Followup|2011-07-30|2011-08-09|Declined|Done||||||||3|3|3|2|2|2|2.5|||||||||3|4|3|3|3|4|3.33||||||4|4|4|4|||||||4|5|4|5|4.5||||||||||4|4|4|4|4|4|3|3.86||||||3|3|3|3|||||3|3|3||||1|1|||||||Red||Volunteer: Lost contact with child/agency|23||1|1|2|2|F|Black||18|No|Mother|28226|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||35|28270|Bachelors Degree|Single|Human Services: Social Worker||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|502183484|31|0|2|501035952|31|0|2|500463671|2||-2||4|3|||-2||-2|0|10|||46|2|||1|161035|161032|4|1|45
502057399|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-02|2011-01-13|Baseline|2010-07-30|2010-08-02|Complete|Done|4|3|4|3|2|4|3.33|||||||||3|3|2|3|3|3|2.83|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|1|2.5|||||2|2|||||||||Green||Volunteer: Time constraint|5.4||2|2|1|1|M|White||20|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28031||Single|Finance||0|0|Recruitment Event|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011639|502057823|1|0|1|502102663|1|0|1|500463696|2||-2||4|1||500005291|-2|500000294|-2|0|4|||7458|9|||1|161076|-1|4|3|44
501872144|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-30|NaT|Followup|2011-07-30|2011-09-01|Complete|Done|4|2|4|3|4|4|3.5|4|4|3|1|3|3|3|16.67|3|4|4|1|3|3|3|2|3|2|1|2|2|2|50|4|4|3|3.67|2|3|2|2.33|57.51|4|3|3|3|3.25|2|2|1|2|1.75|85.71|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|4|3.67|4|4|3|3.67|0|4|4|4|1|1|1|300|2|2|2|2|0|4|4||||Green|||79.5||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown|Y|Yes||Relative|General Community||Match Support|M|White||35|28205|Masters Degree|Married|Tech: Engineer|28115|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501872517|31|31|1|502063676|1|0|1|500460156|2||-2||2|1|||-2||-2|0|3|||46|2|||1|161132|155585|4|3|45
500186352|BBBS of Greater Charlotte|Main Office|C|Completed|2002-07-29|2014-01-02|Followup|2011-07-29|2011-07-29|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|5|3|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child: Graduated|137.2||4|4|2|2|M|Black||21||Mother|28212|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|White||45|28226|Masters Degree|Married|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500187945|31|0|1|500189280|1|0|1|500037290|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|161211||4|3|45
501402710|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-19|2015-06-17|Followup|2011-06-19|2011-06-30|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|4|3|3|3|4|3.17|||||||||4|4|4|4||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Green||Child/Family: Moved|71.9||1|1|1|1|M|Black||18|No|Mother|30058|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28215||Married|Consultant|28285|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501402995|31|0|1|501728845|1|0|1|500368860|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|161219||4|3|45
502145270|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2011-10-26|Followup|2011-07-30|2011-10-14|Expired|Late||||||||3|4|2|1|1|4|2.5|||||||||2|4|3|2|1|3|2.5||||||4|3|4|3.67|||||||3|4|5|4|4||||||||||4|2|4|4|4|4|3|3.57||||||4|4|3|3.67|||||1|1|1||||1|1|||||||Green||Child/Family: Lost contact with volunteer/agency|14.9||1|1|2|2|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|F|Black||39|28262|Masters Degree|Single|Human Services: Psychologist||3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502145699|31|0|2|500189131|31|0|2|500462648|2||-2||4|1|||-2||-2|0|8|||7496|10|||1|161239|159664|4|0|45
502171910|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2015-08-25|Followup|2011-07-12|2011-07-18|Complete|Done|3|1|2|1|1|1|1.5|3|1|2|2|2|3|2.17|-30.88|2|2|1|2|3|3|2.17|2|3|3|4|2|4|3|-27.67|3|4|4|3.67|4|4|4|4|-8.25|4|5|2|3|3.5|4|3|4|3|3.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|4|3.67|4|4|4|4|-8.25|2|2|2|4|4|4|-50|2|2|2|2|0||||||Red|Amachi|Volunteer: Time constraint|60.8||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28214|Some College|Married|Medical||3|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502172339|31|0|1|502141964|31|0|1|500460627|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|5|||7464|9|||1|161269|156504|4|3|45
500910037|BBBS of Greater Charlotte|Main Office|C|Active|2009-06-22|NaT|Followup|2011-06-22|2011-08-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||92.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||46|28277||Married|Business: Mgt, Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|500910307|31|0|1|500856100|1|0|1|500368834|2||-2||2|1|||-2||-2|0|10|||46|2|||1|166251||4|1|45
502247430|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-17|2014-01-23|Baseline|2010-08-02|2010-08-17|Complete|Done|3|1|1|1|2|3|1.83|||||||||2|2|3|1|2|2|2|||||||||4|3|3|3.33||||||2|3|2|4|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|4|3.33||||||2|1|1.5|||||1|1|||||||||Yellow||Child: Lost interest|41.2||1|1|1|1|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||63|28078|Bachelors Degree|Married|Medical: Nurse||10|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502247861|31|0|2|502226106|1|0|2|500465539|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|166252|-1|4|3|44
500395038|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-01|2015-02-20|Followup|2011-08-01|2011-07-18|Complete|Done|4|4|4|4|3|3|3.67|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||5|5|3|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Child: Graduated|102.7||1|1|1|1|M|White||20||Mother|28226|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|M|White||39|28211|Masters Degree|Married|Law: Lawyer|28204|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500395288|1|0|1|500392006|1|0|1|500104016|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|166437||4|3|45
500934906|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-31|2013-02-12|Followup|2011-07-31|2011-09-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Lost contact with child/agency|66.5||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||52|28216|Bachelors Degree|Married|Tech: Engineer||13|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500935173|31|0|2|500859806|31|0|2|500186448|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|166716||4|1|45
501318837|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-04|2013-02-27|Followup|2011-08-04|2011-08-23|Complete|Done|1|2|2|2|2|4|2.17|||||||||3|2|4|2|4|4|3.17|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Time constraint|30.8||2|2|1|1|M|Black||17|No|Mother|28205|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Retail: Sales||0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|501319115|31|0|1|502170420|1|0|1|500459741|2||-2||4|3|||-2||-2|6854|8|||7496|10|||1|166723||4|3|45
502221904|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-06|2013-01-31|Baseline|2010-08-05|2010-08-06|Complete|Done|3|1|2|1|4|3|2.33|||||||||1|1|2|1|2|2|1.5|||||||||4|4|4|4||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||2|4|1|2.33||||||3|3|3|||||2|2|||||||||Red|Amachi|Child/Family: Infraction of match rules/agency policies|29.9||1|1|3|3|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Arby's|Workplace Partner/Business|General Community||Match Support|F|Black||36|28078|Masters Degree|Married|Business: Marketing|28273|1|1|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|277|60|598|500000170|500015820|502222335|31|0|2|502056302|31|0|2|500464397|2||500003586||4|3|500000294||-2|500014505, 500014506|-1|3394|14|||7671|13|||1|167141|-1|4|3|44
501726201|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2015-01-30|Followup|2011-07-08|2011-07-31|Complete|Done|3|2|2|1|2|3|2.17|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2|||||||||Red|Amachi|Child/Family: Moved|66.8||1|1|1|1|F|Black||17|Yes|Mother|28212|One Parent: Female|Unknown||Yes|YeaGod|Faith Organization|General Community|Amachi|Match Support|F|Black||51|28262|PHD|Married|Real Estate: Realtor||0|0|Weeping Willow|Faith Organization|Big|General Community||Enrollment|277|60|598|500000170|500008321|501726541|31|0|2|501734664|31|0|2|500371036|2||-2||4|3|500000294|500000294|-2||-2|5634|9|||9218|7|||1|167309||4|3|45
502221904|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-06|2013-01-31|Followup|2011-08-05|2011-08-04|Complete|Done|3|2|3|1|3|2|2.33|3|1|2|1|4|3|2.33|0|2|3|3|3|3|3|2.83|1|1|2|1|2|2|1.5|88.67|4|3|3|3.33|4|4|4|4|-16.75|3|3|3|3|3|2|2|3|3|2.5|20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|2|4|1|2.33|71.67|3|3|3|3|3|3|0|2|2|2|2|0||||||Red|Amachi|Child/Family: Infraction of match rules/agency policies|29.9||1|1|3|3|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Arby's|Workplace Partner/Business|General Community||Match Support|F|Black||36|28078|Masters Degree|Married|Business: Marketing|28273|1|1|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|277|60|598|500000170|500015820|502222335|31|0|2|502056302|31|0|2|500464397|2||500003586||4|3|500000294||-2|500014505, 500014506|-1|3394|14|||7671|13|||1|167437|167141|4|3|45
500363212|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-24|2012-11-27|Followup|2011-05-24|2011-06-30|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|4|3|3|4|3.5|||||||||4|3|3|3.33||||||4|4|4|4|4|||||||4|4|4|3|3|3|3|3.43||||||||||4|3|3|3.33||||||3|2|2.5|||||2|2|||||||||Green|Amachi|Volunteer: Moved|66.2||2|2|1|1|F|Multi-Race (None of the above)||16||Mother|28025|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||34|28211|Associate Degree|Living w/ Significant Other|Business: Clerical|28211|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188099|7|0|2|500797130|1|0|2|500176231|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|167613||4|3|45
500186953|BBBS of Greater Charlotte|Main Office|C|Completed|2004-05-25|2012-08-09|Followup|2011-05-25|2011-06-30|Complete|Done|3|3|3|2|4|4|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.5||1|1|2|2|M|Black||18|Yes|GrandMother|28214|Other Relative|Unknown||No||Self|General Community|Amachi|Match Support|M|White||45|28207||Single|Unknown|28209|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188126|31|0|1|500189724|1|0|1|500037838|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|167959||4|3|45
500408135|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-25|2015-01-30|Followup|2011-05-25|2011-06-05|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|104.2||1|1|4|4|F|Black||19|Yes|Mother|28083|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500008321|500408385|31|0|2|500189709|31|0|2|500099932|2||500003586||4|1|500000294|500000294|-2|500000294, 500016374|-2|6854|8|||2230|7|||1|167965||4|1|45
501631059|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-26|2012-09-10|Followup|2011-05-26|2011-07-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|39.5||1|1|1|1|F|Black||18|No|Mother|28202|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||29|28216|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501631382|31|0|2|501589359|31|0|2|500364875|2||-2||4|2|||-2|500000294|-2|34|2|||7464|9|||1|168265||4|1|45
501919692|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-13|2012-03-30|Baseline|2010-08-10|2010-08-13|Complete|Done|3|3|3|3|3|4|3.17|||||||||4|1|1|2|4|4|2.67|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Red||Volunteer: Lost contact with child/agency|19.5||1|1|1|1|M|White||16|No|Mother|28270|One Parent: Female|Unknown||No||Self|General Community||Enrollment|M|White||35|28270|Associate Degree|Married|Firefighter||1|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013709|501920088|1|0|1|502219683|1|0|1|500465111|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|168273|-1|4|3|44
502233625|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-13|2011-01-20|Baseline|2010-08-10|2010-08-13|Complete|Done|3|3|3|2|1|3|2.5|||||||||2|3|3|3|4|3|3|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Child/Family: Unrealistic expectations|5.3||3|3|1|1|F|Multi-race (Hispanic & White)||17|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||31|28269|Bachelors Degree|Single|Finance||3|0|Self|Self|Big|General Community||RTBM|277|60|598|500000170|500011639|502234056|35|0|2|502228626|31|0|2|500465112|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|168274|-1|4|3|44
502233621|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-14|2013-04-25|Baseline|2010-08-10|2010-08-13|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|1|4|2|4|4|3.17|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Child/Family: Moved|32.4||1|1|2|2|M|Multi-race (Hispanic & White)||16|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction|28208|1|1|Igniting Breakfast|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500011746|502234052|35|0|1|502255664|1|0|1|500465113|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17266|8|||1|168275|-1|4|3|44
501228176|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-05|2013-08-13|Followup|2011-08-05|2011-07-18|Complete|Early|3|4|4|3|3|4|3.5|||||||||2|3|4|4|3|4|3.33|||||||||4|4|4|4||||||4|3|3|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|4|3.5|||||2|2|||||||||Red||Volunteer: Lost contact with child/agency|60.3||1|1|1|1|M|Black||20|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|28078|Masters Degree|Married|Finance: Auditor|28202|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|501228452|31|0|1|501279790|1|0|1|500279399|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|168648||4|3|45
502193174|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-18|2011-12-28|Baseline|2010-08-11|2010-08-18|Complete|Done|4|1|1|4|2|4|2.67|||||||||1|3|3|2|3|3|2.5|||||||||4|4|4|4||||||4|2|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Lost contact with child/agency|16.3||2|2|1|1|M|Black||16||Mother|28273|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|Black||49|28277|Associate Degree|Married|Tech: Engineer||0|9|Recruitment Event|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|502193603|31|0|1|502187342|31|0|1|500465373|2||-2||4|1|||-2|500000294|-2|0|4|||7443|2|||1|168695|-1|4|3|44
502139829|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-12|2013-08-08|Followup|2011-08-12|2011-08-09|Complete|Done|4|3|4|4|3|4|3.67|3|4|4|4|4|4|3.83|-4.18|2|4|3|3|3|3|3|2|4|4|3|2|4|3.17|-5.36|4|3|4|3.67|4|3|4|3.67|0|4|4|3|2|3.25|5|4|4|4|4.25|-23.53|4|4|4|4|3|1|2|3.14|4|4|4|4|3|3|3|3.57|-12.04|3|3|4|3.33|4|4|3|3.67|-9.26|3|3|3|4|2|3|0|2|2|2|2|0|4|4||||Red||Volunteer: Lost contact with child/agency|35.9||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||30|28226|Masters Degree|Single|Finance: Accountant||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502140258|31|0|1|502178005|1|0|1|500462499|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|169012|159370|4|3|45
500892907|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-29|2012-09-11|Followup|2011-05-29|2011-05-30|Complete|Done|3|4|4|4|3|1|3.17|||||||||2|4|3|3|2|4|3|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|2|2|||||2|2|||||||||Red|Amachi|Child: Graduated|51.4||1|1|3|3|F|Black||22|No|Mother|28216|One Parent: Female|Unknown||No||Faith Organization|General Community|Amachi|Match Support|F|Hispanic||37|28203|Some College|Single|Education: Teacher|28217|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500893173|31|0|2|500188541|3|0|2|500268211|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|169208||4|3|45
500892903|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-29|2012-12-23|Followup|2011-05-29|2011-05-28|Complete|Done|3|4|4|4|4|3|3.67|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||5|2|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|1|2|||||2|2|||||||||Yellow|Amachi|Child: Graduated|54.8||1|1|1|1|F|Black||22|Yes|Mother|28216|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||36|28273|Juris Doctorate (JD)|Single|Law: Lawyer|28052|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500893173|31|0|2|501189856|31|0|2|500268753|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|169211||4|3|45
500910040|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2014-05-08|Followup|2011-05-29|2011-07-15|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|59.3||1|1|1|1|M|White||21|No|Mother|28270|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||31|28209|||Human Services: Non-Profit|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500910310|1|0|1|501600417|1|0|1|500363806|2||||4|3|||-2||-2|0|10|||7464|9|||1|169238||4|1|45
500771746|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2016-06-15|Followup|2011-05-29|2011-07-15|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Child: Graduated|84.6||3|4|1|2|F|Black||19||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||37|28012|Some College|Married|Finance: Banking|28208|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500772014|31|0|2|500996153|1|0|2|500366437|2||500004641||4|1|500004640||-2||-2|0|4|||7464|9|||1|169257||4|1|45
501741559|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-13|2011-10-13|Followup|2011-08-13|2011-09-07|Declined|Done||||||||3|3|3|4|3|3|3.17|||||||||3|3|3|3|2|3|2.83||||||4|4|4|4|||||||4|4|4|3|3.75||||||||||4|4|4|4|3|4|3|3.71||||||3|4|3|3.33|||||4|2|3||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|14||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||32|28208|Bachelors Degree|Married|Tech: Production Line||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501741899|31|0|1|502213067|31|0|1|500464036|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|169387|35898|4|1|45
501919692|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-13|2012-03-30|Followup|2011-08-13|2011-08-12|Complete|Done|4|3|4|3|3|4|3.5|3|3|3|3|3|4|3.17|10.41|3|4|4|4|4|4|3.83|4|1|1|2|4|4|2.67|43.45|4|4|4|4|4|4|4|4|0|4|5|5|4|4.5|5|3|3|4|3.75|20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|3|3|3|16.67|2|2|1|1|100|4|4||||Red||Volunteer: Lost contact with child/agency|19.5||1|1|1|1|M|White||16|No|Mother|28270|One Parent: Female|Unknown||No||Self|General Community||Enrollment|M|White||35|28270|Associate Degree|Married|Firefighter||1|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013709|501920088|1|0|1|502219683|1|0|1|500465111|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|169400|168273|4|3|45
502233621|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-14|2013-04-25|Followup|2011-08-10|2011-08-03|Complete|Done|3|2|3|1|3|3|2.5|3|4|4|4|3|4|3.67|-31.88|2|3|3|2|2|3|2.5|4|1|4|2|4|4|3.17|-21.14|4|4|3|3.67|4|4|4|4|-8.25|3|4|4|3|3.5|5|5|4|5|4.75|-26.32|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|4|4|4|-12.5|2|2|2|2|0||||||Green||Child/Family: Moved|32.4||1|1|2|2|M|Multi-race (Hispanic & White)||16|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction|28208|1|1|Igniting Breakfast|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500011746|502234052|35|0|1|502255664|1|0|1|500465113|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17266|8|||1|169561|168275|4|3|45
501811395|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-10|NaT|Followup|2011-03-10|2011-05-25|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Cabarrus County||84.2||1|1|1|1|F|Black||15|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||60|28213||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501811730|31|0|2|500876892|31|0|2|500436702|2||500016307||2|1|500016374|500016374|-2|500016374|-2|6854|8|||2238|7|||1|169985||4|0|45
502247430|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-17|2014-01-23|Followup|2011-08-17|2011-08-15|Declined|Done||||||||3|1|1|1|2|3|1.83|||||||||2|2|3|1|2|2|2||||||4|3|3|3.33|||||||2|3|2|4|2.75||||||||||4|4|4|4|4|4|3|3.86||||||2|4|4|3.33|||||2|1|1.5||||1|1|||||||Yellow||Child: Lost interest|41.2||1|1|1|1|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||63|28078|Bachelors Degree|Married|Medical: Nurse||10|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502247861|31|0|2|502226106|1|0|2|500465539|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|170099|166252|4|1|45
502193174|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-18|2011-12-28|Followup|2011-08-18|2011-08-10|Complete|Done|4|2|4|2|3|3|3|4|1|1|4|2|4|2.67|12.36|3|3|3|3|3|4|3.17|1|3|3|2|3|3|2.5|26.8|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|2|5|5|4|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|2|2|0|4|4||||Green||Volunteer: Lost contact with child/agency|16.3||2|2|1|1|M|Black||16||Mother|28273|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|Black||49|28277|Associate Degree|Married|Tech: Engineer||0|9|Recruitment Event|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|502193603|31|0|1|502187342|31|0|1|500465373|2||-2||4|1|||-2|500000294|-2|0|4|||7443|2|||1|170466|168695|4|3|45
501725168|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-31|2013-12-18|Followup|2011-08-31|2011-08-10|Complete|Early|3|1|1|1|2|3|1.83|||||||||1|3|3|2|2|4|2.5|||||||||4|4|4|4||||||2|5|5|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|2|2.67||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Moved|51.6||2|2|1|1|F|Multi-Race (None of the above)||15|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28269|Bachelors Degree|Married|Human Services: Non-Profit||2|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017777|501724831|7|0|2|501824761|1|0|2|500381463|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|170564||4|3|45
502260656|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-30|2010-09-22|Baseline|2010-08-19|2010-08-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|0.8||2|2|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28078|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||32|28025|Bachelors Degree|Single|Customer Service||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500002335|502261088|38|0|2|502031924|1|0|2|500466370|2||-2||4|1|||-2||-2|0|10|||46|2|||1|170947|-1|4|1|44
501731841|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-05|2013-08-30|Followup|2011-06-05|2011-06-30|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red|Amachi|Child: Lost interest|50.8||1|1|1|1|F|Black||18|Yes|Father|28210|One Parent: Male|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||49|28277|Bachelors Degree|Single|Business: Mgt, Admin||4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|501732181|31|0|2|501182066|31|0|2|500367022|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||46|2|||1|171130||4|3|45
502064627|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-20|NaT|Followup|2011-08-20|2011-08-11|Complete|Done|2|2|4|1|2|4|2.5|2|2|4|2|3|4|2.83|-11.66|2|3|4|3|2|4|3|3|3|4|3|2|4|3.17|-5.36|4|3|4|3.67|4|3|2|3|22.33|5|4|3|3|3.75|5|3|3|4|3.75|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|2|3|2.67|49.81|3|4|3.5|2|3|2.5|40|2|2|1|1|100|4|4||||Green|||78.9||1|1|2|2|M|Black||16|No|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|502065051|31|0|1|500773055|3|14|1|500462574|2||-2||2|1|||-2||-2|0|10|||46|2|||1|171135|159373|4|3|45
502114704|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-20|2012-01-10|Followup|2011-08-20|2011-11-04|Expired|Late||||||||1|4|2|1|3|3|2.33|||||||||4|4|2|4|4|4|3.67||||||4|4|4|4|||||||5|3|3|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|3|3.5||||1|1|||||||Green||Volunteer: Moved|16.7||1|1|1|1|F|Black||18|No|Mother|28270|One Parent: Female|Unknown||Yes|Radio|Media|General Community||RTBM|F|White||32|28204|Masters Degree|Single|Business: Marketing||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502115131|31|0|2|502130736|1|0|2|500460157|2||-2||4|1|||-2||-2|55|1|||7496|10|||1|171136|148929|4|0|45
501250109|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-11|2013-02-27|Followup|2011-09-11|2011-10-26|Comprehension|Done||||||||3|1|3|1|3|3|2.33|||||||||3|3|3|3|4|3|3.17||||||3|3|3|3|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Red||Volunteer: Lost contact with child/agency|41.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28227|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501250385|31|0|1|501790515|31|0|1|500381167|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|171164|13945|4|2|45
500186435|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-23|2015-08-20|Followup|2011-07-23|2011-08-22|Complete|Done|3|4|4|4|3|3|3.5|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|144.9||1|1|1|1|M|Black||20||Mother|28216|One Parent: Female|Unknown||No|Brochure|Media|General Community||Match Support|M|White||45|28226|Bachelors Degree|Married|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187988|31|0|1|500189358|1|0|1|500037395|2||-2||4|1|||-2||-2|51|1|||7496|10|||1|171222||4|3|45
501457406|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-20|2013-07-16|Followup|2011-08-20|2011-08-26|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|46.9||1|1|1|1|M|Black||21|No|Mother|28269|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28205|||Finance: Banking|28217|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|501457691|31|0|1|501720969|1|0|1|500375964|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|171242||4|3|45
501197292|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-06|2012-03-31|Followup|2011-06-06|2011-07-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|45.8||1|1|1|1|M|White||18|No|Mother|28110|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||50|28112|High School Graduate|Married|Business: Marketing|28105|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501197566|1|0|1|501240286|1|0|1|500269444|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|171361||4|1|45
500393176|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-07|2012-06-21|Followup|2011-06-07|2011-07-06|Complete|Done|3|3|3|2|3|3|2.83|||||||||2|3|2|2|2|2|2.17|||||||||4|3|3|3.33||||||3|3|3|2|2.75|||||||3|4|4|3|3|3|3|3.29||||||||||3|4|3|3.33||||||3|2|2.5|||||1|1|||||||||Green|Amachi|Child: Graduated|72.5||1|1|1|1|F|Black||22||Relative: Other|28216|Other Relative|Unknown||No||Relative|General Community|Amachi|Match Support|F|Black||35|28213||Single|Tech: Engineer||2|0|Bellafonte Presbyter|Faith Organization|Big|General Site|Amachi|Enrollment|277|60|598|500000170|500013781|500187361|31|0|2|500415570|31|0|2|500101074|2||500003586||4|1|500000294|500000294|-2|500000294|-1|0|3|||2238|7|||1|171460||4|3|45
502268597|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-01|2011-10-25|Baseline|2010-08-23|2010-09-01|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|1|3|4|3.17|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1|||||||||Green||Child/Family: Moved|13.8||1|1|1|1|F|Black||16|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||37|28211|Bachelors Degree|Single|Arts, Entertainment, Sports||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|502269029|31|0|2|502097001|1|0|2|500466598|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|171619|-1|4|3|44
502259491|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-25|2012-10-15|Baseline|2010-08-24|2010-08-25|Complete|Done|1|2|1|1|1|1|1.17|||||||||2|1|1|2|3|||||||||||3|2|2|2.33||||||2|2|2|2|2|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Green||Child: Lost interest|25.7||1|1|4|5|F|White||20|No|Mother|28027|Two Parent|Unknown|Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|277|60|598|500000170|500002335|502259924|1|0|2|501306527|1|0|2|500466849|2||-2||4|1|||-2|500014681, 500016374|-2|0|5|||7464|9|||1|172003|-1|4|3|44
502168082|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-05|2012-01-26|Baseline|2010-08-24|2011-01-05|Complete|Done|3|1|1|1|3|2|1.83|||||||||3|4|3|4|3|3|3.33|||||||||4|4|3|3.67||||||4|4|3|2|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2|||||||||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|12.7||1|1|1|1|F|Black||16|No|GrandMother|28208|Grandparents|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|White||43|28210|Bachelors Degree|Single|Business: Sales|6830|3|0|Self|Self|Big|General Community||RTBM|277|60|598|500000170|500013709|502168511|31|0|2|502240884|1|0|2|500505682|2||-2||4|3|500005291|500005291|-2||-2|34|2|||7464|9|||1|172086|-1|4|3|44
500474486|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-23|2015-08-18|Followup|2011-08-23|2011-08-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|107.8||1|1|1|1|M|Black||20||Mother|28214|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||38|28209|Bachelors Degree|Single|Construction|28247|0|2|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500474735|31|0|1|500491064|31|0|1|500118168|2||-2||4|3|||-2||-2|34|2|||7447|3|||1|172482||4|1|45
502259491|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-25|2012-10-15|Followup|2011-08-25|2011-11-09|Expired|Late||||||||1|2|1|1|1|1|1.17|||||||||2|1|1|2|3||||||||3|2|2|2.33|||||||2|2|2|2|2||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||1|1|||||||Green||Child: Lost interest|25.7||1|1|4|5|F|White||20|No|Mother|28027|Two Parent|Unknown|Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|277|60|598|500000170|500002335|502259924|1|0|2|501306527|1|0|2|500466849|2||-2||4|1|||-2|500014681, 500016374|-2|0|5|||7464|9|||1|172592|172003|4|0|45
500761491|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2013-03-22|Followup|2011-08-27|2011-08-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|30.8||3|3|1|1|F|Black||16||Aunt|28213|One Parent: Female|$40,000 to $44,999|Y|No||Self|General Community||Enrollment|F|Black||61|28269|Bachelors Degree|Divorced|Education: Teacher|28215|1|1|LPL Financial|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500761759|31|0|2|502189613|31|0|2|500465204|2||-2||4|1|||-2||-2|0|10|||11247|3|||1|173198||4|1|45
502173588|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2012-08-30|Followup|2011-07-28|2011-07-28|Complete|Done|3|3|3|2|3|2|2.67|3|1|2|1|3|3|2.17|23.04|3|4|4|3|3|4|3.5|2|3|3|2|2|3|2.5|40|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|4|3|3.5|14.29|4|4|4|4|4|4|4|4|2|2|2|1|1|2|1|1.57|154.78|4|4|4|4|4|4|4|4|0|4|4|4|2|1|1.5|166.67|2|2|1|1|100||||||Yellow|Amachi|Volunteer: Lost contact with child/agency|24.1||2|2|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||No|A Child's Place|Service Organization|General Community|Amachi|Enrollment|F|White||29|28217|Bachelors Degree|Single|Customer Service||5|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502174017|31|0|2|502085998|1|0|2|500463449|2||500003586||4|2|500000294|500000294|-2||-2|7016|11|||7496|10|||1|173252|160541|4|3|45
502253085|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-13|2011-10-25|Baseline|2010-08-27|2010-09-13|Complete|Done|3|3|4|3|3|3|3.17|||||||||3|3|4|2|2|4|3|||||||||4|3|4|3.67||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Moved|13.4||1|1|3|3|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||RTBM|M|Black||45|28262|Bachelors Degree|Married|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500011184|502253517|31|0|1|502087592|31|0|1|500467804|2||-2||4|1|||-2|500014505, 500015184|-1|6854|8|||7462|13|||1|173279|-1|4|3|44
502262725|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-30|2011-04-21|Baseline|2010-08-27|2010-08-30|Complete|Done|1|1|1|1|1|1|1|||||||||3|1|4|2|4|3|2.83|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1|||||||||Yellow||Child/Family: Lost contact with volunteer/agency|7.7||1|1|2|2|F|Black||16|No|Mother|28217|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||29|28277|Bachelors Degree|Single|Consultant|28204|0|11|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011639|502263157|31|0|2|502231024|1|0|2|500467811|2||-2||4|2|||-2|500000294|-2|6854|8|||46|2|||1|173285|-1|4|3|44
501332658|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-01-19|Followup|2010-09-29|2010-10-04|Complete|Done|3|3|2|2|3|3|2.67|||||||||3|4|3|2|2|3|2.83|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2|||||||||Green|Amachi|Child: Severity of challenges|87.7||1|1|1|1|M|Black||15|Yes|GrandMother|28213|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||46|28227|High School Graduate|Single|Medical: Healthcare Worker|28269|4|0|Coworker|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500020752|501332937|31|0|1|501814288|1|0|1|500384166|2||-2||4|1|500000294|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||7447|3|||1|173373||4|3|45
501810015|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-19|2012-02-09|Followup|2010-10-19|2010-10-20|Complete|Done|2|2|4|2|4|4|3|||||||||4|4|4|3|4|3|3.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|1|2.67||||||4|4|4|||||2|2|||||||||Green||Child/Family: Unrealistic expectations|27.7||1|1|2|2|M|Hispanic||15|No|Mother|28210|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501810370|3|0|1|501646021|3|0|1|500391598|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|173608||4|3|45
500399525|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-15|2012-08-29|Followup|2011-06-15|2011-08-02|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Agency: Challenges with program/partnership|74.5||1|1|1|1|F|Black||19||Mother|28214|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||46|28217|Some College|Single|Finance: Accountant|28208|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500399775|31|0|2|500416787|31|0|2|500099891|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|173623||4|1|45
502062624|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-30|2012-12-19|Followup|2011-08-30|2011-09-15|Complete|Done|3|3|4|2|2|2|2.67|3|3|3|2|1|4|2.67|0|2|4|3|3|4|3|3.17|2|4|3|3|3|4|3.17|0|4|4|4|4|4|4|4|4|0|3|5|4|5|4.25|3|5|3|5|4|6.25|4|4|4|4|4|3|3|3.71|4|4|4|4|4|4|4|4|-7.25|3|4|4|3.67|4|4|4|4|-8.25|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4||||Yellow||Volunteer: Feels incompatible with child/family|27.7||1|1|1|1|F|Black||16|No|Mother|28081|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||32|28083|Bachelors Degree|Single|Tech: Computer/Programmer|28216|1|7|LPL Financial|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|502063048|31|0|2|502067861|31|0|2|500460279|2||-2||4|2|||-2||-2|0|10|||11247|3|||1|173809|155833|4|3|45
502249063|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-17|2011-01-31|Baseline|2010-08-30|2010-09-16|Complete|Done|3|3|3|4|2|3|3|||||||||3|4|4|3|3|4|3.5|||||||||3|3|3|3||||||4|5|3|5|4.25|||||||4|4|4|4|3|3|2|3.43||||||||||3|4|4|3.67||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Time constraint|4.5||1|1|1|1|M|White||19|No|Mother|28277|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||49|28277|Bachelors Degree|Married|Self-Employed, Entrepreneur|28277|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500010355|502249494|1|0|1|502266549|1|0|1|500468039|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|173810|-1|4|3|44
501157075|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-30|2012-05-23|Followup|2011-08-30|2011-10-10|Complete|Done|3|4|4|3|2|4|3.33|||||||||2|3|3|3|2|3|2.67|||||||||4|4|4|4||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Red|Amachi|Volunteer: Lost contact with child/agency|20.8||3|4|2|2|F|Black||17||Relative: Other|28206|Grandparents|Unknown||Yes||School|General Community|Amachi|Match Support|F|Black||34|28216|Masters Degree|Single|Business|28202|8|7|Self|Self|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|277|60|598|500000170|500008629|501157349|31|0|2|502261758|31|0|2|500467512|2||500003586||4|3|500000294|500000294|-2|500014505, 500014506|-1|0|4|||7464|9|||1|173939||4|3|45
500970267|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-29|NaT|Baseline|2010-08-31|2010-09-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||77.5||1|1|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||61|28204||Divorced|Self-Employed, Entrepreneur||0|0|Billboard|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|2|502084649|1|0|2|500468192|2||500003586||2|1|500000294|500000294|-2|500000294|-2|5635|9|||125|1|||1|174196|-1|4|1|44
501749652|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-01|2013-11-07|Followup|2012-09-01|2012-08-29|Complete|Done|3|2|4|1|4|4|3|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Child/Family: Moved|38.2||1|1|2|2|M|Black||18||Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|Black||52|28107|Some College|Divorced|Tech: Engineer|28262|3|0|Local Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500012459|501749994|31|0|1|501645507|31|0|1|500464305|2||-2||4|2|||-2||-2|0|10|||7437|1|||1|174657|38597|4|3|45
501776333|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-08|2013-07-25|Followup|2011-09-08|2011-08-31|Complete|Done|3|2|1|1|3|3|2.17|3|2|3|2|4|4|3|-27.67|4|4|4|3|4|4|3.83|3|3|3|2|3|3|2.83|35.34|4|4|4|4|3|3|3|3|33.33|4|4|5|4|4.25|4|4|4|4|4|6.25|3|4|4|4|4|4|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|4|4|4|4|-8.25|4|2|3|3|3|3|0|1|1|2|2|-50|4|4||||Green||Volunteer: Moved|46.5||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28210|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|501776688|31|0|1|501832599|31|0|1|500381636|2||-2||4|1|||-2|500000294|-2|34|2|||7464|9|||1|174982|9814|4|3|45
500483980|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-01|2014-03-24|Followup|2011-09-01|2011-09-30|Complete|Done|3|3|3|3|4|4|3.33|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|90.7||1|1|2|2|M|Black||21||Mother|28227|One Parent: Female|$10,000 to $14,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||71|28270||Single|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500484231|31|0|1|500423426|31|0|1|500120592|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|175008||4|3|45
500186765|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-05|2013-08-15|Followup|2011-09-05|2011-11-02|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|107.3||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||46|28078|Masters Degree|Widowed|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500004169|500188083|31|0|2|500189359|31|0|2|500037396|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|175296||4|1|45
500722500|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-20|2011-10-26|Followup|2011-06-20|2011-09-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|52.2||2|2|1|1|F|White||20||Mother|28027||Unknown||No||Service Organization|General Community||Match Support|F|White||34|28083|Bachelors Degree|Single|Education: Teacher Asst/Aid|28147|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|500722767|1|0|2|500830633|1|0|2|500180184|2||-2||4|1|||-2||-2|0|11|||7464|9|||1|175396||4|0|45
500186946|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-20|2012-08-23|Followup|2011-06-20|2011-07-06|Complete|Done|3|2|3|3|3|3|2.83|||||||||2|2|2|1|2|2|1.83|||||||||4|3|2|3||||||3|3|3|3|3|||||||4|4|4|3|3|3|2|3.29||||||||||3|4|3|3.33||||||2|2|2|||||2|2|||||||||Red|Amachi|Volunteer: Lost contact with child/agency|62.1||2|2|1|1|F|Black||19|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||36|28262||Single|Education: Teacher||4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188139|31|0|2|500865596|31|0|2|500181565|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|175399||4|3|45
501257717|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-20|2012-10-30|Followup|2011-06-20|2011-06-30|Complete|Done|4|1|4|1|1|1|2|||||||||4|4|1|1|4|4|3|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||1|4|4|3||||||2|2|2|||||2|2|||||||||Green||Volunteer: Time constraint|52.3||2|2|2|2|F|Black||17|No|GrandMother|28203|Grandparents|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|White||31|28204|Bachelors Degree|Single|Finance: Banking||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|501257994|31|0|2|500839705|1|0|2|500271936|2||-2||4|1|||-2||-2|0|10|||46|2|||1|175421||4|3|45
500383915|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-20|2012-08-30|Followup|2011-06-20|2011-08-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|50.3||2|2|2|2|F|Black||20||GrandMother|28205|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||64|28269||Married|Finance: Economist||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|500384165|31|0|2|500540512|31|0|2|500274279|2||-2||4|1|||-2||-2|6855|8|||7464|9|||1|175425||4|1|45
500186956|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-21|2015-03-04|Followup|2011-06-21|2011-07-06|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|128.4||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28203|Bachelors Degree|Married|Law: Lawyer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|500189727|1|0|1|500037841|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|175500||4|1|45
501721760|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-22|2016-11-01|Followup|2011-06-22|2011-07-15|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|2|3|1|1|3|2|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Volunteer: Infraction of match rules/agency policies|88.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||59|28269|Masters Degree|Married|Clergy||0|0|Coca Cola|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|501722098|31|0|1|501755476|1|0|1|500368545|2||-2||4|1|||-2|500000294|-2|0|10|||9610|3|||1|175627||4|3|45
501212662|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-23|2013-04-22|Followup|2011-06-23|2011-06-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|58||1|1|1|1|M|Multi-Race (None of the above)||16|Yes|Mother|28211|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Multi-Race (None of the above)||34|28205|Bachelors Degree|Single|Business: Sales|28210|0|10|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501212937|7|0|1|501252394|7|0|1|500269647|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|175707||4|1|45
501234601|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-24|2012-08-29|Followup|2011-06-24|2011-08-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|50.2||1|1|2|2|F|Black||23|No|Mother|28215|Grandparents|Unknown||No|TV|Media|General Community||Match Support|F|Black||48|28211|Bachelors Degree|Single|Consultant|28278|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500008629|501234877|31|0|2|501223094|31|0|2|500271822|2||-2||4|2|||-2|500014505, 500015184|-1|56|1|||7462|13|||1|176034||4|1|45
502245018|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-21|2011-02-16|Baseline|2010-09-10|2010-09-21|Complete|Done|3|4|4|4|3|3|3.5|||||||||2|3|2|3|3|2|2.5|||||||||4|3|3|3.33||||||2|3|4|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2|||||||||Green||Volunteer: Moved|4.9||1|1|3|3|M|Hispanic||20|No|Mother|28217|One Parent: Female|Unknown||No|Radio|Media|General Community||Match Support|M|White||36|28202|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500010765|502245449|3|0|1|501811850|1|0|1|500469733|2||-2||4|1|||-2||-2|55|1|||7464|9|||1|176909|-1|4|3|44
500402676|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-27|2012-02-29|Followup|2011-06-27|2011-06-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Graduated|68.1||1|1|1|1|M|White||24|||28211|One Parent: Female|Unknown||No||Therapist/Counselor|General Community|Amachi|Match Support|M|White||36|28208|Bachelors Degree|Single|Business: Mgt, Admin|28203|2|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500402926|1|0|1|500339569|1|0|1|500102368|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|5|||2238|7|||1|177190||4|1|45
500186374|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-28|2012-01-10|Followup|2011-06-28|2011-08-12|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|66.4||2|2|1|1|F|Black||22||Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||55|28269|High School Graduate|Single|Business: Human Resources|28202|5|0|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008629|500187968|31|0|2|500419439|31|0|2|500102160|2||-2||4|2|||-2||-2|0|10|||6247|12|||1|177333||4|1|45
500402978|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-29|2012-05-08|Followup|2011-06-29|2011-06-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Time constraints|70.3||1|1|1|1|M|White||22||Mother|28211|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||33|28203|Bachelors Degree|Single|Business: Sales|27609|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500402926|1|0|1|500414710|1|0|1|500103314|2||-2||4|2|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|177432||4|1|45
502211307|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-03|2014-04-24|Baseline|2010-09-13|2011-02-03|Complete|Done|4|4|4|3|4|3|3.67|||||||||4|3|3|4|3|3|3.33|||||||||4|4|4|4||||||4|4|4|||||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4|||||||3||||||2|2|||||||||Yellow|Amachi|Volunteer: Time constraint|38.6||1|1|1|1|M|Black||16|Yes|Mother|28278|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||51|28214|Bachelors Degree|Single|Business: Sales|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502211737|31|0|1|502371462|1|0|1|500512414|2||-2||4|2|500000294|500000294|-2|500000294|-2|7016|11|||7496|10|||1|177660|-1|4|3|44
502265907|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-31|2012-02-22|Baseline|2010-09-13|2011-01-31|Complete|Done|4|4|4|4|3|4|3.83|||||||||2|2|3|4|2|4|2.83|||||||||4|4|4|4||||||3|5|3|4|3.75|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|4|4||||||4|4|4|||||1|1|||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|12.7||1|1|1|1|F|Black||19|Yes|Mother|28210|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||37|28209|PHD|Single|Medical: Doctor, Provider|28210|2|3|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502266339|31|0|2|501332017|1|0|2|500512367|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|177670|-1|4|3|44
500539341|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-24|2012-01-27|Followup|2011-09-24|2011-09-19|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|3|3|3|2.83|||||||||4|3|3|3.33||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Child: Family structure changed|64.1||1|1|2|2|M|White||19|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||44|28205||Single|Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|500539592|1|0|1|500191356|1|0|1|500123020|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|178178||4|3|45
501101149|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-01|NaT|Followup|2011-07-01|2011-07-16|Complete|Done|3|4|4|4|1|2|3|||||||||2|1|4|4|2|4|2.83|||||||||4|4|4|4||||||4|4|5|3|4|||||||4|4|4|4|4|4|4|4||||||||||3|1|1|1.67||||||4|4|4|||||2|2|||||||||Yellow|||104.5||1|2|1|2|F|White||16||Mother|28270|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||55|28277|Masters Degree|Widowed|Consultant||5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|501101423|1|0|2|500834694|1|0|2|500276073|2||-2||2|2|||-2||-2|0|4|||7671|13|||1|178305||4|3|45
502264006|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-22|2017-02-26|Baseline|2010-09-16|2010-09-22|Complete|Done|2|1|3|1|2|3|2|||||||||1|3|2|2|1|3|2|||||||||4|4|4|4||||||4|2|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|3|3.5|||||1|1|||||||||Red||Child: Lost interest|77.2||1|1|1|1|F|Hispanic||16|No|Mother|28211|One Parent: Female|Unknown||Yes|Spanish Print|Media|General Community||Match Support|F|Hispanic||38|28202|Bachelors Degree|Single|Tech: Engineer|28202|12|0|Big Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020753|502264438|3|0|2|502274748|3|0|2|500470897|2||-2||4|3|||-2||-2|7063|1|||7456|8|||1|178842|-1|4|3|44
500187075|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-21|2014-01-16|Followup|2011-09-21|2011-09-19|Complete|Done|3|3|3|3|3|3|3|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||2|3|3|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|111.8||1|1|6|6|F|Black||21||Mother|28205|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||38|28209|Bachelors Degree|Single|Human Services: Non-Profit||0|0|Recruitment Event|Self|Big|General Site||Match Support|277|60|598|500000170|500012459|500188223|31|0|2|500189550|1|0|2|500037643|2||-2||4|1|||-2||-1|0|10|||7458|9|||1|178914||4|3|45
500896018|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-03|2014-08-14|Followup|2011-07-03|2011-09-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|73.4||1|1|1|1|F|Black||20|Yes|Mother|28027|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||40|28027|Bachelors Degree|Separated|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500896288|31|0|2|501225232|31|0|2|500269506|2||-2||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|179197||4|0|45
501750505|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-31|2012-06-28|Followup|2011-07-31|2011-09-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|34.9||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|Black||32|28205|Bachelors Degree|Single|Finance: Banking||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501750847|31|0|1|501777375|31|0|1|500375403|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|179613||4|1|45
502290880|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-20|2014-03-31|Baseline|2010-09-20|2010-10-20|Complete|Done|4|3|3|1|4|4|3.17|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2|||||||||Green|Project Big|Child/Family: Time constraints|41.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|M|White||35|28202|Bachelors Degree|Single|Real Estate: Realtor|28208|2|10|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502291312|31|0|1|502261364|1|0|1|500471473|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7496|10|||1|179708|-1|4|3|44
501234604|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-23|2012-09-06|Followup|2011-07-23|2011-09-06|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Severity of challenges|49.5||1|1|1|1|F|Black||19|No|Mother|28215|Grandparents|Unknown||No||Self|General Community||Match Support|F|Black||38|28213|Masters Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008629|501234880|31|0|2|501165150|31|0|2|500278984|2||-2||4|2|||-2||-2|0|10|||46|2|||1|180204||4|1|45
500186277|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2014-07-16|Followup|2011-07-08|2011-07-07|Complete|Done|4|1|1|1|2|3|2|||||||||2|4|4|4|1|4|3.17|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2|||||||||Red||Child/Family: Moved|60.3||3|4|2|3|F|Black||18||Mother|28206|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||39|28210|Bachelors Degree|Married|Business: Sales||8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500187876|31|0|2|500188587|1|0|2|500373187|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|180205||4|3|45
501791428|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-29|2012-09-06|Followup|2011-07-29|2011-09-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|37.3||1|1|1|1|M|Black||19|No|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Multi-Race (None of the above)||33|28273|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501163776|31|0|1|501726049|7|0|1|500374912|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|180206||4|1|45
500185647|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-09|2013-10-31|Followup|2011-07-09|2011-07-19|Complete|Done|3|2|4|3|4|4|3.33|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2|||||||||Green|Amachi|Child: Graduated|123.8||1|2|1|2|F|Black||21|Yes|Mother|28217|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||38|28269|Bachelors Degree|Married|Unknown|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187284|31|0|2|500188649|31|0|2|500038124|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|180208||4|3|45
501240369|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-10-09|Followup|2011-07-10|2011-08-09|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|75||1|1|1|1|M|Black||20|Yes|Mother|28214|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||43|28269|Masters Degree|Single|Business: Mgt, Admin|28202|3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501240645|31|0|1|501240602|1|0|1|500272039|2||500003586||4|1|500000294|500000294|-2||-2|0|3|||131|1|||1|180210||4|1|45
500186682|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2015-07-22|Followup|2011-07-20|2011-08-09|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|96.1||3|4|1|1|M|Black||20|Yes|Mother|28227|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|M|Black||57|28262||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|500887363|31|0|1|500184396|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|180211||4|1|45
500186960|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-31|2013-08-15|Followup|2011-07-31|2011-08-09|Complete|Done|3|3|3|3|3|4|3.17|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||3|4|4|4|3|3|3|3.43||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|72.5||2|2|1|1|M|White||19|Yes|Mother|28227|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||40|28105|Some College|Married|Military|28112|11|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188147|1|0|1|500738970|1|0|1|500186719|2||500003586||4|3|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|180212||4|3|45
500417281|BBBS of Greater Charlotte|Main Office|C|Completed|2006-07-31|2013-01-31|Followup|2011-07-31|2011-08-09|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|78.1|Y|1|1|1|1|F|White||16||Mother|28211|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||48|28211|Masters Degree|Married|Finance: Banking|28202|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500402926|1|0|2|500349297|1|0|1|500112798|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|180213||4|3|45
501078559|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-04|2012-06-21|Followup|2011-08-04|2011-08-09|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|46.6||1|1|1|1|M|Black||22|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||37|28269|Bachelors Degree|Single|Medical: Admin|19380|0|9||Relative|Big|General Community||Match Support|277|60|598|500000170|500013781|501078832|31|0|1|501262050|1|0|1|500279449|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||0|11|||1|180214||4|3|45
501347097|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-30|2014-10-16|Followup|2011-07-30|2011-07-18|Complete|Done|3|4|4|4|3|4|3.67|||||||||1|3|2|4|2|3|2.5|||||||||3|4|4|3.67||||||3|4|2|2|2.75|||||||4|3|4|4|3|4|4|3.71||||||||||3|4|4|3.67||||||4|4|4|||||2|2|||||||||Yellow||Volunteer: Time constraint|74.5||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||35|28078|Bachelors Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501347376|31|0|2|501099568|1|0|2|500278256|2||-2||4|2|||-2||-2|0|10|||46|2|||1|180335||4|3|45
501641337|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-07|2015-03-13|Followup|2011-08-07|2011-08-04|Complete|Done|4|4|4|2|4|3|3.5|||||||||3|4|4|4|3|4|3.67|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|3|4|3|3|3|3.43||||||||||3|4|3|3.33||||||3|2|2.5|||||1|1|||||||||Green||Volunteer: Moved|67.2||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||31|28269|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|2|500835981|31|0|2|500373972|2||-2||4|1||500000294|-2|500000294|-2|0|10|||46|2|||1|180346||4|3|45
502264006|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-22|2017-02-26|Followup|2011-09-22|2011-10-02|Complete|Done|4|3|3|3|3|4|3.33|2|1|3|1|2|3|2|66.5|3|4|4|4|3|4|3.67|1|3|2|2|1|3|2|83.5|4|4|4|4|4|4|4|4|0|4|||3||4|2|3|4|3.25||4|4|4|4||4|4||4|4|4|4|4|4|4|4||4|4|4|4|3|4|3|3.33|20.12|4|4|4|4|3|3.5|14.29|1|1|1|1|0|4|4||||Red||Child: Lost interest|77.2||1|1|1|1|F|Hispanic||16|No|Mother|28211|One Parent: Female|Unknown||Yes|Spanish Print|Media|General Community||Match Support|F|Hispanic||38|28202|Bachelors Degree|Single|Tech: Engineer|28202|12|0|Big Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020753|502264438|3|0|2|502274748|3|0|2|500470897|2||-2||4|3|||-2||-2|7063|1|||7456|8|||1|180643|178842|4|3|45
502269033|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-29|2011-03-29|Baseline|2010-09-22|2010-09-29|Complete|Done|4|4|4|2|3|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|Amachi, Project Big, Project Big AND Amachi|Child/Family: Unrealistic expectations|5.9||1|1|2|2|F|Multi-race (Black & White)||17|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Relative|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community|Project Big AND Amachi|Match Support|277|60|598|500000170|500011184|502265485|36|0|2|502208867|31|0|2|500472485|2||500004772||4|1|500000294, 500004640, 500004901|500004640, 500004901|-2|500004901|-2|0|3|||7464|9|||1|180839|-1|4|3|44
502248736|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-11|2011-02-08|Baseline|2010-09-22|2010-10-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Health|3.9||1|1|1|1|M|Black||16|No|Mother|28027|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|Black||61|28027||Single|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|502249167|31|0|1|502266779|31|0|1|500472618|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|180971|-1|4|1|44
502230729|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-09|2012-08-27|Baseline|2010-09-23|2011-03-09|Complete|Done|4|2|3|2|3|4|3|||||||||2|4|3|3|3|3|3|||||||||3|3|2|2.67||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Moved|17.6||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||36|28277|Bachelors Degree|Single|Student: College|28205|0|4|Recruitment Event|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|277|60|598|500000170|500012459|502231160|1|0|1|502483362|1|0|1|500518850|2||-2||4|2|500005291|500005291|-2|500000294, 500005291|-2|34|2|||7459|10|||1|181484|-1|4|3|44
500970267|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-29|NaT|Followup|2011-09-29|2011-10-25|Complete|Done|4|4|4|1|4|4|3.5|||||||||1|3|3|2|4|3|2.67|||||||||4|4|4|4||||||2|4|2|5|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green|Amachi||77.5||1|1|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||61|28204||Divorced|Self-Employed, Entrepreneur||0|0|Billboard|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|2|502084649|1|0|2|500468192|2||500003586||2|1|500000294|500000294|-2|500000294|-2|5635|9|||125|1|||1|183843|174196|4|3|45
502172536|BBBS of Greater Charlotte|Main Office|C|Active|2010-10-13|NaT|Baseline|2010-09-30|2010-10-13|Complete|Done|3|2|4|3|1|1|2.33|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|2|3|||||2|2|||||||||Green|||77.1||1|1|1|1|F|Black||17|No|Mother|28269|Two Parent|Unknown||Yes||Relative|General Community||Match Support|F|Multi-race (Asian & White)||33|28205|Masters Degree|Married|Finance: Economist|28223|7|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502172965|31|0|2|501279665|37|0|2|500475431|2||-2||2|1|||-2||-2|0|3|||129|1|||1|184611|-1|4|3|44
501627668|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2012-09-14|Followup|2011-01-26|2011-01-04|Complete|Early|3|2|3|3|3|3|2.83|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Moved|31.6||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||38|28209|Bachelors Degree|Single|Business|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|501627988|31|0|1|501865457|1|0|1|500423715|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|185079||4|3|45
501641325|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-24|2015-08-03|Followup|2011-06-24|2011-08-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|73.3||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Multi-race (Asian & White)||34|28205|Bachelors Degree|Single|Tech: Research/Design|28255|3|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|1|501715652|37|0|1|500366872|2||-2||4|1||500000294|-2|500000294|-2|6854|8|||7464|9|||1|185082||4|1|45
500728622|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-16|2012-05-23|Followup|2011-08-16|2011-10-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|57.2||1|2|1|2|M|Black||18|No|Mother|28205|One Parent: Female|Unknown||No||School|General Site||Match Support|M|Black||78|28216||Married|Retired||20|0|Other|BBBS Board/Staff|Big|General Site||Match Support|277|60|598|500000170|500008629|500730811|31|0|1|500546003|31|0|1|500188249|2||-2||4|2|||-1||-1|0|4|||7671|13|||1|185242||4|1|45
500186665|BBBS of Greater Charlotte|Main Office|C|Completed|2004-07-20|2013-02-28|Followup|2011-07-20|2011-09-13|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|103.3||1|1|1|1|M|Black||21||Mother|28202|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|Black||40|28207||Single|Medical: Nurse||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500188050|31|0|1|500189566|31|0|1|500037664|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|185916||4|1|45
500948385|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-28|2013-01-09|Followup|2011-08-28|2011-10-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|64.4||1|1|1|1|F|Black||17|No|Mother|28214|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Asian|Chinese|32|28216|||Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|500948655|31|0|2|500885771|4|16|2|500187434|2||-2||4|2|||-2||-2|34|2|||46|2|||1|186212||4|1|45
501300101|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-14|2015-05-11|Followup|2011-08-14|2011-08-15|Complete|Done|4|2|4|3|3|3|3.17|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|2|3|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2|||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|80.9||1|1|4|4|F|Black||19|Yes|GrandMother|28273|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501300379|31|0|2|500346193|31|0|2|500281421|2||500003586||4|2|500000294|500000294|-2||-2|7294|13|||46|2|||1|186213||4|3|45
500465521|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-21|2012-05-31|Followup|2011-08-21|2011-08-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|69.3||1|1|1|1|F|Black||23|Yes|Mother|28262|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|F|White||42|28209|Masters Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|2|500542558|1|0|2|500118432|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|186217||4|1|45
500465511|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-21|2013-10-31|Followup|2011-08-21|2011-08-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Graduated|86.3||1|1|1|1|M|Black||21|Yes|Mother|28262|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|M|White||54|28210|Masters Degree|Married|Finance: Accountant||0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500527675|1|0|1|500118120|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|4|||2230|7|||1|186218||4|1|45
500465506|BBBS of Greater Charlotte|Main Office|C|Active|2006-08-21|NaT|Followup|2011-08-21|2011-08-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi||126.8||1|1|1|1|M|Black||16|Yes|Mother|28262|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||54|28226|Bachelors Degree|Married|Arts, Entertainment, Sports||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500496966|1|0|1|500118121|2||500003586||2|2|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|186219||4|1|45
500186675|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-23|2013-08-29|Followup|2011-08-23|2011-09-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|72.2||4|4|1|1|F|Black||20|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||38|28221||Single|Human Services: Youth Worker||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188055|31|0|2|500865601|31|0|2|500185332|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|186220||4|1|45
500186938|BBBS of Greater Charlotte|Main Office|C|Completed|2004-08-24|2011-12-21|Followup|2011-08-24|2011-09-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Lost contact with child/agency|87.9||1|1|1|1|F|Black||21||Mother|28215|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||40|28217|Bachelors Degree|Single|Finance: Accountant|28277|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188131|31|0|2|500189708|31|0|2|500037821|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|186221||4|1|45
501825910|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-24|2016-09-23|Followup|2011-08-24|2011-09-07|Complete|Done|3|3|4|3|4|4|3.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|85||1|1|1|1|M|Black||16|Yes|Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|White||51|28214|Masters Degree|Married|Business: Sales|94108|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|501196986|1|0|1|500380446|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||7496|10|||1|186222||4|3|45
501332658|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-01-19|Followup|2011-09-29|2011-10-10|Complete|Done|3|3|2|3|3|2|2.67|||||||||1|4|4|4|4|4|3.5|||||||||3|2|4|3||||||5|5|5|5|5|||||||3|4|4|4|4|4|4|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Severity of challenges|87.7||1|1|1|1|M|Black||15|Yes|GrandMother|28213|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||46|28227|High School Graduate|Single|Medical: Healthcare Worker|28269|4|0|Coworker|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500020752|501332937|31|0|1|501814288|1|0|1|500384166|2||-2||4|1|500000294|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||7447|3|||1|186225||4|3|45
501645192|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-21|2016-08-19|Followup|2011-07-21|2011-10-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|85||1|1|2|2|M|Hispanic||19|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501645515|3|0|1|501519306|1|0|1|500374818|2||-2||4|3||500016374|-2|500016374|-2|0|10|||7464|9|||1|186437||4|0|45
500267459|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-19|2013-02-27|Followup|2011-09-19|2011-09-20|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|77.3||1|1|1|1|M|Black||16||Mother|28203|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28202|Bachelors Degree|Single|Finance: Accountant||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|500187395|31|0|1|500464544|1|0|1|500121193|2||-2||4|3|||-2||-2|0|10|||46|2|||1|186502||4|1|45
501597228|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-04|NaT|Followup|2011-09-04|2011-09-07|Complete|Done|3|3|3|3|3|3|3|||||||||2|2|2|4|3|3|2.67|||||||||4|3|1|2.67||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi||90.3||1|1|1|1|F|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||40|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28204|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501597548|31|0|2|501397328|31|0|2|500379964|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|186505||4|3|45
502278018|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-25|2011-03-30|Baseline|2010-10-07|2010-10-25|Complete|Done|3|4|4|4|2|3|3.33|||||||||4|4|3|4|4|3|3.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|2|3|3|3.43||||||||||3|4|1|2.67||||||4|1|2.5|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|5.1||2|2|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||26|28215|High School Graduate|Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|502278450|31|0|1|502227238|1|0|1|500477903|2||-2||4|2|||-2||-2|0|10|||46|2|||1|187800|-1|4|3|44
501811375|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-27|2013-08-28|Followup|2011-07-27|2011-10-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|49.1||1|1|3|3|F|Black||21|No|Mother|28027|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||41|28027|PHD|Single|Medical: Doctor, Provider|28075|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|501811730|31|0|2|501391123|31|0|2|500374230|2||-2||4|2|||-2|500016374|-2|0|8|||7464|9|||1|188871||4|0|45
500970264|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2013-06-17|Baseline|2010-10-11|2010-10-27|Complete|Done|4|3|3|2|3|3|3|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4||||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red|Amachi|Volunteer: Lost contact with child/agency|31.7||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Enrollment|M|Black||44|28269|Some High School|Single|Insurance||0|2|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|1|502250629|31|0|1|500478922|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||12183|14|1209|1|1|189150|-1|4|3|44
502063945|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-21|2016-08-05|Baseline|2010-10-11|2010-10-21|Complete|Done|3|3|3|2|2|3|2.67|||||||||2|3|3|1|3|2|2.33|||||||||3|2|2|2.33||||||3|2|4|2|2.75|||||||4|4|4|4|4|3|2|3.57||||||||||3|4|3|3.33||||||1|4|2.5|||||2|2|||||||||Yellow||Volunteer: Time constraint|69.5||1|1|1|1|M|White||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community||Match Support|M|White||37|28205||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502064367|1|0|1|502295138|1|0|1|500478943|2||500004641||4|2|||-2||-2|0|5|||7496|10|||1|189168|-1|4|3|44
502063943|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-20|2012-10-31|Baseline|2010-10-11|2012-06-19|Complete|Done|4|4|4|3|3|4|3.67|||||||||2|4|4|3|2|3|3|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||1|1||||4|4||||Red||Child: Severity of challenges|4.4||1|1|1|1|M|White||19|No|Mother|28213|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community||Match Support|M|White||62|28209|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502064367|1|0|1|502890782|1|0|1|500617038|2||-2||4|3|||-2||-2|0|5|||7439|1|1209|1|1|189170|-1|4|3|44
500186174|BBBS of Greater Charlotte|Main Office|C|Completed|2005-07-28|2012-10-31|Followup|2011-07-28|2011-08-03|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|2|2|3|2.5|||||||||4|4|2|3.33||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red||Volunteer: Lost contact with child/agency|87.1||2|2|2|2|F|Black||18||Mother|28208|One Parent: Female|Unknown||No||Self|General Community||Enrollment|F|Black||48|29715|Some College|Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500187758|31|0|2|500189225|31|0|2|500038037|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|189334||4|3|45
502172536|BBBS of Greater Charlotte|Main Office|C|Active|2010-10-13|NaT|Followup|2011-10-13|2011-09-13|Complete|Early|4|4|4|2|3|4|3.5|3|2|4|3|1|1|2.33|50.21|3|3|3|3|3|4|3.17|2|4|4|2|2|4|3|5.67|4|4|4|4|4|4|4|4|0|4|4|3|4|3.75|5|4|4|4|4.25|-11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|4|4|4|4|2|3|33.33|2|2|2|2|0|4|4||||Green|||77.1||1|1|1|1|F|Black||17|No|Mother|28269|Two Parent|Unknown||Yes||Relative|General Community||Match Support|F|Multi-race (Asian & White)||33|28205|Masters Degree|Married|Finance: Economist|28223|7|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502172965|31|0|2|501279665|37|0|2|500475431|2||-2||2|1|||-2||-2|0|3|||129|1|||1|190348|184611|4|3|45
501201092|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-26|2012-04-30|Followup|2011-08-26|2011-08-29|Complete|Done|3|2|4|2|2|4|2.83|||||||||3|3|3|4|4|4|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Red||Volunteer: Moved|44.1||1|1|1|1|M|White||20|No|Mother|28105|One Parent: Female|Unknown||No||Relative|General Community||Match Support|M|White||35|28270|Bachelors Degree|Single|Tech: Engineer|48121|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501201366|1|0|1|501285276|1|0|1|500280817|2||-2||4|3|||-2||-2|0|3|||7464|9|||1|191026||4|3|45
501670169|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-30|2012-04-04|Followup|2011-09-30|2011-09-13|Complete|Early|4|2|4|2|3|3|3|4|4|4|4|4|4|4|-25|2|2|3|2|3|3|2.5|2||4|||4|||4|4|4|4|4|4|3|3.67|8.99|3|3|3|4|3.25|4|2|4|5|3.75|-13.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3.67|8.99|3|3|3|4|2|3|0|2|2|1|1|100|4|4||||Green||Volunteer: Time constraint|30.1||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||Neighbor/Friend|General Community||Match Support|F|Black||32|28269||Single|Consultant|28209|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501670507|31|0|2|501466072|31|0|2|500379969|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|191050|2678|4|3|45
502188863|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2013-10-31|Baseline|2010-10-15|2010-12-31|Complete|Done|4|2|3|2|3|3|2.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1|||||||||Red|Project Big|Volunteer: Moved|34||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|M|Some Other Race||30|28202|Some College|Single|Tech: Support, Writing|28210|0|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502189292|31|0|1|502288935|41|0|1|500498784|2||-2||4|3|500004640|500004640|-2|500004640|-2|0|10|||46|2|||1|191872|-1|4|3|44
502358538|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-17|2011-10-26|Baseline|2010-10-15|2010-11-17|Complete|Done|4|4|4|4|3|3|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green||Child/Family: Moved|11.3||1|1|1|1|M|White||18|No|Mother|28025|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||68|28107||Married|Retired||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500002335|501519460|1|0|1|502078043|1|0|1|500481260|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|192065|-1|4|3|44
501829369|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-03|2012-01-10|Followup|2011-08-03|2011-10-18|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|29.2|Y|1|1|1|1|M|White||16|No|Mother|28027|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||61|28025||Married|Medical: Doctor, Provider||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|501829737|1|0|1|501687434|1|0|1|500376549|2||500003586||4|1|||-2||-2|0|10|||7464|9|||1|192340||4|0|45
502260656|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-18|2013-03-19|Followup|2011-10-18|2011-12-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Moved|29||2|2|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28078|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||33|28078|Associate Degree|Married|Education: Teacher Asst/Aid||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502261088|38|0|2|502249984|1|0|2|500475564|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|192420|170947|4|1|45
502185085|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-30|2011-05-02|Baseline|2010-10-19|2010-10-30|Complete|Done|4|2|3|2|3|3|2.83|||||||||4|4|4|4|4|3|3.83|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow||Child: Lost interest|6||1|1|2|2|M|White||16|No|Mother|28031|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||53|28117|Bachelors Degree|Married|Real Estate: Realtor|28031|0|0|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|277|60|598|500000170|500010355|502185514|1|0|1|502335257|1|0|1|500482493|2||-2||4|2|||-2|500000294, 500004901|-2|6854|8|||7464|9|||1|193379|-1|4|3|44
501810015|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-19|2012-02-09|Followup|2011-10-19|2011-11-03|Complete|Done|2|2|4|1|3|3|2.5|||||||||3|4|3|3|3|3|3.17|||||||||3|3|3|3||||||3|4|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|3|3.5|||||1|1||||4|4||||Green||Child/Family: Unrealistic expectations|27.7||1|1|2|2|M|Hispanic||15|No|Mother|28210|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501810370|3|0|1|501646021|3|0|1|500391598|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|194045||4|3|45
502338222|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2012-09-26|Baseline|2010-10-20|2010-10-27|Complete|Done|4|3|3|2|4|4|3.33|||||||||3|3|3|3|3|3|3|||||||||3|3|3|3||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1|||||||||Red|Project Big|Volunteer: Lost contact with child/agency|23||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Enrollment|F|Black||43|28105|Some College|Single|Business: Mgt, Admin|28226|11|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502338658|31|0|2|502255795|31|0|2|500483087|2||500004641||4|3|500004640|500004640|-2|500004640|-2|0|4|||7496|10|||1|194047|-1|4|3|44
500382177|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-18|2015-08-25|Followup|2011-09-18|2011-09-26|Complete|Done|3|2|2|3|3|3|2.67|||||||||3|4|4|3|2|3|3.17|||||||||4|4|4|4||||||3|3|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|107.2||1|1|2|2|M|Black||16||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||43|28215|Bachelors Degree|Single|Finance: Banking|28262|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|500382427|31|0|1|500188566|31|0|1|500122093|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|194049||4|3|45
502290880|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-20|2014-03-31|Followup|2011-10-20|2012-01-04|Expired|Late||||||||4|3|3|1|4|4|3.17|||||||||3|4|4|3|3|4|3.5||||||4|4|4|4|||||||5|4|5|4|4.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|4|3||||2|2|||||||Green|Project Big|Child/Family: Time constraints|41.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|M|White||35|28202|Bachelors Degree|Single|Real Estate: Realtor|28208|2|10|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502291312|31|0|1|502261364|1|0|1|500471473|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7496|10|||1|194052|179708|4|0|45
502338225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2016-05-26|Baseline|2010-10-20|2010-10-27|Complete|Done|3|2|3|1|4|4|2.83|||||||||2|3|2|2|3|3|2.5|||||||||3|3|3|3||||||2|3|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1|||||||||Yellow|Project Big|Volunteer: Lost contact with child/agency|67||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|White||33|28227|Bachelors Degree|Single|Unknown||9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502338658|31|0|2|502312449|1|0|2|500483095|2||500004641||4|2|500004640|500004640|-2|500004640|-2|0|4|||7496|10|||1|194054|-1|4|3|44
501123191|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-20|2015-12-21|Followup|2011-10-20|2011-11-09|Complete|Done|4|4|4|2|4|4|3.67|||||||||2|4|3|4|2|2|2.83|||||||||4|4|4|4||||||5|2|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||2|4|3|3||||||4|2|3|||||1|1||||4|4||||Green||Child/Family: Moved|62||2|2|1|1|F|Black||15|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||48|28210|Some College|Single|Human Services||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500915629|31|0|2|502153920|1|0|2|500478644|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|194321||4|3|45
502307545|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2011-10-25|Baseline|2010-10-20|2010-10-27|Complete|Done|3|3|3|2|3|3|2.83|||||||||2|3|3|3|3|3|2.83|||||||||3|3|3|3||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|1|1.5|||||1|1|||||||||Yellow|Project Big|Volunteer: Lost contact with child/agency|11.9||2|2|1|1|F|Hispanic||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Hispanic||33|28216|Some College|Widowed|Retail: Mgt||5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011184|502307977|3|0|2|502172480|3|0|2|500483395|2||500004641||4|2|500004640|500004640|-2|500004640|-2|0|4|||7496|10|||1|194334|-1|4|3|44
502304267|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-28|2012-10-10|Baseline|2010-10-20|2010-10-28|Complete|Done|3|1|2|1|1|2|1.67|||||||||2|2|3|4|2|3|2.67|||||||||3|4|2|3||||||5|4|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|2|2.5|||||1|1|||||||||Red||Volunteer: Moved|23.4||2|2|1|1|M|White||16|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||32|28270|Masters Degree|Living w/ Significant Other|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|502304699|1|0|1|502301421|1|0|1|500483429|2||-2||4|3|||-2||-2|0|10|||46|2|||1|194371|-1|4|3|44
502063945|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-21|2016-08-05|Followup|2011-10-21|2012-01-05|Expired|Late||||||||3|3|3|2|2|3|2.67|||||||||2|3|3|1|3|2|2.33||||||3|2|2|2.33|||||||3|2|4|2|2.75||||||||||4|4|4|4|4|3|2|3.57||||||3|4|3|3.33|||||1|4|2.5||||2|2|||||||Yellow||Volunteer: Time constraint|69.5||1|1|1|1|M|White||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community||Match Support|M|White||37|28205||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502064367|1|0|1|502295138|1|0|1|500478943|2||500004641||4|2|||-2||-2|0|5|||7496|10|||1|194859|189168|4|0|45
502310004|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-26|2014-05-01|Baseline|2010-10-21|2010-10-26|Complete|Done|4|4|4|4|3|3|3.67|||||||||2|3|4|4|3|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Yellow|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|42.2||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||No||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Enrollment|F|White||37|28078||Single|Business||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502310436|31|0|2|502331000|1|0|2|500483762|2||500003586||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7496|10|||1|194875|-1|4|3|44
502247579|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-30|2011-10-25|Baseline|2010-10-21|2010-10-30|Complete|Done|4|3|3|2|3|4|3.17|||||||||2|3|2|2|2|3|2.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Yellow|Amachi, Project Big, Project Big AND Amachi|Volunteer: Lost contact with child/agency|11.8||2|2|1|1|F|Black||15|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||29|28203||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011184|502248010|31|0|2|502322424|1|0|2|500483853|2||500004772||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7496|10|||1|194970|-1|4|3|44
502307478|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2012-04-30|Baseline|2010-10-21|2010-12-31|Complete|Done|3|2|3|2|3|3|2.67|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||1|1|1|1|1|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Red|Project Big|Volunteer: Moved|16||1|1|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Enrollment|M|Black||40|28215|Some College|Married|Transport: Driver||3|0|Michael Baisden|Media|Big|General Community||Match Support|277|60|598|500000170|500013709|502307910|31|0|1|502035292|31|0|1|500503967|2||||4|3|500004640|500004640|-2||-2|0|4|||11146|1|||1|195055|-1|4|3|44
500186133|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-14|2016-06-28|Followup|2011-10-14|2011-12-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|140.5||1|1|1|1|M|White||18||Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||51|28262|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500187724|1|0|1|500188930|1|0|1|500036930|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|195764||4|1|45
501575257|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-18|2013-09-24|Followup|2011-03-18|2011-03-11|Complete|Done|3|1|1|1|2|3|1.83|||||||||2|4|3|1|4|3|2.83|||||||||4|4|4|4||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|54.2||1|1|1|1|M|Black||15|No|Mother|28079|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||38|28079||Married|Law: Police Officer|28211|5|0|Recruitment Event|Self|Big|General Community||Enrollment|277|60|598|500000170|500004169|501575553|31|0|1|501234758|1|0|1|500348757|2||-2||4|3|||-2||-2|0|10|||7458|9|||1|196101||4|3|45
500185628|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-09|2012-08-30|Followup|2011-08-09|2011-08-22|Complete|Done|3|4|4|4|3|3|3.5|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||4|3|2|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|72.7||2|2|2|2|M|American Indian or Alaska Native||22||Mother|28031|Other/Unknown|Unknown||No||Neighbor/Friend|General Community||Match Support|M|White||51|28078|Bachelors Degree|Married|Business: Sales|28269|0|6|Igniting Breakfast|Special Event|Big|General Community|mentor2.0, mentor2.0 2015|RTBM|277|60|598|500000170|500008321|500187262|6|0|1|500190654|1|0|1|500117464|2||||4|3|||-2|500014505, 500015184|-2|0|8|||17266|8|||1|196238||4|3|45
501611456|BBBS of Greater Charlotte|Main Office|C|Active|2010-05-28|NaT|Followup|2011-05-28|2011-06-27|Complete|Done|4|4|4|1|4|4|3.5|||||||||1|4|4|2|2|4|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|||81.6||1|1|1|1|M|Black||15|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black|Other African|32|28262||Married|Law: Police Officer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501611776|31|0|1|501876475|31|31|1|500450969|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|196311||4|3|45
502307352|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-22|2011-07-28|Baseline|2010-10-25|2010-11-22|Complete|Done|3|3|3|3|3|3|3|||||||||3|3|3|3|3|3|3|||||||||3|4|3|3.33||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Green|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|8.1||2|2|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big AND Amachi|Match Support|F|Black||34|28208|PHD|Single|Medical: Doctor, Provider||1|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011184|502307784|31|0|2|502217265|31|0|2|500485187|2||500004772||4|1|500000294, 500004640, 500004901|500004901|-2|500004640|-2|0|4|||7464|9|||1|196663|-1|4|3|44
502310004|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-26|2014-05-01|Followup|2011-10-26|2011-12-13|Declined|Late||||||||4|4|4|4|3|3|3.67|||||||||2|3|4|4|3|4|3.33||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Yellow|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|42.2||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||No||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Enrollment|F|White||37|28078||Single|Business||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502310436|31|0|2|502331000|1|0|2|500483762|2||500003586||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7496|10|||1|197128|194875|4|1|45
501669649|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-26|2012-03-31|Followup|2011-10-26|2011-12-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|29.1||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Enrollment|M|Black||67|28262||Married|Business: Mgt, Admin||32|0|Mayfield Memorial|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013709|501669987|31|0|1|501818546|31|0|1|500388262|2||-2||4|3|||-2||-2|6854|8|||9212|7|||1|197586||4|1|45
500186428|BBBS of Greater Charlotte|Main Office|C|Completed|2005-10-03|2013-09-30|Followup|2011-10-03|2011-10-28|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|95.9||1|2|2|3|M|Black||21||Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||40|28211|Bachelors Degree|Single|Unknown||0|0|Brochure|Media|Big|General Community||Match Support|277|60|598|500000170|500004169|500187986|31|0|1|500189441|1|0|1|500044683|2||-2||4|1|||-2||-2|0|10|||127|1|||1|197588||4|1|45
500826594|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-21|2016-06-15|Followup|2011-08-21|2011-08-15|Complete|Done|3|2|3|2|3|2|2.5|||||||||3|3|3|3|3|3|3|||||||||4|4|3|3.67||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|105.8||1|1|1|1|M|Black||18|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Some Other Race||36|28209|||Business: Sales||0|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|1|500920342|41|0|1|500185735|2||-2||4|1|||-2||-2|0|5|||6450|12|||1|197658||4|3|45
500185734|BBBS of Greater Charlotte|Main Office|C|Completed|2003-10-15|2013-08-15|Followup|2011-10-15|2011-10-19|Complete|Done|2|2|3|2|3|3|2.5|||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||3|3|3|3|||||||||||||2|2|||||||||Red||Child: Graduated|118||1|1|1|1|F|Black||21||Mother|28203|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|White||45|28202|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187476|31|0|2|500188688|1|0|2|500036688|2||-2||4|3|||-2||-2|0|8|||7464|9|||1|197675||4|3|45
500970264|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2013-06-17|Followup|2011-10-27|2012-01-05|Declined|Late||||||||4|3|3|2|3|3|3|||||||||2|4|3|3|2|3|2.83||||||4|4|4|4|||||||2|3|3|3|2.75||||||||||4|4|4|4|4|4||||||||4|4|4|4|||||3|3|3||||2|2|||||||Red|Amachi|Volunteer: Lost contact with child/agency|31.7||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Enrollment|M|Black||44|28269|Some High School|Single|Insurance||0|2|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|1|502250629|31|0|1|500478922|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||12183|14|1209|1|1|198038|189150|4|1|45
502338222|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2012-09-26|Followup|2011-10-27|2012-01-11|Expired|Late||||||||4|3|3|2|4|4|3.33|||||||||3|3|3|3|3|3|3||||||3|3|3|3|||||||3|3|4|3|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|2|2||||1|1|||||||Red|Project Big|Volunteer: Lost contact with child/agency|23||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Enrollment|F|Black||43|28105|Some College|Single|Business: Mgt, Admin|28226|11|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502338658|31|0|2|502255795|31|0|2|500483087|2||500004641||4|3|500004640|500004640|-2|500004640|-2|0|4|||7496|10|||1|198421|194047|4|0|45
502338225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2016-05-26|Followup|2011-10-27|2012-01-11|Expired|Late||||||||3|2|3|1|4|4|2.83|||||||||2|3|2|2|3|3|2.5||||||3|3|3|3|||||||2|3|2|3|2.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|3|2.5||||1|1|||||||Yellow|Project Big|Volunteer: Lost contact with child/agency|67||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|White||33|28227|Bachelors Degree|Single|Unknown||9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502338658|31|0|2|502312449|1|0|2|500483095|2||500004641||4|2|500004640|500004640|-2|500004640|-2|0|4|||7496|10|||1|198431|194054|4|0|45
500930976|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-13|2013-04-26|Followup|2011-08-13|2011-10-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|56.4||1|1|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|Y|No||Service Organization|General Community||Match Support|F|Black||66|28205|Masters Degree|Single|Self-Employed, Entrepreneur||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500931243|31|0|2|501176751|31|0|2|500280106|2||-2||4|1|||-2||-2|0|11|||46|2|||1|198657||4|1|45
502304267|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-28|2012-10-10|Followup|2011-10-28|2011-10-03|Complete|Early|4|2|4|2|3|3|3|3|1|2|1|1|2|1.67|79.64|4|4|4|2|3|4|3.5|2|2|3|4|2|3|2.67|31.09|2|4|4|3.33|3|4|2|3|11|3|4|4|4|3.75|5|4|3|4|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|4|3|3.5|3|2|2.5|40|1|1|1|1|0|4|4||||Red||Volunteer: Moved|23.4||2|2|1|1|M|White||16|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||32|28270|Masters Degree|Living w/ Significant Other|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|502304699|1|0|1|502301421|1|0|1|500483429|2||-2||4|3|||-2||-2|0|10|||46|2|||1|198914|194371|4|3|45
502374716|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-11|2012-09-27|Baseline|2010-10-28|2010-11-11|Complete|Done|4|4|4|3|2|3|3.33|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2|||||||||Green|Project Big|Volunteer: Moved|22.5||2|2|1|1|M|Hispanic|Mexican|16|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Hispanic||38|28204||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502375154|3|10|1|502014837|3|0|1|500491463|2||500004641||4|1|500004640||-2|500004640|-2|0|4|||7496|10|||1|199086|-1|4|3|44
502255225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-08|2016-08-26|Baseline|2010-10-28|2010-11-08|Complete|Done|2|2|2|4|1|4|2.5|||||||||2|3|3|2|2|3|2.5|||||||||4|3|3|3.33||||||5|3|5|3|4|||||||4|3|4|4|4|4|4|3.86||||||||||4|4|4|4||||||1|1|1|||||1|1|||||||||Red||Volunteer: Moved|69.6||1|1|1|1|M|Hispanic||15||Mother|28212|One Parent: Female|Unknown||No|Spanish Radio|Media|General Community||Match Support|M|White||33|28226|Bachelors Degree|Single|Education: Teacher||3|0|Spanish Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502255655|3|0|1|502312682|1|0|1|500487118|2||-2||4|3|||-2||-2|7068|1|||11662|1|||1|199091|-1|4|3|44
502307403|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-30|2011-02-16|Baseline|2010-10-28|2010-11-30|Complete|Done|4|3|4|2|4|3|3.33|||||||||2|2|3|3|3|3|2.67|||||||||3|3|3|3||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Project Big|Volunteer: Moved|2.6||2|2|1|1|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Asian||28|28202|Bachelors Degree|Single|Finance|28202|0|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502307835|31|0|1|502312010|4|0|1|500487319|2||500004641||4|1|500004640|500004640, 500005291|-2||-2|0|4|||7462|13|||1|199366|-1|4|3|44
501300013|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-14|2012-05-01|Followup|2011-08-14|2011-10-29|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Agency: Challenges with program/partnership|44.6||2|2|2|2|F|Black||17|Yes|GrandMother|28273|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||40|28277|Associate Degree|Single|Unknown||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500003657|500561354|31|0|2|500188952|31|0|2|500281427|2||-2||4|1|500000294|500000294|-2||-2|7294|13|||7464|9|||1|199573||4|0|45
500970495|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-10|2017-03-09|Followup|2011-09-10|2011-09-06|Complete|Done|3|2|2|2|3|2|2.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|101.9||3|3|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$35,000 to $39,999||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black|Other African|44|28212||Single|Consultant||1|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500970766|31|0|2|500965698|31|31|2|500285645|2||-2||4|2|||-2||-2|7294|13|||46|2|||1|199909||4|3|45
501201068|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2012-08-29|Followup|2011-10-30|2011-12-15|Complete|Late|3|3|4|3|4|4|3.5|3|2|3|2|4|4|3|16.67|2|4|3|3|3|4|3.17|2|4|4|2|2|4|3|5.67|4|3|3|3.33|4|4|4|4|-16.75|4|4|5|4|4.25|4|4|5|3|4|6.25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|3|3|3|2|2|2|50|2|2|1|1|100|4|4||||Green||Child/Family: Lost contact with volunteer/agency|34||1|1|1|1|M|Black||21|No|Mother|28215|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||60|28262|Masters Degree|Single|Tech: Engineer||5|0|AA Task Force|Service Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501201342|31|0|1|501771844|31|0|1|500396764|2||-2||4|1|||-2|500000294|-2|6854|8|||9226|6|||1|199936|5730|4|3|45
500186853|BBBS of Greater Charlotte|Main Office|C|Completed|2004-11-04|2012-01-27|Followup|2011-11-04|2011-12-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|86.7||1|1|1|1|M|Black||21||Mother|28210|Other/Unknown|Unknown||No||Self|General Community||Match Support|M|Black||36|28203|Bachelors Degree||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500264223|31|0|1|500189632|31|0|1|500037741|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|199999||4|1|45
501342393|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-22|2014-06-06|Followup|2011-10-22|2011-11-11|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|2|2|||||2|2||||4|4||||Green||Child: Lost interest|67.4||1|1|1|1|F|White||19|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Business: Sales||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501342672|1|0|2|501210017|1|0|2|500293459|2||-2||4|1|||-2||-2|0|10|||46|2|||1|200029||4|3|45
501309634|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-12|NaT|Followup|2011-09-12|2011-09-13|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||102.1||1|1|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||46|27704|Associate Degree|Divorced|Medical: Admin||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501309912|31|0|2|501046221|31|0|2|500281317|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7462|13|||1|200293||4|3|45
500741571|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-15|2012-01-10|Followup|2011-08-15|2011-10-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|52.9||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Some Other Race||31|28262|||Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500002335|500724899|31|0|1|500938541|41|0|1|500187546|2||-2||4|1|||-2||-2|0|10|||46|2|||1|200544||4|0|45
501195410|BBBS of Greater Charlotte|Main Office|C|Active|2008-08-15|NaT|Followup|2011-08-15|2011-08-15|Complete|Done|4|3|3|2|3|||||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|||103||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Asian||35|28210|Bachelors Degree|Married|Business: Sales|28217|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501195684|31|0|1|501277677|4|0|1|500278978|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|200552||4|3|45
501234606|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-16|NaT|Followup|2011-09-16|2011-11-01|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||101.9||1|1|1|1|F|Black||16|No|Mother|28216|Grandparents|Unknown||No|TV|Media|General Community||Match Support|F|Black||42|28212|Bachelors Degree|Single|Unknown|28202|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501234882|31|0|2|501233675|31|0|2|500287478|2||-2||2|1|||-2||-2|56|1|||7464|9|||1|201197||4|1|45
501023408|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-05|NaT|Followup|2011-11-05|2011-10-18|Complete|Early|4|1|4|2|3|3|2.83|||||||||4|3|4|3|4|4|3.67|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||100.3||1|1|1|1|M|Hispanic|Other South American|17|No|Mother|28273|One Parent: Female|Less than $10,000||Yes||Self|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501023677|3|15|1|501356600|1|0|1|500296545|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|201433||4|3|45
500399844|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-20|2017-02-24|Followup|2011-08-20|2011-09-17|Complete|Done|4|1|4|1|4|4|3|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|1|3||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|114.2||1|2|1|2|F|Black||16||Mother|28208|One Parent: Female|Unknown||No||School|General Site||Match Support|F|White||35|28210|Bachelors Degree|Single|Business: Mgt, Admin|29715|0|0|Radio|Media|Big|General Site||Match Support|277|60|598|500000170|500008321|500400094|31|0|2|500188569|1|0|2|500190707|2||-2||4|3|||-1||-1|0|4|||131|1|||1|203376||4|3|45
501809541|BBBS of Greater Charlotte|Main Office|C|Active|2009-08-07|NaT|Followup|2011-08-07|2011-08-07|Complete|Done|4|2|4|2|4|4|3.33|||||||||3|3|4|3|3|3|3.17|||||||||4|3|3|3.33||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||91.3||1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||49|28031|Bachelors Degree|Married|Transport: Pilot|40223|9|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501809896|36|0|1|501620528|1|0|1|500375025|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|204813||4|3|45
502255225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-08|2016-08-26|Followup|2011-11-08|2011-11-06|Complete|Done|4|1|3|1|4|4|2.83|2|2|2|4|1|4|2.5|13.2|1|2|4|3|3|4|2.83|2|3|3|2|2|3|2.5|13.2|4|4|2|3.33|4|3|3|3.33|0|5|3|5|3|4|5|3|5|3|4|0|2|4|4|4|4|4|4|3.71|4|3|4|4|4|4|4|3.86|-3.89|4|4|4|4|4|4|4|4|0|2|2|2|1|1|1|100|1|1|1|1|0|4|4||||Red||Volunteer: Moved|69.6||1|1|1|1|M|Hispanic||15||Mother|28212|One Parent: Female|Unknown||No|Spanish Radio|Media|General Community||Match Support|M|White||33|28226|Bachelors Degree|Single|Education: Teacher||3|0|Spanish Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502255655|3|0|1|502312682|1|0|1|500487118|2||-2||4|3|||-2||-2|7068|1|||11662|1|||1|204974|199091|4|3|45
502295599|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2012-01-13|Baseline|2010-11-08|2010-11-18|Complete|Done|4|2|4|2|4|4|3.33|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||2|4|3|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||4|3|3.5|||||1|1|||||||||Red||Volunteer: Lost contact with child/agency|13.8||1|1|1|1|F|Black||17|No|Mother|28211|One Parent: Female|Unknown||No|AARTF|BBBS Board/Staff|General Community||Enrollment|F|White||28|28277||Single|Finance: Accountant||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502296031|31|0|2|502306663|1|0|2|500491842|2||-2||4|3|||-2||-2|7294|13|||7496|10|||1|205074|-1|4|3|44
501101153|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-30|2013-08-30|Followup|2011-09-30|2011-10-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Severity of challenges|59||1|2|2|3|M|Black||19||Mother|28205|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||62|28214|Bachelors Degree|Married|Human Services: Non-Profit|28214|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501101427|31|0|1|500789916|1|0|1|500293277|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|205256||4|1|45
501092957|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-09|2014-05-15|Followup|2011-11-09|2012-01-17|Blank|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|42.2||2|2|1|1|M|Black||17|No|Mother|28027|One Parent: Female|$30,000 to $34,999||No|Radio|Media|General Community||Match Support|M|White||44|28269||Married|Finance: Banking||5|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|501093231|31|0|1|502294662|1|0|1|500484597|2||-2||4|1|||-2||-2|55|1|||7459|10|||1|205698||4|3|45
500998929|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-19|2011-08-30|Baseline|2010-11-09|2010-11-19|Complete|Done|4|4|4|2|4|4|3.67|||||||||1|3|2|2|1|3|2|||||||||4|4|4|4||||||1|5|2|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|2|2|||||1|1|||||||||Green|Amachi|Volunteer: Moved|9.3||1|1|1|1|F|Black||21|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|F|White||29|28204|Bachelors Degree|Single|Medical: Nurse|28202|0|0|Big Champions|Other Big|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008629|500999202|31|0|2|502332678|1|0|2|500497432|2||-2||4|1|500000294|500000294|-2|500000294, 500004640|-2|0|10|||7461|12|||1|205735|-1|4|3|44
502308593|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-23|2015-05-28|Baseline|2010-11-10|2010-11-23|Complete|Done|4|2|3|1|3|4|2.83|||||||||3|3|4|4|3|3|3.33|||||||||3|2|3|2.67||||||3|4|5|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|3|2.5|||||1|1|||||||||Red||Child/Family: Moved|54.1||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||40|28278|Bachelors Degree|Married|Tech: Computer/Programmer||3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502309025|31|0|1|502262702|31|0|1|500492994|2||-2||4|3|||-2||-2|0|10|||12183|14|1209|1|1|206463|-1|4|3|44
500185630|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-26|2012-09-06|Followup|2011-09-26|2011-09-26|Complete|Done|4|4|3|3|3|4|3.5|||||||||2|4|3|3|4|4|3.33|||||||||4|4|4|4||||||2|5|3|4|3.5|||||||3|3|4|3|4|4|4|3.57||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child/Family: Time constraints|71.4||3|3|2|2|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||39|28211|High School Graduate|Single|Finance: Banking|28208|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008629|500187264|31|0|2|500542491|31|0|2|500122710|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|206663||4|3|45
500867579|BBBS of Greater Charlotte|Main Office|C|Completed|2007-09-22|2013-04-02|Followup|2011-09-22|2011-11-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|66.3||1|1|1|1|M|Black||23|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|No||Faith Organization|General Community|Amachi|Match Support|M|Black||42|28269||Single|Finance: Banking||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|500867843|31|0|1|500577903|31|0|1|500195387|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|206665||4|1|45
501288021|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-27|2016-02-01|Followup|2011-08-27|2011-11-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|89.2||1|1|1|1|F|Black||16|No|Mother|28211|Two Parent|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28027|PHD|Single|Education: College Professor|27411|1|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501288299|31|0|2|501249338|31|0|2|500281778|2||-2||4|1|||-2||-2|0|10|||46|2|||1|207115||4|0|45
502374716|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-11|2012-09-27|Followup|2011-11-11|2011-11-13|Complete|Done|2|1|3|2|3|4|2.5|4|4|4|3|2|3|3.33|-24.92|2|3|4|1|2|4|2.67|2|3|3|2|2|3|2.5|6.8|4|3|3|3.33|4|4|4|4|-16.75|4|3|3|3|3.25|3|3|4|3|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|4|4|3.67|-9.26|4|4|4|4|4|4|0|1|1|2|2|-50|4|4||||Green|Project Big|Volunteer: Moved|22.5||2|2|1|1|M|Hispanic|Mexican|16|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Hispanic||38|28204||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502375154|3|10|1|502014837|3|0|1|500491463|2||500004641||4|1|500004640||-2|500004640|-2|0|4|||7496|10|||1|207512|199086|4|3|45
501614040|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-11|2013-02-28|Followup|2011-11-11|2011-11-11|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|5|2|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|39.6||1|1|1|1|M|Hispanic||16|No|Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||29|28273|||Facilities/Maintenance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|501614360|3|0|1|501864748|1|0|1|500404360|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|208113||4|3|45
500867581|BBBS of Greater Charlotte|Main Office|C|Completed|2007-09-28|2014-02-06|Followup|2011-09-28|2011-11-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|76.3||1|1|2|2|M|Black||21|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999||No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||40|28269|Masters Degree|Single|Finance: Accountant|28255|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|500867843|31|0|1|500708515|1|0|1|500195388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|208337||4|1|45
501365904|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-20|2012-09-05|Followup|2011-04-20|2011-05-02|Complete|Done|3|3|3|1|4|3|2.83|||||||||3|4|4|2|3|4|3.33|||||||||4|4|3|3.67||||||4|5|4|5|4.5|||||||4|4|4|3|3|3|2|3.29||||||||||3|4|3|3.33||||||2|2|2|||||1|1|||||||||Yellow||Child/Family: Moved|40.5||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown|Y|No||Self|General Community||Enrollment|M|Black||48|28269|Some College|Married|Business: Engineer|28262|20|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501366183|31|0|1|501459709|31|0|1|500353421|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|208662||4|3|45
500186926|BBBS of Greater Charlotte|Main Office|C|Completed|2004-08-30|2011-12-21|Followup|2011-08-30|2011-09-07|Complete|Done|3|3|3|3|3|3|3|||||||||3|3|3|3|4|3|3.17|||||||||4|3|3|3.33||||||3|4|3|3|3.25|||||||4|4|4|3|3|4|3|3.57||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Volunteer: Lost contact with child/agency|87.7||1|1|1|1|M|Some Other Race||23|Yes|Mother|28213|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||60|28277|Bachelors Degree|Married|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500003657|500188133|41|0|1|500189699|31|0|1|500037812|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|208671||4|3|45
500383923|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-30|2012-08-30|Followup|2011-08-30|2011-10-19|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|72||1|1|2|2|M|Black||18||GrandMother|28205|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||66|28269||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500384165|31|0|1|500540549|31|0|1|500118470|2||-2||4|1|||-2||-2|0|8|||7464|9|||1|208682||4|1|45
501129781|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-15|2015-01-15|Followup|2011-11-15|2011-11-15|Complete|Done|4|1|4|1|4|4|3|||||||||3|4|4|4|1|4|3.33|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Green||Child: Family structure changed|50||1|2|4|6|F|Black||17||Mother|28217|Two Parent|Unknown||No||School|General Community||Match Support|F|Black||48|28273|Bachelors Degree|Married|Business: Mgt, Admin|28273|4|0|Recruitment Event|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500018987|501130055|31|0|2|500189245|31|0|2|500494855|2||-2||4|1|||-2||-2|0|4|||7459|10|||1|209384||4|3|45
500185972|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-01|2012-12-21|Followup|2011-09-01|2011-09-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|75.7||2|3|1|1|F|Black||22|Yes|Mother|28206|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|F|Black||38|28213|Bachelors Degree|Single|Education: Teacher|28202|2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187610|31|0|2|500492482|31|0|2|500120588|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|209649||4|1|45
502177629|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-30|2011-10-25|Baseline|2010-11-17|2010-11-30|Complete|Done|3|4|4|3|1|4|3.17|||||||||1|4|4|2|4|4|3.17|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1|||||||||Yellow||Volunteer: Lost contact with child/agency|10.8||1|1|1|1|M|Black||16|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||RTBM|M|White||59|28277|Associate Degree|Divorced|Unknown||0|0|CIAA Tournament|Special Event|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500011184|502178058|31|0|1|502247130|1|0|1|500495930|2||-2||4|2|||-2|500000294, 500004640|-2|0|10|||11248|8|||1|210517|-1|4|3|44
502295599|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2012-01-13|Followup|2011-11-18|2011-11-13|Complete|Done|4|3|4|1|3|4|3.17|4|2|4|2|4|4|3.33|-4.8|4|1|4|4|4|4|3.5|2|4|3|4|4|3|3.33|5.11|4|4|4|4|4|4|4|4|0|5|2|4|5|4|2|4|3|3|3|33.33|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3.5|14.29|1|1|1|1|0|4|4||||Red||Volunteer: Lost contact with child/agency|13.8||1|1|1|1|F|Black||17|No|Mother|28211|One Parent: Female|Unknown||No|AARTF|BBBS Board/Staff|General Community||Enrollment|F|White||28|28277||Single|Finance: Accountant||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502296031|31|0|2|502306663|1|0|2|500491842|2||-2||4|3|||-2||-2|7294|13|||7496|10|||1|211544|205074|4|3|45
502173821|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2014-08-29|Followup|2011-11-18|2012-01-05|Declined|Late||||||||4|1|1|1|4|4|2.5|||||||||3|4|4|3|3|4|3.5||||||4|4|4|4|||||||5|5|4|4|4.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|2|2||||1|1|||||||Red|Amachi|Volunteer: Time constraint|45.3||2|2|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||32|28262|Masters Degree|Single|Finance: Banking|28262|3|11|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502174240|31|0|2|502264706|1|0|2|500491573|2||500003586||4|3|500000294|500000294|-2|500000294, 500004640|-2|7016|11|||7464|9|||1|211735|148526|4|1|45
500186192|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2014-10-13|Followup|2011-11-18|2011-12-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|46.8||2|2|1|1|F|Black||20||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|Black||33|28208||Single|Service: Restaurant||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187762|31|0|2|502323059|31|0|2|500490136|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|211741||4|1|45
500998933|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-19|2013-12-06|Followup|2011-11-19|2012-01-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|36.6||1|1|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|F|White||37|28210|Masters Degree|Single|Medical|28210|1|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500015820|500999202|31|0|2|502274159|1|0|2|500497430|2||500003586||4|3|500000294|500000294|-2|500000294, 500004640|-2|0|10|||7496|10|||1|212848||4|1|45
500185723|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-05|2015-06-25|Followup|2011-09-05|2011-10-19|Complete|Done|4|2|4|4|3|4|3.5|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|81.6||2|2|1|1|M|Black||19||Mother|28214|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|M|Black||36|28214|Bachelors Degree|Single|Tech: Computer/Programmer|28147|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187335|31|0|1|501310677|31|0|1|500284133|2||-2||4|3|||-2||-2|6855|8|||7464|9|||1|212898||4|3|45
501716720|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-02|2017-02-06|Followup|2011-03-02|2011-05-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Cabarrus County|Child/Family: Lost contact with volunteer/agency|83.2||1|1|1|1|M|Black||15|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||52|28075||Married|Medical: Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501716992|31|0|1|501878786|31|0|1|500435676|2||500016307||4|3|500016374|500016374|-2|500016374|-2|6854|8|||7464|9|||1|213037||4|0|45
500931662|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-07|NaT|Followup|2011-09-07|2011-10-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||114.3||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$60,000 to $74,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||58|28270|Bachelors Degree|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500931932|31|0|1|500894084|1|0|1|500193824|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|213228||4|1|45
500480596|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-13|2014-01-16|Followup|2011-09-13|2011-09-15|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|Amachi|Child: Graduated|88.1||1|1|1|1|M|Black||21|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Married|Business: Sales|28203|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500480847|31|0|1|500491267|1|0|1|500120915|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|213342||4|3|45
500185846|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-28|2014-10-23|Followup|2011-09-28|2011-11-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|120.8||1|2|1|2|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||65|28256|Bachelors Degree||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187437|31|0|2|500188764|31|0|2|500038142|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|213343||4|1|45
500191820|BBBS of Greater Charlotte|Main Office|C|Completed|2005-09-30|2013-08-29|Followup|2011-09-30|2011-11-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|94.9|Y|2|2|2|2|M|Black||19||Mother|28227||Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||72|28214||Married|Retired||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500191823|31|0|1|500191501|31|0|1|500044434|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|213345||4|1|45
500871683|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-01|2016-02-22|Followup|2011-10-01|2011-11-21|Complete|Late|3|3|4|3|3|3|3.17|||||||||3|3|3|3|3|3|3|||||||||4|3|3|3.33||||||4|3|4|3|3.5|||||||4|4|4|3|3|3|3|3.43||||||||||4|4|3|3.67||||||2|2|2|||||1|1||||4|4||||Green|Amachi|Child: Graduated|100.7||1|1|1|1|M|Black||19|Yes|Aunt|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|M|White||46|28209|Masters Degree|Single|Self-Employed, Entrepreneur|28209|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500871952|31|0|1|500933829|1|0|1|500199601|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|213346||4|3|45
501340102|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-03|2013-04-25|Followup|2011-10-03|2011-11-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Time constraints|54.7||1|1|1|1|M|Multi-race (Black & Hispanic)||18|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||50|28269|Masters Degree|Married|Customer Service|28269|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340381|38|0|1|501316292|1|0|1|500287888|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|213347||4|1|45
501114443|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-08|2013-07-25|Followup|2011-10-08|2011-11-21|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|57.5||1|1|2|2|M|Black||22|No|Uncle|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||34|28205|Juris Doctorate (JD)|Married|Law: Lawyer||0|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501114708|31|0|1|501180846|1|0|1|500290376|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||46|2|||1|213348||4|3|45
501068953|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-06|2012-03-31|Followup|2011-10-06|2011-12-21|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|29.8||2|2|2|2|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||40|28262|Bachelors Degree|Married|Law: Paralegal|28280|4|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008629|501060469|31|0|2|500874318|31|0|2|500380111|2||-2||4|1|||-2||-2|34|2|||46|2|||1|214170||4|0|45
500826592|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-08|2016-10-18|Followup|2011-10-08|2011-11-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|84.3||3|3|1|1|F|Black||20|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|F|White||33|28277|Bachelors Degree|Living w/ Significant Other|Unknown|28209|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|2|501314246|1|0|2|500382768|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|214173||4|1|45
500713817|BBBS of Greater Charlotte|Main Office|C|Active|2009-10-30|NaT|Followup|2011-10-30|2011-11-11|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||2|4|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||88.5||2|2|1|1|M|Black||16||Mother|28216|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28078|||Medical: Pharmacist|28210|10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|500714084|31|0|1|501834795|1|0|1|500396466|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|214325||4|3|45
502308593|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-23|2015-05-28|Followup|2011-11-23|2012-01-05|Declined|Done||||||||4|2|3|1|3|4|2.83|||||||||3|3|4|4|3|3|3.33||||||3|2|3|2.67|||||||3|4|5|2|3.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|3|2.5||||1|1|||||||Red||Child/Family: Moved|54.1||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||40|28278|Bachelors Degree|Married|Tech: Computer/Programmer||3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502309025|31|0|1|502262702|31|0|1|500492994|2||-2||4|3|||-2||-2|0|10|||12183|14|1209|1|1|214453|206463|4|1|45
502294587|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-07|2011-03-04|Baseline|2010-11-24|2010-12-07|Complete|Done|2|4|4|4|3|3|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|3|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|1|2.67||||||3|4|3.5|||||2|2|||||||||Green||Volunteer: Moved|2.9||1|1|1|1|M|Black||21|No|Mother|28215|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||31|28204|Juris Doctorate (JD)|Single|Law: Lawyer|28280|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500010765|501712404|31|0|1|502389185|1|0|1|500499438|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|214956|-1|4|3|44
502274030|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-18|2012-05-31|Followup|2011-10-18|2012-01-02|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Moved|19.4||1|1|1|1|F|White||15|No|Mother|28270|One Parent: Female|Unknown||Yes||Relative|General Community||Enrollment|F|White||38|28205|Bachelors Degree|Married|Tech: Engineer||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502274462|1|0|2|502133187|1|0|2|500477736|2||-2||4|3|||-2||-2|0|3|||7464|9|||1|215294||4|0|45
500186692|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-11|2012-06-30|Followup|2011-09-11|2011-09-13|Complete|Done|3|3|4|2|3|3|3|||||||||3|3|3|3|4|4|3.33|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|33.6||7|8|1|1|F|Black||19|No|Mother|28270|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|White||50|28270|Some College|Single|Finance: Banking|28217|1|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500188059|31|0|2|501582415|1|0|2|500381441|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|215361||4|3|45
500186190|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-13|2014-08-20|Followup|2011-10-13|2011-11-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|118.2||1|1|2|2|F|Black||20||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187761|31|0|2|500189140|31|0|2|500037140|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|215390||4|1|45
500336002|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-29|2012-03-31|Followup|2011-11-29|2012-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Lost contact with child/agency|16||4|5|2|3|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|F|White||33|28202||Single|Business: Marketing||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013709|500293247|31|0|2|500801056|1|0|2|500490281|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|215749||4|1|45
501224282|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-16|2012-06-14|Followup|2011-10-16|2011-11-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Feels incompatible with child/family|43.9||2|2|1|1|F|Black||15|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||35|28215|Bachelors Degree|Single|Finance: Banking|28262|2|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501224558|31|0|2|501389463|31|0|2|500296679|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||7453|7|||1|215811||4|1|45
501253195|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-24|NaT|Followup|2011-10-24|2011-11-21|Complete|Done|3|2|2|2|3|2|2.33|||||||||3|3|3|3|3|3|3|||||||||4|4|3|3.67||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi||100.7||1|1|2|2|M|Black||15|Yes|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28203|Masters Degree|Single|Medical: Doctor, Provider|28211|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501253471|31|0|1|500395148|1|0|1|500282924|2||500003586||2|1|500000294||-2||-2|0|10|||7464|9|||1|215814||4|3|45
500185907|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2015-02-18|Followup|2011-10-29|2011-11-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|99.7||2|3|1|1|F|Black||19|Yes|Mother|28262|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||48|28212||Single|Medical: Healthcare Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187470|31|0|2|500697782|31|0|2|500134557|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|215818||4|1|45
501224287|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-30|2014-01-23|Followup|2011-10-30|2011-11-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|62.8||1|1|1|1|M|Black||19|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||43|28262|Bachelors Degree|Married|Customer Service|28211|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501224558|31|0|1|501343190|31|0|1|500298289|2||-2||4|3|500000294|500000294|-2|500000294|-2|5635|9|||2230|7|||1|215820||4|1|45
500252077|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-24|2016-01-20|Followup|2011-11-24|2011-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|85.8||3|3|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Tech: Computer/Programmer||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501750989|31|0|1|501365749|1|0|1|500317108|2||500003586||4|3|500000294|500000294|-2||-2|7295|11|||46|2|||1|215822||4|1|45
502280284|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-13|2013-07-31|Baseline|2010-11-30|2010-12-13|Complete|Done|4|3|3|2|4|4|3.33|||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Red|Project Big|Volunteer: Lost contact with child/agency|31.6||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|White||31|28205|Associate Degree|Married|Business: Human Resources||3|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502280719|31|0|2|502241391|1|0|2|500500329|2||500004641||4|3|500004640|500004640|-2|500004640|-2|0|10|||46|2|||1|216597|-1|4|3|44
500829028|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-30|NaT|Followup|2011-11-30|2011-11-10|Complete|Early|4|1|4|1|4|4|3|||||||||2|2|4|2|2|4|2.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||75.5||3|3|2|2|F|Black||17|No|Mother|28209|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||39|28210|Masters Degree|Single|Education|28212|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502254499|31|0|2|501978180|1|0|2|500498594|2||-2||2|1|||-2|500000294, 500004640|-2|0|10|||7464|9|||1|217216||4|3|45
502256918|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-07|2013-04-25|Baseline|2010-12-01|2010-12-07|Complete|Done|4|4|4|1|3|4|3.33|||||||||3|3|4|2|4|3|3.17|||||||||4|4|4|4||||||3|3|2|5|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|3|3|||||2|2|||||||||Red||Child/Family: Moved|28.6||1|1|1|1|M|Hispanic||16|No|Mother|28212|One Parent: Female|Unknown||No|Spanish Print|Media|General Community||Match Support|M|White||38|28209|Juris Doctorate (JD)|Single|Law||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502257350|3|0|1|502143354|1|0|1|500501039|2||-2||4|3|||-2||-2|7063|1|||7464|9|||1|217658|-1|4|3|44
501086649|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-20|2013-01-09|Followup|2011-11-20|2011-12-30|Declined|Done||||||||4|3|4|2|3|4|3.33|||||||||4|4|4|4|3|3|3.67||||||4|3|3|3.33|||||||5|4|4|5|4.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||4|4|4||||2|2|||||||Red||Volunteer: Feels incompatible with child/family|37.7||1|1|1|1|M|Black||21|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Relative|General Community||Match Support|M|White||39|28205|Bachelors Degree|Single|Transport: Pilot|30320|2|0|Other Church Partner|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500004169|501086923|31|0|1|501833794|1|0|1|500399391|2||-2||4|3|||-2||-2|0|3|||7453|7|||1|217677|385|4|1|45
500801567|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-26|2013-12-12|Followup|2011-10-26|2011-12-15|Complete|Late|3|4|3|3|3|3|3.17|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|49.5||2|2|1|1|M|Black||20||Mother|28213|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||62|28078|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500801835|31|0|1|501834907|1|0|1|500391790|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|217680||4|3|45
500970181|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-31|2012-08-29|Followup|2011-10-31|2011-10-20|Complete|Done|3|3|3|3|3|3|3|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||3|3||||Red||Child: Severity of challenges|58||1|1|1|1|M|Black|Other African|20|No|Mother|28208|One Parent: Female|$15,000 to $19,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||37|28210|Bachelors Degree|Single|Finance: Accountant||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|500970452|31|31|1|500969057|1|0|1|500203109|2||-2||4|3|||-2||-2|34|2|||46|2|||1|217732||4|3|45
500897065|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-17|2012-05-23|Followup|2011-09-17|2011-11-01|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|32.2||3|4|2|3|F|Black||18|Yes|Mother|28269|Other/Unknown|Unknown||No||Service Organization|General Community||Match Support|F|Black||34|28105|Bachelors Degree|Married|Education: Admin|28202|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500897335|31|0|2|501454753|31|0|2|500384418|2||-2||4|1|||-2||-2|0|11|||7464|9|||1|218019||4|1|45
502270499|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-28|2011-03-29|Baseline|2010-12-03|2010-12-21|Complete|Done|4|2|1|1|3|4|2.5|||||||||2|4|4|2|1|3|2.67|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Time constraint|3||2|2|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||67|28207|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011184|502231230|31|0|2|502376097|1|0|2|500501731|2||500003586||4|1||500000294|-2|500000294|-2|5635|9|||7464|9|||1|218599|-1|4|3|44
502307481|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2012-01-27|Baseline|2010-12-03|2010-12-31|Complete|Done|4|3|3|2|4|4|3.33|||||||||3|3|2|2|3|3|2.67|||||||||4|4|4|4||||||3|2|2|3|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Red|Project Big|Volunteer: Time constraint|12.9||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|RTBM|M|White||38|28205|Bachelors Degree|Married|Business: Sales||4|0|Other|Service Organization|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013709|502307910|31|0|1|502212397|1|0|1|500501813|2||500004641||4|3|500004640|500004640|-2|500004640|-2|0|4|||7452|6|||1|218679|-1|4|3|44
500958307|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-19|NaT|Followup|2011-09-19|2011-12-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi, Cabarrus County||113.9|Y|1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$40,000 to $44,999|Y|No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|Black||62|28213||Married|Finance: Economist||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500958577|31|0|1|500876132|31|0|1|500193868|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|219033||4|0|45
500186646|BBBS of Greater Charlotte|Main Office|C|Completed|2005-10-20|2013-09-23|Followup|2011-10-20|2011-12-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|95.1||3|3|3|3|F|Some Other Race||21||Mother|28217|Other/Unknown|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||39|28216|Some College||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500188044|41|0|2|500189263|31|0|2|500047741|2||-2||4|2|||-2||-2|0|8|||7464|9|||1|219104||4|1|45
501725162|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2016-10-14|Followup|2011-10-29|2011-12-06|Complete|Done|2|1|3|1|4|4|2.5|4|1|2|1|4|4|2.67|-6.37|2|4|3|3|3|2|2.83|3|4|2|3|3|3|3|-5.67|3|2|3|2.67|1|4|4|3|-11|2|5|3|4|3.5|5|1|5|5|4|-12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|2|3|4|4|2|3.33|-9.91|4|3|3.5|4|3|3.5|0|2|2|2|2|0|4|4||||Green||Agency: Challenges with program/partnership|83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501724831|39|0|1|501833178|1|0|1|500394157|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|219462|16143|4|3|45
500185721|BBBS of Greater Charlotte|Main Office|C|Completed|2003-12-03|2012-05-25|Followup|2011-12-03|2011-12-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|101.7||1|1|1|1|M|Black||22||Mother|28054|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||43|28207||Single|Unknown||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|500187333|31|0|1|500188678|1|0|1|500036678|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|219464||4|1|45
502256918|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-07|2013-04-25|Followup|2011-12-07|2011-12-05|Complete|Done|2|4|3|1|3|4|2.83|4|4|4|1|3|4|3.33|-15.02|2|3|3|2|3|3|2.67|3|3|4|2|4|3|3.17|-15.77|4|4|4|4|4|4|4|4|0|1|5|4|4|3.5|3|3|2|5|3.25|7.69|4|4|4|4|4|3|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|3|3|3.33|4|3|4|3.67|-9.26|4|4|4|3|3|3|33.33|1|1|2|2|-50|4|4||||Red||Child/Family: Moved|28.6||1|1|1|1|M|Hispanic||16|No|Mother|28212|One Parent: Female|Unknown||No|Spanish Print|Media|General Community||Match Support|M|White||38|28209|Juris Doctorate (JD)|Single|Law||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502257350|3|0|1|502143354|1|0|1|500501039|2||-2||4|3|||-2||-2|7063|1|||7464|9|||1|220020|217658|4|3|45
502138562|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-14|2013-06-06|Baseline|2010-12-07|2010-12-14|Complete|Done|2|3|4|3|1|1|2.33|||||||||1|2|1|4|4|4|2.67|||||||||3|3|3|3||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2|||||||||Green||Child: Lost interest|29.7||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||38|28216|Masters Degree|Single|Finance: Auditor|28217|3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500011746|502138991|31|0|1|502380370|31|0|1|500502780|2||-2||4|1|||-2||-2|0|10|||12183|14|||1|220057|-1|4|3|44
502129650|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-17|2012-09-27|Baseline|2010-12-07|2010-12-17|Complete|Done|4|4|4|4|4|4|4|||||||||1|4|3|4|1|4|2.83|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Yellow||Volunteer: Lost contact with child/agency|21.4||2|2|1|1|F|Black||17|No|GrandMother|28027|Grandparents|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|Black||29|28027|||Customer Service||0|0||High School Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|502130079|31|0|2|501733783|31|0|2|500502959|2||-2||4|2||500016374|-2||-2|0|10|||0|4|||1|220242|-1|4|3|44
502083429|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-11|2016-08-19|Baseline|2010-12-07|2012-02-11|Complete|Done|4|2|4|3|2|4|3.17|||||||||4|4|4|1|4|4|3.5|||||||||4|3|3|3.33||||||3|5|4|4|4|||||||4|2|4|4|4|4|3|3.57||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Moved|54.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Cabarrus County|Match Support|F|Black||29|28027|Bachelors Degree|Single|Education: Teacher||1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|502083853|31|0|2|502653045|31|0|2|500590992|2||-2||4|3||500016374|-2|500016374|-2|7016|11|||7464|9|||1|220254|-1|4|3|44
500186742|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-08|2016-06-30|Followup|2011-12-08|2011-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|66.7||4|4|1|1|M|Black||19|Yes|Mother|28227|One Parent: Female|Unknown|Y|No||School|General Community|Amachi|Match Support|M|Black||52|28227|Masters Degree|Married|Education: Teacher|28227|2|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|502397541|31|0|1|500501282|2||500003586||4|1|500000294|500000294|-2|500000294, 500004640|-2|0|4|||12183|14|635|1|1|220663||4|1|45
500717519|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-08|2013-08-29|Followup|2011-12-08|2012-02-10|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Lost interest|80.7||1|1|2|2|M|Black||20||Mother|28205|One Parent: Female|$20,000 to $24,999|Y|No||School|General Community||Match Support|M|Black||37|28269|Bachelors Degree|Married|Education: Admin||0|0|Yahoo!|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|500717786|31|0|1|500188838|31|0|1|500145722|2||-2||4|2|||-2||-2|0|4|||32|2|||1|221471||4|1|45
501796006|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-03|2011-12-20|Followup|2011-11-03|2011-12-20|Declined|Late||||||||3|4|4|2|3|4|3.33|||||||||2|4|4|4|2|4|3.33||||||4|4|4|4||||||||3|3|5|||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||4|2|3||||2|2|||||||Green||Volunteer: Time constraint|25.5||3|3|1|1|F|Black||17|No|Mother|28031|Two Parent|Unknown|Y|Yes||School|General Community||Match Support|F|White||37|28078|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011639|501489205|31|0|2|501621517|1|0|2|500396069|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|221480|6008|4|1|45
501347056|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2015-10-12|Followup|2011-12-12|2012-02-01|Complete|Late|4|4|4|2|3|4|3.5|||||||||1|4|4|1|4|2|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Child: Graduated|82||1|1|1|1|M|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28226|Bachelors Degree|Married|Tech: Engineer|28202|2|8|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|501347335|31|0|1|501217000|1|0|1|500322327|2||-2||4|2|||-2||-2|34|2|||7446|3|||1|221498||4|3|45
501363890|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-21|2012-08-29|Followup|2011-11-21|2012-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|45.2||1|1|2|2|M|Black||21|No|Mother|28216|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|M|Black||37|28213|Masters Degree|Single|Medical: Healthcare Worker||2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501356607|31|0|1|500189279|31|0|1|500315105|2||-2||4|2|||-2|500000294|-2|0|8|||7464|9|||1|221515||4|1|45
502290482|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-18|2011-10-25|Baseline|2010-12-09|2010-12-18|Complete|Done|4|1|4|1|4|4|3|||||||||3|4|3|2|4|4|3.33|||||||||4|4|4|4||||||2|3|4|2|2.75|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|3|2.5|||||2|2|||||||||Green||Volunteer: Moved|10.2||2|2|1|1|F|Black||18|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28202|Masters Degree||Finance: Banking||0|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500011184|502290914|31|0|2|501861156|1|0|2|500503975|2||-2||4|1|||-2|500000294, 500004640|-2|0|10|||7464|9|||1|221593|-1|4|3|44
501247286|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-14|2016-11-08|Followup|2011-05-14|2011-07-29|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|101.8||1|1|1|1|M|White||15|No|Father|28025|One Parent: Male|Unknown||No||Self|General Community|Cabarrus County|Enrollment|M|White||49|27103|Masters Degree|Single|Education: Teacher|27282|0|0|Other|Service Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500341682|1|0|1|501247141|1|0|1|500264655|2||-2||4|1||500016374|-2|500016374|-2|0|10|||7452|6|||1|221844||4|0|45
500337327|BBBS of Greater Charlotte|Main Office|C|Active|2006-12-14|NaT|Followup|2011-12-14|2012-01-23|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||123||2|3|4|5|M|Black||16||GrandMother|28208|Grandparents|Unknown||No||School|General Site||Match Support|M|Black||49|28217|Associate Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site||Match Support|277|60|598|500000170|500017732|500251937|31|0|1|500189300|31|0|1|500148262|2||-2||2|1|||-1||-1|0|4|||7464|9|||1|222171||4|3|45
501860373|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-16|2011-08-25|Baseline|2010-12-13|2010-12-16|Complete|Done|4|3|4|3|4|4|3.67|||||||||2|3|4|3|2|3|2.83|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|4|3|||||2|2|||||||||Green||Volunteer: Time constraint|8.3||1|1|2|2|F|Black||20|No|GrandMother|28025|Grandparents|Unknown||Yes|Brochure|Media|General Community||Match Support|F|Black||35|28083|Bachelors Degree|Single|Customer Service||5|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500002335|501860746|31|0|2|502078407|31|0|2|500505055|2||-2||4|1|||-2|500000294|-2|51|1|||7464|9|||1|223006|-1|4|3|44
502280284|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-13|2013-07-31|Followup|2011-12-13|2011-12-14|Complete|Done|1|3|4|4|4|4|3.33|4|3|3|2|4|4|3.33|0|2|4|3|3|2|4|3|3|4|4|2|3|4|3.33|-9.91|4|4|4|4|4|4|4|4|0|5|4|2|3|3.5|3|3|3|3|3|16.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|1|1|100|4|4||||Red|Project Big|Volunteer: Lost contact with child/agency|31.6||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|White||31|28205|Associate Degree|Married|Business: Human Resources||3|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502280719|31|0|2|502241391|1|0|2|500500329|2||500004641||4|3|500004640|500004640|-2|500004640|-2|0|10|||46|2|||1|223211|216597|4|3|45
501729405|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-14|2013-06-16|Followup|2011-12-14|2011-12-06|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|1|2|3|2.5|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|30.1||2|2|1|1|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|RTBM|F|White||33|28204|Bachelors Degree|Single|Business: Sales|28210|0|7|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501729745|31|0|2|502361956|1|0|2|500501689|2||500004772||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|4|||7464|9|||1|223589||4|3|45
500185865|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-15|2014-08-20|Followup|2011-12-15|2012-01-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|68.1||2|2|2|2|F|Black||19||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187761|31|0|2|500189140|31|0|2|500326656|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|223629||4|1|45
501788773|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-27|2012-06-28|Followup|2011-10-27|2011-12-13|Declined|Late||||||||3|2|2|1|4|4|2.67|||||||||2|4|3|4|4|3|3.33||||||4|4|3|3.67|||||||3|4|4|5|4||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||2|2|2||||2|2|||||||Green|Amachi|Volunteer: Moved|32||1|1|1|1|M|Black||18|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|RTBM|M|White||33|28202|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501789128|31|0|1|501845020|1|0|1|500393644|2||-2||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|223672|7735|4|1|45
502138562|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-14|2013-06-06|Followup|2011-12-14|2011-11-06|Complete|Early|2|2|4|4|4|4|3.33|2|3|4|3|1|1|2.33|42.92|3|4|4|1|3|4|3.17|1|2|1|4|4|4|2.67|18.73|4|2|3|3|3|3|3|3|0|5|4|5|4|4.5|5|4|4|5|4.5|0|4|4|4|3|3|4|3|3.57|4|4|4|4|4|4|4|4|-10.75|4|4|4|4|4|4|4|4|0|4|2|3|4|2|3|0|1|1|2|2|-50|4|4||||Green||Child: Lost interest|29.7||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||38|28216|Masters Degree|Single|Finance: Auditor|28217|3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500011746|502138991|31|0|1|502380370|31|0|1|500502780|2||-2||4|1|||-2||-2|0|10|||12183|14|||1|223775|220057|4|3|45
500243491|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-16|2012-05-09|Followup|2011-12-16|2011-12-29|Complete|Done|2|2|4|4|4|4|3.33|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|16.8||4|4|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|F|Black||35|28270||Single|Business: Mgt, Admin||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500013781|500188056|31|0|2|501689965|31|0|2|500505331|2||500003586||4|3|500000294|500000294|-2|500000294, 500004640|-2|0|4|||7496|10|||1|224960||4|3|45
502129650|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-17|2012-09-27|Followup|2011-12-17|2011-12-05|Complete|Done|4|4|4|3|3|4|3.67|4|4|4|4|4|4|4|-8.25|2|3|4|2|4|4|3.17|1|4|3|4|1|4|2.83|12.01|4|4|4|4|4|4|4|4|0|4|5|5|5|4.75|5|4|5|4|4.5|5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4||||Yellow||Volunteer: Lost contact with child/agency|21.4||2|2|1|1|F|Black||17|No|GrandMother|28027|Grandparents|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|Black||29|28027|||Customer Service||0|0||High School Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|502130079|31|0|2|501733783|31|0|2|500502959|2||-2||4|2||500016374|-2||-2|0|10|||0|4|||1|225758|220242|4|3|45
500187090|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-04|2013-08-29|Followup|2011-10-04|2011-09-19|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||3|4|4|4|4|4|3|3.71||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green||Child: Graduated|82.8||2|2|3|3|F|Black||20||Mother|28216|Two Parent|Unknown||No||School|General Community||Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|500188103|31|0|2|500189320|31|0|2|500125754|2||-2||4|1|||-2|500016374|-2|0|4|||7464|9|||1|225971||4|3|45
501390345|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-26|2011-09-02|Followup|2011-02-26|2011-03-21|Complete|Done|4|3|1|1|4|4|2.83|||||||||1|4|2|1|1|4|2.17|||||||||4|4|4|4||||||1|4|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||2|2|4|2.67||||||4|4|4|||||2|2|||||||||Green|Amachi|Volunteer: Moved|30.2||2|2|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||29|28206|Some College|Single|Retail: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011184|501390617|31|0|1|501474303|1|0|1|500342705|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|226036||4|3|45
501390344|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-26|NaT|Followup|2011-02-26|2011-05-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||96.6||1|1|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Single|Tech: Computer/Programmer||0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|501390617|31|0|1|501380163|1|0|1|500342682|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|226061||4|0|45
500186800|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-06|2012-07-25|Followup|2011-10-06|2011-09-19|Complete|Early|4|3|4|4|4|4|3.83|||||||||2|4|4|1|4|4|3.17|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|93.6||1|1|3|3|F|Black||22||Mother|28216|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|500188103|31|0|2|500189320|31|0|2|500037337|2||-2||4|1|||-2|500016374|-2|0|4|||7464|9|||1|226798||4|3|45
500340183|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-18|2013-08-30|Followup|2011-12-18|2012-01-20|Complete|Done|3|3|4|3|3|4|3.33|||||||||2|3|3|3|2|4|2.83|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Yellow||Volunteer: Lost contact with child/agency|44.4||3|3|1|1|M|Black||17|No|Relative: Other|28208|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction||0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|500340317|31|0|1|501933993|1|0|1|500419988|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|226941||4|3|45
500914579|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-16|2014-12-04|Followup|2011-12-16|2012-01-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Severity of challenges|71.6||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|M|White||32|28277|Bachelors Degree|Single|Tech: Engineer|28117|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500914849|31|0|1|501345550|1|0|1|500323102|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|228485||4|1|45
502198485|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-12|2012-10-17|Baseline|2010-12-28|2011-01-12|Complete|Done|3|2|3|2|1|3|2.33|||||||||2|2|3|3|4|4|3|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|21.2||1|1|2|2|M|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||Yes||School|General Community|Amachi|Match Support|M|Black||53|28262|Some College|Married|Business: Clerical||0|0|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500012459|502198914|31|0|1|500188656|31|0|1|500508298|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|228625|-1|4|3|44
500186106|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-18|2015-08-13|Followup|2011-10-18|2011-09-15|Complete|Early|3|1|3|1|3|3|2.33|||||||||2|3|3|3|3|4|3|||||||||4|4||||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|93.8||2|2|1|1|F|Black||20||Mother|28217|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||35|28211|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187698|31|0|2|500778380|1|0|2|500202993|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|228924||4|3|45
502180724|BBBS of Greater Charlotte|Main Office|C|Active|2010-12-30|NaT|Followup|2011-12-30|2011-12-27|Complete|Done|4|4|4|4|4|4|4|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||74.5|Y|2|2|2|2|M|Black||15|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502181148|31|0|1|502391505|31|0|2|500505039|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7438|1|||1|229235||4|3|45
501967613|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2013-02-26|Followup|2011-12-31|2011-12-28|Complete|Done|4|4|4|4|1|4|3.5|4|3|3|3|3|4|3.33|5.11|1|2|3|2|1|3|2|3|4|3|3|3|2|3|-33.33|4|4|4|4|4|3|3|3.33|20.12|2|3|2|4|2.75|3|4|4|3|3.5|-21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4||||Yellow||Volunteer: Time constraint|25.9||1|1|1|1|F|Black||20|No|Mother|28273|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Finance: Accountant|28277|3|5|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500012459|501968011|31|0|2|502311344|1|0|2|500498762|2||-2||4|2|||-2|500000294, 500004640|-2|34|2|||7496|10|||1|229477|148519|4|3|45
502188863|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2013-10-31|Followup|2011-12-31|2012-01-24|Complete|Done|3|2|2|3|3|3|2.67|4|2|3|2|3|3|2.83|-5.65|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|4|5|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|2|3|33.33|2|2|1|1|100|4|4||||Red|Project Big|Volunteer: Moved|34||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|M|Some Other Race||30|28202|Some College|Single|Tech: Support, Writing|28210|0|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502189292|31|0|1|502288935|41|0|1|500498784|2||-2||4|3|500004640|500004640|-2|500004640|-2|0|10|||46|2|||1|229478|191872|4|3|45
502307478|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2012-04-30|Followup|2011-12-31|2012-01-04|Declined|Done||||||||3|2|3|2|3|3|2.67|||||||||2|4|3|2|3|3|2.83||||||4|4|4|4|||||||1|1|1|1|1||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|2|2.5||||2|2|||||||Red|Project Big|Volunteer: Moved|16||1|1|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Enrollment|M|Black||40|28215|Some College|Married|Transport: Driver||3|0|Michael Baisden|Media|Big|General Community||Match Support|277|60|598|500000170|500013709|502307910|31|0|1|502035292|31|0|1|500503967|2||||4|3|500004640|500004640|-2||-2|0|4|||11146|1|||1|229483|195055|4|1|45
501831581|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-29|NaT|Followup|2011-09-29|2011-09-08|Complete|Early|3|3|1|1|1|3|2|||||||||2|3|4|2|2|4|2.83|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|4|3.67||||||2|2|2|||||2|2||||4|4||||Green|Amachi||89.5||1|1|2|3|F|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||38|28273||Single|Tech: Engineer||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501831944|31|0|2|500715453|31|0|2|500387624|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|229998||4|3|45
501176569|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-08|2012-02-29|Followup|2012-01-08|2012-01-23|Complete|Done|4|2|4|2|4|4|3.33|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green||Child/Family: Moved|37.7||1|1|1|1|M|Multi-race (Black & White)||18||Mother|28031|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28078|Bachelors Degree|Living w/ Significant Other|Education: Admin|28035|2|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501176843|36|0|1|501457533|1|0|1|500327489|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|230071||4|3|45
501516900|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-28|2015-08-27|Followup|2012-01-28|2012-01-26|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|4|4|4|3|4|3.67|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|78.9||1|1|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||39|28212|Bachelors Degree|Single|Medical: Healthcare Worker|28210|1|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500018987|501517192|31|0|2|501438601|31|0|2|500332399|2||-2||4|1|||-2||-2|6854|8|||7462|13|||1|230077||4|3|45
501904094|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-15|2013-06-19|Followup|2012-01-15|2012-01-23|Complete|Done|3|2|4|1|4|3|2.83|4|1|4|2|4|4|3.17|-10.73|3|4|4|3|3|4|3.5|2|4|4|3|4|4|3.5|0|4|4|4|4|4|4|4|4|0|5|4|4|5|4.5|3|4|2|5|3.5|28.57|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|2|3|2.5|4|4|4|-37.5|2|2|2|2|0|4|4||||Red||Volunteer: Lost contact with child/agency|41.1||1|1|1|1|F|Black||16|No|Mother|28214|One Parent: Female|Unknown|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||56|28208|Some College|Single|Finance: Accountant|28203|19|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500004169|501904482|31|0|2|501342148|31|0|2|500420809|2||-2||4|3|||-2|500000294|-2|34|2|||7446|3|||1|230080|23717|4|3|45
501428903|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-21|2015-02-25|Followup|2012-01-21|2012-01-20|Complete|Done|3|4|4|2|3|3|3.17|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|73.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|White||53|15001|Masters Degree|Single|Consultant|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501429188|31|0|1|501441245|1|0|1|500331206|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|230081||4|3|45
501627668|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2012-09-14|Followup|2012-01-26|2012-01-12|Complete|Done|3|1|4|2|4|4|3|||||||||4|3|4|4|2|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Yellow||Volunteer: Moved|31.6||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||38|28209|Bachelors Degree|Single|Business|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|501627988|31|0|1|501865457|1|0|1|500423715|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|230082||4|3|45
501735420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2015-08-13|Followup|2012-01-26|2012-02-13|Complete|Done|3|2|3|3|3|3|2.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green||Child: Lost interest|66.5||2|2|2|2|F|Black||16||GrandMother|28215|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||41|28277|Bachelors Degree|Single|Business: Mgt, Admin||9|0|General|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500017732|501735760|31|0|2|500956022|1|0|2|500428818|2||-2||4|1|||-2||-2|6854|8|||6450|12|||1|230085||4|3|45
502177920|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-14|2012-05-23|Baseline|2011-01-06|2011-01-14|Complete|Done|4|3|4|1|3|4|3.17|||||||||3|4|4|2|4|4|3.5|||||||||3|4|4|3.67||||||4|5|5|2|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2|||||||||Red||Volunteer: Lost contact with child/agency|16.3||1|1|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||59|28212|Associate Degree|Divorced|Transport: Driver|28269|0|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||RTBM|277|60|598|500000170|500011746|502178349|31|0|1|502387867|31|0|1|500509427|2||-2||4|3||500005291|-2||-2|34|2|||12183|14|||1|230935|-1|4|3|44
501744683|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-06|2012-11-28|Followup|2011-11-06|2011-12-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|36.7||1|1|1|1|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||56|28270|Some College|Separated|Unknown|28277|7|7|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500013781|501745023|31|0|1|501863268|31|0|1|500405317|2||-2||4|1|||-2||-2|0|10|||46|2|||1|230948||4|1|45
502365086|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-13|2011-10-25|Baseline|2011-01-06|2011-01-13|Complete|Done|3|4|2|4|3|3|3.17|||||||||3|3|4|4|4|4|3.67|||||||||4|4|3|3.67||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|4|3.33||||||3|2|2.5|||||2|2|||||||||Yellow|Amachi|Child: Lost interest|9.4||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||Yes|TV|Media|General Community|Amachi|Match Support|M|Black||34|28269|Masters Degree|Married|Tech: Research/Design|19355|1|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011184|502365524|31|0|1|502426330|31|0|1|500509521|2||500003586||4|2|500000294|500000294|-2|500000294|-2|56|1|||7446|3|||1|231016|-1|4|3|44
502118927|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-23|2012-05-23|Followup|2011-06-23|2011-09-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|23||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||38|28202||Single|Customer Service||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500008629|502099867|31|0|2|502069043|31|0|2|500455591|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|231113||4|0|45
500496598|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-23|NaT|Followup|2011-10-23|2012-01-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi, Cabarrus County||100.7||2|2|1|1|M|White||15|Yes|Mother|28083|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi, Cabarrus County|Match Support|M|White||35|28083|Masters Degree|Single|Business: Mgt, Admin|28027|2|3|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500496849|1|0|1|501383928|1|0|1|500299090|2||500003586||2|2|500000294, 500016374|500000294, 500016374|-2|500016374|-2|34|2|||7464|9|||1|231179||4|0|45
502312413|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-18|2013-01-03|Baseline|2011-01-07|2011-01-18|Complete|Done|4|2|4|1|1|1|2.17|||||||||2|2|3|4|1|4|2.67|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|4|2.5|||||1|1|||||||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|23.5||1|1|1|1|M|Black||17|Yes|Mother|28211|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||33|28209|Bachelors Degree|Single|Finance: Economist|60602|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011349|502312845|31|0|1|502410938|1|0|1|500509858|2||500003586||4|1|500000294|500000294|-2||-2|7295|11|||7496|10|||1|231459|-1|4|3|44
502312421|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-18|2012-08-29|Baseline|2011-01-12|2011-01-18|Complete|Done|3|3|2|1|1|3|2.17|||||||||4|4|4|1|1|4|3|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1|||||||||Green|Amachi|Volunteer: Moved|19.4||1|1|1|1|M|Black||19|Yes|Mother|28211|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||33|28210|Bachelors Degree|Single|Construction|28269|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502312845|31|0|1|502402041|1|0|1|500510430|2||-2||4|1|500000294|500000294|-2||-2|7295|11|||7496|10|||1|232682|-1|4|3|44
500414909|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-12|2012-07-30|Followup|2012-01-12|2012-03-28|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|2010-2012 OJJDP JJI|Child: Graduated|18.6||3|3|3|3|M|White||22|No|Mother|28027|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||56|28078|Bachelors Degree|Single|Business: Sales|28027|14|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500002335|500415159|1|0|1|500188447|1|0|1|500510533|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7446|3|||1|232791||4|0|45
502198485|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-12|2012-10-17|Followup|2012-01-12|2012-01-03|Complete|Done|4|2|4|1|2|3|2.67|3|2|3|2|1|3|2.33|14.59|3|4|4|3|4|4|3.67|2|2|3|3|4|4|3|22.33|4|4|4|4|4|4|4|4|0|4|4|4|3|3.75|3|4|5|5|4.25|-11.76|2|4|4|4|4|4|4|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|3|3.67|4|4|4|4|-8.25|4|4|4|4|4|4|0|2|2|2|2|0|4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|21.2||1|1|2|2|M|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||Yes||School|General Community|Amachi|Match Support|M|Black||53|28262|Some College|Married|Business: Clerical||0|0|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500012459|502198914|31|0|1|500188656|31|0|1|500508298|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|232809|228625|4|3|45
502443215|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-09|2012-06-30|Baseline|2011-01-12|2011-02-09|Complete|Done|4|2|2|2|3|3|2.67|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|16.7||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black|Other African|50|28215|Bachelors Degree|Divorced|Govt|28208|17|8|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013709|502443662|31|0|2|502348503|31|31|2|500510587|2||-2||4|3|500005291|500005291|-2|500000294|-2|0|10|||7464|9|||1|232852|-1|4|3|44
501853848|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-30|2014-08-29|Followup|2011-11-30|2011-12-20|Complete|Done|4|1|4|1|3|4|2.83|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|56.9||1|1|1|1|M|Black||15|Yes|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|M|Black||33|28273|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501854219|31|0|1|501839466|31|0|1|500405366|2||-2||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|232858||4|3|45
500186260|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-29|2015-12-17|Followup|2011-10-29|2012-01-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|133.6||3|3|1|1|M|Black||19|No|Mother|28025|One Parent: Female|Unknown||No||Self|General Site||Match Support|M|Black||42|28025|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|500187857|31|0|1|500189139|31|0|1|500037139|2||-2||4|2|||-1||-2|0|10|||7464|9|||1|233038||4|0|45
500545326|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2016-09-02|Followup|2011-10-29|2011-12-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|118.1|Y|1|1|1|1|M|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|Black||55|28214||Married|Clergy||12|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|1|500697845|31|0|1|500134545|2||-2||4|3|||-2||-2|0|10|||2238|7|||1|233043||4|1|45
500997812|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-12|2012-11-16|Followup|2012-01-12|2012-03-01|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|46.1||1|1|1|1|M|Black||20|No|Mother|28266|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community||Match Support|M|White||40|28203|Bachelors Degree|Single|Transport: Pilot||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|500998085|31|0|1|501429055|1|0|1|500329285|2||-2||4|1|||-2|500000294|-2|0|10|||7496|10|||1|233391||4|1|45
501686310|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2013-03-13|Followup|2011-10-30|2011-12-13|Declined|Done||||||||3|4|4|4|3|4|3.67|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||4|5|5|5|4.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|4|4||||1|1|||||||Red||Child/Family: Lost contact with volunteer/agency|40.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28211|One Parent: Female|Unknown||No|Radio|Media|General Community||Match Support|M|Black||34|28202|Juris Doctorate (JD)|Single|Law: Lawyer||1|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501686648|36|0|1|501818631|31|0|1|500392214|2||-2||4|3|||-2||-2|55|1|||7446|3|||1|233559|14832|4|1|45
502177920|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-14|2012-05-23|Followup|2012-01-14|2012-02-10|Declined|Done||||||||4|3|4|1|3|4|3.17|||||||||3|4|4|2|4|4|3.5||||||3|4|4|3.67|||||||4|5|5|2|4||||||||||4|4|4|4|3|4|3|3.71||||||4|4|3|3.67|||||3|2|2.5||||2|2|||||||Red||Volunteer: Lost contact with child/agency|16.3||1|1|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||59|28212|Associate Degree|Divorced|Transport: Driver|28269|0|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||RTBM|277|60|598|500000170|500011746|502178349|31|0|1|502387867|31|0|1|500509427|2||-2||4|3||500005291|-2||-2|34|2|||12183|14|||1|233594|230935|4|1|45
502244776|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-19|NaT|Baseline|2011-01-14|2011-01-19|Complete|Done|4|2|2|1|3|4|2.67|||||||||2|3|3|2|3|2|2.5|||||||||4|3|2|3||||||2|3|3|4|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI||73.9||1|1|2|2|F|Black||16|No|Mother|28216|Two Parent|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28209|Bachelors Degree|Single|Law|28273|5|0|Relative|Relative|Big|General Community|Amachi|Match Support|277|60|598|500000170|500021785|502245202|31|0|2|502143351|1|0|2|500511171|2||-2||2|1|500005291|500005291|-2|500000294|-2|0|4|||17161|11|||1|233727|-1|4|3|44
501529924|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2017-02-28|Followup|2011-08-27|2011-08-26|Complete|Done|2|2|2|1|3|2|2|||||||||2|3|2|1|2|2|2|||||||||4|4|4|4||||||2|2|2|2|2|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|78.1||2|2|1|1|F|Black||15|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||30|28209|Bachelors Degree|Single|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501530213|31|0|2|502199360|1|0|2|500465517|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|234032||4|3|45
501261979|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-22|2014-10-13|Followup|2011-07-22|2011-09-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|74.7||1|1|3|3|F|Black||15|No|Mother|28134|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||55|28173||Married|Human Services: Non-Profit|28205|0|0|Coworker|Workplace Partner|Big|General Community|VOL - Maximizing Match Impact|Match Support|277|60|598|500000170|500011349|501262256|31|0|2|500418936|31|0|2|500278634|2||-2||4|1|||-2|500011314|-2|0|10|||7447|3|||1|234112||4|1|45
500897083|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-13|2012-11-19|Followup|2011-11-13|2012-01-03|Declined|Late||||||||4|1|4|1|3|4|2.83|||||||||3|3|3|4|4|4|3.5||||||4|4|4|4|||||||3|3|4|3|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Red|Amachi|Child/Family: Infraction of match rules/agency policies|36.2||1|1|1|1|M|Black||21|Yes|Mother|28269|One Parent: Female|Unknown|Y|No||Service Organization|General Community|Amachi|Match Support|M|White||54|28210||Married|Self-Employed, Entrepreneur||0|0|Holy Comforter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|500897335|31|0|1|501862348|1|0|1|500407273|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|11|||9216|7|||1|234194|268|4|1|45
500186325|BBBS of Greater Charlotte|Main Office|C|Completed|2003-11-19|2012-11-29|Followup|2011-11-19|2012-01-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|108.4||2|2|2|3|M|Black||22||Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28202|Bachelors Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187951|31|0|1|500189265|1|0|1|500047102|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|234195||4|1|45
501356328|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-21|2012-09-06|Followup|2011-11-21|2012-02-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|45.5||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||33|28269|Masters Degree|Single|Finance: Banking|28255|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501356607|31|0|2|501371070|31|0|2|500315101|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|234196||4|0|45
500185729|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-26|2012-09-05|Followup|2011-11-26|2012-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|57.3||2|2|2|2|M|Black||22||Relative: Other|28208|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||35|2109||Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500187496|31|0|1|500188672|1|0|1|500223221|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|234198||4|1|45
502312413|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-18|2013-01-03|Followup|2012-01-18|2012-03-14|Declined|Late||||||||4|2|4|1|1|1|2.17|||||||||2|2|3|4|1|4|2.67||||||4|4|4|4|||||||4|3|5|5|4.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||1|4|2.5||||1|1|||||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|23.5||1|1|1|1|M|Black||17|Yes|Mother|28211|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||33|28209|Bachelors Degree|Single|Finance: Economist|60602|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011349|502312845|31|0|1|502410938|1|0|1|500509858|2||500003586||4|1|500000294|500000294|-2||-2|7295|11|||7496|10|||1|234325|231459|4|1|45
502312421|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-18|2012-08-29|Followup|2012-01-18|2012-03-14|Declined|Late||||||||3|3|2|1|1|3|2.17|||||||||4|4|4|1|1|4|3||||||4|4|4|4|||||||5|4|4|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||1|1|||||||Green|Amachi|Volunteer: Moved|19.4||1|1|1|1|M|Black||19|Yes|Mother|28211|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||33|28210|Bachelors Degree|Single|Construction|28269|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502312845|31|0|1|502402041|1|0|1|500510430|2||-2||4|1|500000294|500000294|-2||-2|7295|11|||7496|10|||1|234331|232682|4|1|45
501313839|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-11|2013-06-18|Followup|2011-11-11|2011-12-23|Declined|Done||||||||3|2|3|3|4|4|3.17|||||||||2|3|4|4|2|4|3.17||||||3|4|4|3.67|||||||4|5|5|5|4.75||||||||||4|4|4|3|2|2|1|2.86||||||3|4|3|3.33|||||3|3|3||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|43.2||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||36|28204|Bachelors Degree|Single|Consultant||4|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501314117|31|0|1|501788563|1|0|1|500396680|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|234464|590|4|1|45
502244776|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-19|NaT|Followup|2012-01-19|2012-01-23|Complete|Done|3|3|4|1|4|4|3.17|4|2|2|1|3|4|2.67|18.73|4|3|4|4|3|4|3.67|2|3|3|2|3|2|2.5|46.8|4|4|4|4|4|3|2|3|33.33|5|3|5|4|4.25|2|3|3|4|3|41.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|2|2|2|2|4|3|-33.33|1|1|2|2|-50|4|4|4|4|0|Green|2010-2012 OJJDP JJI||73.9||1|1|2|2|F|Black||16|No|Mother|28216|Two Parent|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28209|Bachelors Degree|Single|Law|28273|5|0|Relative|Relative|Big|General Community|Amachi|Match Support|277|60|598|500000170|500021785|502245202|31|0|2|502143351|1|0|2|500511171|2||-2||2|1|500005291|500005291|-2|500000294|-2|0|4|||17161|11|||1|234769|233727|4|3|45
502275241|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-21|2015-10-15|Baseline|2011-01-20|2011-03-21|Complete|Done|4|3|3|3|4|3|3.33|||||||||3|3|4|3|3|2|3|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|||||||||||||3|3|3|3||||||3|3|3|||||2|2|||||||||Green|Amachi|Child: Lost interest|54.8||1|1|1|1|F|Black||17|No|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||26|28031|Bachelors Degree|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|502275673|31|0|2|502394690|1|0|2|500521625|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7496|10|||1|235273|-1|4|3|44
502255150|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-14|NaT|Baseline|2011-01-20|2011-02-14|Complete|Done|1|2|1|1|1|4|1.67|||||||||1|4|3|1|1|3|2.17|||||||||4|4|4|4||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||1|1|1|||||2|2|||||||||Green|Amachi||73||1|1|1|1|F|Black||17|Yes|Relative: Other|28227|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||34|28212|Masters Degree|Single|Education: Teacher|28216|6|3|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020752|502255582|31|0|2|502392989|1|0|2|500512287|2||500003586||2|1|500000294|500000294|-2|500000294, 500004640|-2|0|5|||7464|9|||1|235505|-1|4|3|44
500474841|BBBS of Greater Charlotte|Main Office|C|Completed|2006-11-18|2012-01-17|Followup|2011-11-18|2011-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|62||1|1|2|2|F|Black||15||Mother|28208|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Multi-Race (None of the above)||52|28227|Bachelors Degree|Single|Education: Admin||4|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500013709|500474737|31|0|2|500370830|7|0|2|500133665|2||-2||4|2|||-2||-2|34|2|||46|2|||1|235954||4|1|45
501249455|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-03|2012-08-30|Followup|2011-12-03|2011-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|44.9||1|1|1|1|M|Black||22|No|Mother|28269|One Parent: Female|Unknown||Yes|Brochure|Media|General Community||Match Support|M|Black||36|28262|Masters Degree|Single|Finance: Banking||6|6|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|501249731|31|0|1|501488627|31|0|1|500317964|2||-2||4|3|||-2||-2|51|1|||7464|9|||1|235955||4|1|45
501201377|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-31|2016-08-26|Followup|2012-01-31|2012-02-01|Complete|Done|4|2|1|1|1|3|2|||||||||2|2|3|2|2|3|2.33|||||||||3|3|2|2.67||||||1|3|2|4|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2||||4|4||||Red||Child: Graduated|90.8||1|1|1|1|F|Hispanic||18|No|Mother|28212|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community||Match Support|F|Hispanic||65|28269|Masters Degree|Single|Medical: Admin|28262|8|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500017777|501201651|3|0|2|501497622|3|0|2|500331903|2||-2||4|3|||-2||-2|7016|11|||7446|3|||1|236513||4|3|45
501060196|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-26|2015-08-03|Followup|2011-11-26|2012-01-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|92.2||1|1|1|1|M|Black||19|No|Mother|28205|One Parent: Female|$15,000 to $19,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28226|Masters Degree|Single|Finance: Accountant||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501060469|31|0|1|501036081|1|0|1|500223215|2||-2||4|1|||-2||-2|34|2|||46|2|||1|237159||4|1|45
500191327|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-07|2012-09-05|Followup|2011-12-07|2012-01-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Family structure changed|69||2|2|1|1|M|Black||19||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28212||Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008629|500191330|31|0|1|500547393|31|0|1|500144146|2||-2||4|1|||-2||-2|0|10|||46|2|||1|237167||4|1|45
501454635|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-19|2013-09-30|Followup|2012-01-19|2012-01-23|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|44.4||1|1|2|2|M|Black||15|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Some Other Race||40|28216|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|501454920|31|0|1|500188923|41|0|1|500424889|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|238463||4|3|45
501936316|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-28|2016-08-29|Followup|2012-01-28|2012-03-09|Declined|Done||||||||3|3|3|2|2|2|2.5|||||||||3|3||3|3|3|||||||3|3|3|3|||||||4|5|4|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Child/Family: Lost contact with volunteer/agency|79||1|1|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||54|28203|||Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|501936714|31|0|1|501872326|1|0|1|500428557|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|238799|28181|4|1|45
501771263|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-02-28|Followup|2011-09-29|2011-10-03|Complete|Done|3|3|4|3|3|3|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|89||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||31|28262|Bachelors Degree|Single|Medical: Admin|28216|0|8|Recruitment Event|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501741899|31|0|2|501622704|31|0|2|500379993|2||-2||4|1|||-2||-2|0|10|||7443|2|||1|239277||4|3|45
501185592|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-23|2016-03-03|Followup|2011-06-23|2011-07-21|Complete|Done|4|1|4|3|4|4|3.33|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2|||||||||Green||Child: Family structure changed|92.3|Y|1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||45|28211||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501255830|1|0|1|500270254|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|239281||4|3|45
502431042|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-10|2013-12-20|Baseline|2011-02-03|2011-02-10|Complete|Done|3|4|2|3|4|4|3.33|||||||||2|3|3|3|4|3|3|||||||||4|4|4|4||||||3|4|5|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|34.3||1|1|1|1|F|Black||17|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||34|28226|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502431483|31|0|2|502447496|1|0|2|500515174|2||-2||4|2|500005291|500005291|-2||-2|0|10|||7464|9|||1|240749|-1|4|3|44
502211307|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-03|2014-04-24|Followup|2012-02-03|2012-01-27|Complete|Done|4|4|4|2|4|4|3.67|4|4|4|3|4|3|3.67|0|2|3|4|2|2|3|2.67|4|3|3|4|3|3|3.33|-19.82|4|4|4|4|4|4|4|4|0|5|4|4|3|4|4|4|4||||4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4||3|||1|1|2|2|-50|4|4||||Yellow|Amachi|Volunteer: Time constraint|38.6||1|1|1|1|M|Black||16|Yes|Mother|28278|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||51|28214|Bachelors Degree|Single|Business: Sales|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502211737|31|0|1|502371462|1|0|1|500512414|2||-2||4|2|500000294|500000294|-2|500000294|-2|7016|11|||7496|10|||1|240822|177660|4|3|45
502197477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-10|2016-10-03|Baseline|2011-02-04|2011-02-10|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|3|3|4|3|3|3|||||||||3|3|3|3||||||5|3|3|5|4|||||||4|4|4|3|3|4|4|3.71||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Moved|67.7||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28202|Bachelors Degree|Single|Business: Sales|27560|1|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017732|502197915|31|0|1|502422929|1|0|1|500515536|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|4|||7464|9|||1|241218|-1|4|3|44
501860404|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-21|2012-07-31|Followup|2012-01-21|2012-01-23|Complete|Done|4|3|4|4|4|4|3.83|3|1|4|2|4|4|3|27.67|2|3|3|3|3|3|2.83|2|4|2||4|3|||4|4|4|4|4|4|4|4|0|3|4|3|2|3|5|3|2|4|3.5|-14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|3|3.67|4|4|3|3.67|0|3|3|3|4|1|2.5|20|2|2|2|2|0|4|4||||Green||Volunteer: Moved|30.3||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Enrollment|M|White||30|28202||Single|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501860777|31|31|1|501893096|1|0|1|500425993|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|242250|26821|4|3|45
500936718|BBBS of Greater Charlotte|Main Office|C|Completed|2007-12-20|2016-06-16|Followup|2011-12-20|2011-12-15|Complete|Done|4|1|4|4|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Agency: Challenges with program/partnership|101.9||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28210|Bachelors Degree|Married|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500017732|500915629|31|0|1|501027885|1|0|1|500224574|2||-2||4|1|||-2|500014505, 500015184|-1|34|2|||46|2|||1|242254||4|3|45
500261295|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-21|2017-03-09|Followup|2011-12-21|2012-01-27|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|2|3|3|3|3|2.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green||Child: Graduated|134.6||1|1|1|1|M|White||20||Mother|28104|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||60|28270|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500261310|1|0|1|500188435|1|0|1|500073081|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|242255||4|3|45
501296349|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-01|2014-02-27|Followup|2011-12-01|2011-12-30|Complete|Done|3|3|3|3|3|3|3|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child: Graduated|62.9||1|1|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||42|28214|Bachelors Degree|Single|Business: Mgt, Admin|28205|3|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501296627|31|0|2|501471640|31|0|2|500318555|2||||4|2|||-2|500000294|-2|0|4|||7464|9|||1|242260||4|3|45
501340105|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2013-06-27|Followup|2011-12-12|2011-12-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Graduated|54.5||1|1|1|1|F|Multi-race (Black & Hispanic)||21|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||53|28269||Married|Medical: Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340376|38|0|2|501514453|1|0|2|500322778|2||-2||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|242308||4|1|45
500733695|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-26|2015-03-03|Followup|2011-12-26|2011-12-29|Complete|Done|4|2|4|4|4|4|3.67|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.2||1|1|1|1|F|Black||19|Yes|GrandMother|28217|Grandparents|Less than $10,000|Y|No|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||34|28210|Bachelors Degree|Married|Finance: Accountant|28202|0|2|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500733962|31|0|2|500307108|1|0|2|500150172|2||500003586||4|3|500000294|500000294|-2||-2|7294|13|||2238|7|||1|242309||4|3|45
501114434|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-23|2014-06-12|Followup|2011-12-23|2011-12-30|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|65.6||1|1|1|1|M|Black||20|No|Uncle|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||33|28207|Masters Degree|Single|Finance: Accountant|28244|0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501114708|31|0|1|501315131|1|0|1|500324423|2||-2||4|3|500000294|500000294|-2||-2|0|10|||130|1|11|3|1|242310||4|3|45
501292079|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-11|2013-07-18|Followup|2011-12-11|2011-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Lost interest|55.2||1|1|1|1|F|Black||17|Yes|GrandMother|28214|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||31|28203|Bachelors Degree|Single|Consultant|28204|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501292357|31|0|2|501519897|1|0|2|500323243|2||500003586||4|1|500000294|500000294|-2||-2|7294|13|||7464|9|||1|242311||4|1|45
500636617|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-10|2013-08-20|Followup|2012-01-10|2012-02-12|Complete|Done|2|4|4|3|4|4|3.5|||||||||4|4|4|1|3|4|3.33|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|79.3||2|2|1|1|M|Black||17||Mother|28269|One Parent: Female|$20,000 to $24,999|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28262||Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500636863|31|0|1|500756919|31|0|1|500151137|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|242415||4|3|45
502443215|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-09|2012-06-30|Followup|2012-02-09|2012-04-25|Expired|Late||||||||4|2|2|2|3|3|2.67|||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||2|3|3|3|2.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|16.7||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black|Other African|50|28215|Bachelors Degree|Divorced|Govt|28208|17|8|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013709|502443662|31|0|2|502348503|31|31|2|500510587|2||-2||4|3|500005291|500005291|-2|500000294|-2|0|10|||7464|9|||1|242665|232852|4|0|45
502197477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-10|2016-10-03|Followup|2012-02-10|2012-01-20|Complete|Early|3|2|2|2|3|3|2.5|4|3|4|4|4|4|3.83|-34.73|2|3|3|3|3|3|2.83|2|3|3|4|3|3|3|-5.67|4|4|4|4|3|3|3|3|33.33|2|2|3|3|2.5|5|3|3|5|4|-37.5|4|4|4|4|4|4|4|4|4|4|4|3|3|4|4|3.71|7.82|4|4|4|4|4|4|3|3.67|8.99|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Moved|67.7||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28202|Bachelors Degree|Single|Business: Sales|27560|1|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017732|502197915|31|0|1|502422929|1|0|1|500515536|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|4|||7464|9|||1|243075|241218|4|3|45
502272172|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-23|2012-06-28|Baseline|2011-02-10|2011-02-23|Complete|Done|3|4|4|1|4|4|3.33|||||||||2|4|2|1|3|3|2.5|||||||||4|4|4|4||||||2|3|3|4|3|||||||4|4|4|4|4|4|4|4||||||||||1|1|1|1||||||4|3|3.5|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Moved|16.1||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||29|28277||Single|Student: College||0|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502272604|31|0|2|502296220|1|0|2|500516654|2||-2||4|3|500005291||-2|500004640|-2|6854|8|||7464|9|||1|243094|-1|4|3|44
502290600|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-18|2012-04-30|Baseline|2011-02-10|2011-02-18|Complete|Done|4|4|4|3|3|4|3.67|||||||||3|4|3|4|4|3|3.5|||||||||4|3|3|3.33||||||4|5|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1|||||||||Yellow|Amachi|Volunteer: Lost contact with child/agency|14.4||1|1|1|1|M|Black||17|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Radio|Media|General Community|Amachi|Enrollment|M|Some Other Race||52|28031|Some College|Married|Govt|28031|17|0|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|502291037|31|0|1|502450688|41|0|1|500516671|2||-2||4|2|500000294|500000294|-2||-2|55|1|||7452|6|||1|243116|-1|4|3|44
502431042|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-10|2013-12-20|Followup|2012-02-10|2012-01-09|Complete|Early|3|3|4|2|4|4|3.33|3|4|2|3|4|4|3.33|0|3|3|4|4|4|4|3.67|2|3|3|3|4|3|3|22.33|4|4|4|4|4|4|4|4|0|4|5|5|4|4.5|3|4|5|3|3.75|20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|1|1|1|1|0|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|34.3||1|1|1|1|F|Black||17|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||34|28226|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502431483|31|0|2|502447496|1|0|2|500515174|2||-2||4|2|500005291|500005291|-2||-2|0|10|||7464|9|||1|243200|240749|4|3|45
500185637|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-29|2014-12-11|Followup|2011-12-29|2011-12-15|Complete|Done|3|2|4|4|3|3|3.17|||||||||3|4|3|3|2|3|3|||||||||4|4||||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|107.4||1|1|2|2|M|Black||20||Mother|28206|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Black||55|28297|Masters Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500187271|31|0|1|500189284|31|0|1|500073080|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|243575||4|3|45
500185601|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-28|2015-07-23|Followup|2012-01-28|2012-01-26|Complete|Done|3|2|4|2|4|4|3.17|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green||Child: Graduated|89.8||2|2|1|1|M|Black||20||Mother|28210|Other/Unknown|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28078|High School Graduate|Single|Finance: Accountant|28202|0|4|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500187235|31|0|1|501082220|1|0|1|500236473|2||-2||4|1|||-2||-2|6854|8|||7458|9|||1|243578||4|3|45
501070152|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-29|2012-04-17|Followup|2011-11-29|2011-12-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|52.6||1|1|2|2|M|Black||20|Yes|Mother|28212|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community|Amachi|Match Support|M|Black||45|28079|Bachelors Degree|Married|Business||13|6|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500001281|501070425|31|0|1|501052547|31|0|1|500224306|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||7671|13|||1|243579||4|1|45
501045214|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-30|2015-12-16|Followup|2011-11-30|2012-02-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|96.5||1|1|2|2|F|Black||20|No|Relative: Other|28269|Grandparents|$20,000 to $24,999||Yes||BBBS Board/Staff|General Community||Match Support|F|Black||35|28213|Masters Degree|Single|Business||4|0|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|277|60|598|500000170|500002335|501045484|31|0|2|500953330|31|0|2|500217682|2||-2||4|1|||-2|500014505, 500016394|-1|0|13|||46|2|||1|243980||4|0|45
502255150|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-14|NaT|Followup|2012-02-14|2012-04-30|Expired|Late||||||||1|2|1|1|1|4|1.67|||||||||1|4|3|1|1|3|2.17||||||4|4|4|4|||||||2|3|3|2|2.5||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||1|1|1||||2|2|||||||Green|Amachi||73||1|1|1|1|F|Black||17|Yes|Relative: Other|28227|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||34|28212|Masters Degree|Single|Education: Teacher|28216|6|3|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020752|502255582|31|0|2|502392989|1|0|2|500512287|2||500003586||2|1|500000294|500000294|-2|500000294, 500004640|-2|0|5|||7464|9|||1|244181|235505|4|0|45
502136043|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-21|2013-06-06|Baseline|2011-02-14|2011-02-21|Complete|Done|4|1|4|4|3|4|3.33|||||||||3|4|2|1|3|3|2.67|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|3|4|3.86||||||||||4|4|3|3.67||||||3|4|3.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Moved|27.5||1|1|2|2|M|Black||19|No|GrandMother|28227|Other Relative|Unknown||Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502136472|31|0|1|502459922|1|0|1|500517447|2||-2||4|1|500005291|500005291|-2|500004640|-2|56|1|||7464|9|||1|244354|-1|4|3|44
502421176|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-10|2013-03-21|Baseline|2011-02-14|2011-03-10|Complete|Done|3|3|3|2|3|2|2.67|||||||||2|2|4|2|4|4|3|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|24.4||2|2|1|1|F|Black||18|No|GrandMother|28214|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||33|28273|Bachelors Degree|Single|Insurance||0|0|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500004169|502421614|31|0|2|502419727|31|0|2|500517478|2||-2||4|3|500005291||-2|500000294, 500004640|-2|0|4|||46|2|||1|244394|-1|4|3|44
501185594|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-29|2016-06-15|Followup|2012-03-01|2012-02-21|Complete|Done|4|3|4|3|3|3|3.33|||||||||2|3|4|2|2|4|2.83|||||||||4|4|4|4||||||3|2|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|99.5||1|1|1|1|M|Multi-race (Black & White)||19|No|Mother|28227|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Consultant|28226|0|8|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501153366|1|0|1|500248756|2||-2||4|1|||-2||-2|0|4|||7452|6|||1|245056||4|3|45
500185897|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-05|2014-01-31|Followup|2012-02-05|2012-02-02|Complete|Done|2|4|4|4|4|4|3.67|||||||||1|1|4|4|4|3|2.83|||||||||3|4|4|3.67||||||2|3|4|4|3.25|||||||4|4|4|4|3|4|4|3.86||||||||||3|3|1|2.33||||||3|4|3.5|||||2|2||||4|4||||Red|Project Big|Child: Graduated|83.8||2|2|1|1|M|Black||21|No|Relative: Other|28208|Other Relative|Unknown||No||Self|General Community||Match Support|M|White||39|28277|Bachelors Degree|Single|Tech: Computer/Programmer||4|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500008321|500187458|31|0|1|500549520|1|0|1|500155451|2||500004641||4|3|500004640||-2||-2|0|10|||46|2|||1|245259||4|3|45
502472483|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2014-08-28|Baseline|2011-02-16|2011-02-28|Complete|Done|3|1|4|4|1|1|2.33|||||||||2|2|3|3|4|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|3|2.5|||||1|1|||||||||Red|Amachi|Volunteer: Time constraint|42||1|1|1|1|F|Black||18|Yes|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi|Match Support|F|White||33|28202|Bachelors Degree|Single|Education|28208|4|10|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013781|502472930|31|0|2|502453698|1|0|2|500518061|2||500003586||4|3|500000294|500000294|-2|500004640|-2|0|10|||7464|9|||1|245268|-1|4|3|44
500796255|BBBS of Greater Charlotte|Main Office|C|Active|2010-01-20|NaT|Followup|2012-01-20|2012-01-26|Complete|Done|4|2|2|2|4|4|3|||||||||2|4|4|3|3|3|3.17|||||||||4|4|3|3.67||||||3|3|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|4|3.5|||||2|2||||4|4||||Green|||85.8||3|3|1|1|M|White||18|No|Mother|28031|One Parent: Male|$20,000 to $24,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||60|28269|||Medical: Admin|28207|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500796529|1|0|1|501846438|1|0|1|500424314|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|245286||4|3|45
502378719|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-24|2012-06-29|Baseline|2011-02-16|2011-02-24|Complete|Done|4|3|4|1|4|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|3|3|3.33||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|16.1||1|1|1|1|F|Black||15|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|F|White||30|28202|Bachelors Degree|Single|Business: Marketing||1|0|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500001281|502379157|31|0|2|502454212|1|0|2|500518127|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|10|||46|2|||1|245362|-1|4|3|44
502316483|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-25|2012-09-27|Baseline|2011-02-17|2011-02-25|Complete|Done|4|2|4|4|3|4|3.5|||||||||2|3|3|3|4|1|2.67|||||||||3|3|2|2.67||||||3|2|3|2|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|4|3.67||||||4|4|4|||||1|1|||||||||Yellow|Project Big AND Amachi|Child: Lost interest|19.1||1|1|1|1|M|Black||19|Yes|Mother|28208|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|M|Black||32|28269|Bachelors Degree|Single|Medical: Pharmacist|27511|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|501467438|31|0|1|502428948|31|0|1|500518256|2||500003586||4|2|500004901|500000294|-2|500000294|-2|0|4|||7496|10|||1|245665|-1|4|3|44
502290600|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-18|2012-04-30|Followup|2012-02-18|2012-01-27|Complete|Early|4|2|4|1|4|4|3.17|4|4|4|3|3|4|3.67|-13.62|2|4|4|4|2|4|3.33|3|4|3|4|4|3|3.5|-4.86|4|4|4|4|4|3|3|3.33|20.12|3|5|5|2|3.75|4|5|3|3|3.75|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|3|3.67|8.99|4|2|3|4|4|4|-25|1|1|1|1|0|4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|14.4||1|1|1|1|M|Black||17|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Radio|Media|General Community|Amachi|Enrollment|M|Some Other Race||52|28031|Some College|Married|Govt|28031|17|0|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|502291037|31|0|1|502450688|41|0|1|500516671|2||-2||4|2|500000294|500000294|-2||-2|55|1|||7452|6|||1|246061|243116|4|3|45
502291098|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-03|2011-10-25|Baseline|2011-02-18|2011-03-03|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|4|4|4|4|3|3.67|||||||||4|4|4|4||||||3|4|2|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|7.8||2|2|4|4|F|Black||20|No|Mother|28203|One Parent: Female|Unknown||Yes|Brochure|Media|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||38|28219||Single|Finance: Banking|28273|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011184|502291530|31|0|2|500459674|31|0|2|500518681|2||-2||4|2|500005291|500005291|-2|500000294|-2|51|1|||2238|7|||1|246279|-1|4|3|44
502136043|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-21|2013-06-06|Followup|2012-02-21|2012-02-16|Complete|Done|3|3|4|3|4|3|3.33|4|1|4|4|3|4|3.33|0|3|4|3|2|2|3|2.83|3|4|2|1|3|3|2.67|5.99|4|4|4|4|4|4|4|4|0|2|4|3|3|3|3|5|5|4|4.25|-29.41|4|4|4|4|4|3|4|3.86|4|4|4|4|4|3|4|3.86|0|4|4|4|4|4|4|3|3.67|8.99|2|4|3|3|4|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Moved|27.5||1|1|2|2|M|Black||19|No|GrandMother|28227|Other Relative|Unknown||Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502136472|31|0|1|502459922|1|0|1|500517447|2||-2||4|1|500005291|500005291|-2|500004640|-2|56|1|||7464|9|||1|246927|244354|4|3|45
501247269|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-21|NaT|Followup|2012-02-21|2012-04-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|2010-2012 OJJDP JJI, Cabarrus County||72.8||2|2|1|1|F|White||15|No|Father|28025|One Parent: Male|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|White||43|28027|Associate Degree|Married|Student: College||4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500341682|1|0|2|501914025|1|0|2|500515263|2||500016307||2|1|500005291, 500016374|500016374|-2|500016374|-2|0|10|||7496|10|||1|246967||4|1|45
501526664|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-25|2013-02-19|Followup|2011-02-25|2011-05-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Moved|47.8||1|1|1|1|F|White||15|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|F|White||35|28269|Bachelors Degree|Single|Business: Sales|33609|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|501526956|1|0|2|501233757|1|0|2|500332719|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7496|10|||1|247011||4|0|45
500918264|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-13|2012-02-28|Followup|2012-02-13|2012-02-13|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Severity of challenges|48.5||1|1|1|1|M|Multi-Race (None of the above)||16|No|Mother|28227|Two Mothers|$45,000 to $49,999||No||Self|General Community||Match Support|M|Black||33|28269|Some College|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500001281|500918534|7|0|1|501074231|31|0|1|500236477|2||-2||4|2|||-2||-2|0|10|||46|2|||1|247181||4|1|45
502495214|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2012-03-29|Baseline|2011-02-23|2011-02-28|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|3|2|4|3|3|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Time constraint|13||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||61|28056||Married|Medical: Pharmacist||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|502495663|31|0|2|502346954|31|0|2|500519656|2||500004772||4|2|500000294, 500004640, 500004901, 500005291|500004640, 500005291|-2||-2|0|4|459|3|10326|3|||1|248006|-1|4|3|44
502272172|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-23|2012-06-28|Followup|2012-02-23|2012-03-01|Complete|Done|3|2|3|2|4|4|3|3|4|4|1|4|4|3.33|-9.91|2|4|4|2|2|4|3|2|4|2|1|3|3|2.5|20|4|4|4|4|4|4|4|4|0|1|5|5|5|4|2|3|3|4|3|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|1|1|1|1|267|2|4|3|4|3|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Moved|16.1||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||29|28277||Single|Student: College||0|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502272604|31|0|2|502296220|1|0|2|500516654|2||-2||4|3|500005291||-2|500004640|-2|6854|8|||7464|9|||1|248067|243094|4|3|45
502378719|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-24|2012-06-29|Followup|2012-02-24|2012-03-08|Complete|Done|4|1|4|4|3|4|3.33|4|3|4|1|4|4|3.33|0|2|3|4|4|4|3|3.33|4|4|4|4|4|4|4|-16.75|4|4|4|4|4|3|3|3.33|20.12|4|4|5|5|4.5|4|5|4|5|4.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|2|4|3|0|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|16.1||1|1|1|1|F|Black||15|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|F|White||30|28202|Bachelors Degree|Single|Business: Marketing||1|0|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500001281|502379157|31|0|2|502454212|1|0|2|500518127|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|10|||46|2|||1|248427|245362|4|3|45
502462646|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-18|2013-02-28|Baseline|2011-02-24|2011-03-18|Complete|Done|3|3|3|2|4|4|3.17|||||||||3|4|4|2|2|4|3.17|||||||||4|4|4|4||||||4|5|3|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Child: Lost interest|23.4||1|1|1|1|F|Black||19|No|Mother|28262|One Parent: Female|$25,000 to $29,999||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||36|28269|PHD|Living w/ Significant Other|Medical: Pharmacist|28217|4|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|502463093|31|0|2|502431913|31|0|2|500520035|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|248602|-1|4|3|44
501536733|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-26|2017-02-06|Followup|2011-11-26|2012-02-07|Complete|Late|2|1|2|1|1|2|1.5|||||||||1|3|2|2|2|3|2.17|||||||||4|4|4|4||||||1|4|5|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Red|Cabarrus County|Child: Severity of challenges|98.4||3|3|1|1|F|White||15||Father|28025|One Parent: Male|Unknown||No||School|General Site|Cabarrus County|Match Support|F|White||44|28037|Bachelors Degree|Married|Business: Sales|28027|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501537025|1|0|2|501418563|1|0|2|500320917|2||500016307||4|3|500016374|500016374|-1|500016374|-2|0|4|||7464|9|||1|248763||4|3|45
502316483|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-25|2012-09-27|Followup|2012-02-25|2012-03-08|Complete|Done|3|2|2|2|3|3|2.5|4|2|4|4|3|4|3.5|-28.57|2|3|2|2|4|3|2.67|2|3|3|3|4|1|2.67|0|4|4|4|4|3|3|2|2.67|49.81|3|3|4|3|3.25|3|2|3|2|2.5|30|3|4|4|4|4|4|4|3.86|4|4|4|4|4|4|3|3.86|0|3|3|3|3|4|3|4|3.67|-18.26|2|3|2.5|4|4|4|-37.5|2|2|1|1|100|3|3||||Yellow|Project Big AND Amachi|Child: Lost interest|19.1||1|1|1|1|M|Black||19|Yes|Mother|28208|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|M|Black||32|28269|Bachelors Degree|Single|Medical: Pharmacist|27511|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|501467438|31|0|1|502428948|31|0|1|500518256|2||500003586||4|2|500004901|500000294|-2|500000294|-2|0|4|||7496|10|||1|248881|245665|4|3|45
500961274|BBBS of Greater Charlotte|Main Office|C|Active|2007-08-27|NaT|Followup|2011-08-27|2011-09-07|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||114.6||1|1|2|2|F|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28216|Bachelors Degree|Divorced|Business: Clerical|28204|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500934638|31|0|2|500403000|31|0|2|500186952|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|249281||4|3|45
500186071|BBBS of Greater Charlotte|Main Office|C|Completed|2004-01-05|2014-04-30|Followup|2012-01-05|2012-02-09|Complete|Done|4|2|4|3|3|3|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green||Child: Graduated|123.8||1|1|1|1|M|White||21|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||40|28277|Masters Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187670|1|0|1|500189012|1|0|1|500037012|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|249730||4|3|45
500186327|BBBS of Greater Charlotte|Main Office|C|Completed|2003-01-11|2012-11-30|Followup|2012-01-11|2012-03-27|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|118.6||1|1|1|1|M|Black||22||Mother|28208|One Parent: Female|Unknown|Y|No||School|General Community||Match Support|M|White||63|28211|Some College|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|500187974|31|0|1|500189289|1|0|1|500037301|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|249732||4|0|45
501833031|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2015-11-04|Followup|2012-02-28|2012-03-14|Complete|Done|3|4|2|1|4|4|3|3|3|1|4|4|4|3.17|-5.36|2|4|4|1|2|3|2.67|2|2|3|2|4|4|2.83|-5.65|4|4|4|4|4|4|4|4|0|4|5|4|5|4.5|4|4|4|4|4|12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|4|4|4|4|-8.25|4|4|4|4|2|3|33.33|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Moved|56.2||1|1|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28205|Masters Degree|Single|Medical: Doctor, Provider|28277|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502427342|1|0|2|500518294|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|249812|157600|4|3|45
502495214|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2012-03-29|Followup|2012-02-28|2012-02-20|Complete|Done|4|4|4|4|3|4|3.83|4|4|4|4|4|4|4|-4.25|2|4|3|2|4|4|3.17|2|4|3|2|4|3|3|5.67|4|4|4|4|4|4|4|4|0|4|3|4|4|3.75|3|4|5|5|4.25|-11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Time constraint|13||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||61|28056||Married|Medical: Pharmacist||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|502495663|31|0|2|502346954|31|0|2|500519656|2||500004772||4|2|500000294, 500004640, 500004901, 500005291|500004640, 500005291|-2||-2|0|4|459|3|10326|3|||1|250135|248006|4|3|45
502472483|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2014-08-28|Followup|2012-02-28|2012-02-13|Complete|Done|3|2|4|4|1|1|2.5|3|1|4|4|1|1|2.33|7.3|2|2|3|3|4|3|2.83|2|2|3|3|4|3|2.83|0|4|4|4|4|4|4|4|4|0|2|4|4|3|3.25|3|3|3|3|3|8.33|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|3|4|4|3.67|4|4|4|4|-8.25|4|4|4|2|3|2.5|60|2|2|1|1|100|4|4||||Red|Amachi|Volunteer: Time constraint|42||1|1|1|1|F|Black||18|Yes|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi|Match Support|F|White||33|28202|Bachelors Degree|Single|Education|28208|4|10|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013781|502472930|31|0|2|502453698|1|0|2|500518061|2||500003586||4|3|500000294|500000294|-2|500004640|-2|0|10|||7464|9|||1|250273|245268|4|3|45
502057399|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2014-03-31|Followup|2012-02-28|2012-02-29|Complete|Done|3|2|2|2|3|3|2.5|4|3|4|3|2|4|3.33|-24.92|2|4|4|1|3|3|2.83|3|3|2|3|3|3|2.83|0|4|4|4|4|4|4|4|4|0|4|3|3|4|3.5|4|5|5|4|4.5|-22.22|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|4|1|2.5|60|2|2|2|2|0|4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|37||2|2|1|1|M|White||20|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||50|28078|Bachelors Degree|Single|Arts, Entertainment, Sports|28078|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502057823|1|0|1|502389976|1|0|1|500516780|2||-2||4|2|500005291|500005291|-2||-2|0|4|||7464|9|||1|250292|161076|4|3|45
502233625|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-02|2012-06-29|Followup|2012-03-02|2012-03-03|Complete|Done|3|1|3|1|4|4|2.67|3|3|3|2|1|3|2.5|6.8|2|3|4|4|4|4|3.5|2|3|3|3|4|3|3|16.67|4|4|4|4|4|4|4|4|0|4|5|4|5|4.5|3|5|4|4|4|12.5|4|3|4|4|4|4|4|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|4|3|4|4|4|-25|2|2|2|2|0|4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Moved|15.9||3|3|1|1|F|Multi-race (Hispanic & White)||17|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||29|28262|Bachelors Degree|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502234056|35|0|2|502381327|1|0|2|500519189|2||-2||4|2|500005291||-2||-2|0|10|||7464|9|||1|250961|168274|4|3|45
501833026|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-02|2016-09-30|Followup|2012-03-02|2012-02-29|Complete|Done|4|4|4|4|3|4|3.83|2|4|4|3|1|3|2.83|35.34|2|4|4|2|2|3|2.83|2|1|3|2|3|2|2.17|30.41|4|4|4|4|4|4|4|4|0|3|4|2|3|3|3|4|3|3|3.25|-7.69|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|2|3|33.33|4|4|4|2|4|3|33.33|2|2|1|1|100|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|67||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28205|Masters Degree|Single|Education: Teacher|2122|1|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502451325|1|0|2|500518305|2||-2||4|2|500005291|500005291|-2|500000294|-2|0|10|||7464|9|||1|250987|157601|4|3|45
501525308|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-16|2015-06-18|Followup|2012-02-16|2012-02-23|Complete|Done|4|4|4|2|1|4|3.17|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|76||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28205|Some College|Married|Retail: Sales|28206|1|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|501525600|31|0|1|501536144|1|0|1|500335230|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|251041||4|3|45
502307585|BBBS of Greater Charlotte|Main Office|C|Active|2011-03-21|NaT|Baseline|2011-03-02|2011-03-21|Complete|Done|4|1|2|1|1|1|1.67|||||||||2|2|4|1|2|3|2.33|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Amachi, Project Big, Project Big AND Amachi||71.9||1|1|1|1|F|Black||17|Yes|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||53|28031||Divorced|Medical: Admin|28207|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500020910|502308017|31|0|2|501519450|1|0|2|500521250|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|4|||7446|3|||1|251051|-1|4|3|44
501989028|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-16|2012-03-27|Baseline|2011-03-04|2011-03-16|Complete|Done|4|1|4|1|4|4|3|||||||||2|3|4|3|4|4|3.33|||||||||4|3|4|3.67||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|12.4||2|2|1|1|M|Black||15|No|Mother|28273|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black|Other African|44|28212|Bachelors Degree|Married|Business: Marketing||12|0|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|502425720|31|0|1|502346780|31|31|1|500521737|2||-2||4|3|500005291|500005291|-2|500000294|-2|6855|8|||7671|13|||1|251884|-1|4|3|44
501378357|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-13|NaT|Followup|2012-02-13|2012-02-20|Complete|Done|1|4|4|4|3|4|3.33|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||97||1|1|2|2|M|Multi-race (Black & White)||18|No|Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Mgt, Admin|28215|10|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501378636|36|0|1|501174997|31|0|1|500339619|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|251953||4|3|45
502183217|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-05|NaT|Followup|2011-08-05|2011-07-19|Complete|Early|1|4|4|4|4|1|3|||||||||4|4|4|2|3|4|3.5|||||||||4|4|4|4||||||4|2|3|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|1|1.5|||||2|2|||||||||Green|Amachi||79.3||1|1|2|2|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|Black||50|28078|||Service: Restaurant|28082|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502183646|31|0|1|501733851|31|0|1|500462588|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|253562||4|3|45
502137968|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-08|2013-01-08|Followup|2012-02-29|2012-04-16|Declined|Late||||||||3|4|3|1|3|4|3|||||||||3|3|4|3|2|4|3.17||||||4|4|4|4|||||||4|5|5|4|4.5||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||4|4|4||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|22.1||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||41|28078|Bachelors Degree|Married|Govt|28262|7|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500011746|502138397|31|0|1|502417993|1|0|1|500521032|2||-2||4|3|500005291|500005291|-2|500000294, 500004640|-2|34|2|||7464|9|||1|254289|159363|4|1|45
502419933|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-28|2011-10-25|Baseline|2011-03-08|2011-03-28|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|3|3|2|3|4|3|||||||||4|4|4|4||||||4|4|4|4|4||||||||4|4|4|4|4|4|||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|6.9||2|2|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$40,000 to $44,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||59|28204|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011184|502371107|31|0|1|502442556|1|0|1|500523858|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|254462|-1|4|3|44
502393980|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-30|2012-04-30|Baseline|2011-03-08|2011-09-29|Complete|Done|3|1|1|1|3|3|2|||||||||2|3|2|2|2|3|2.33|||||||||4|4|4|4||||||2|3|5|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||1|4|1|2||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|7||2|2|1|1|F|Multi-race (Black & White)||16|Yes|Aunt|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||31|28078|Some College|Married|Medical: Healthcare Worker|28262|0|6|Big Champions|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|502394418|36|0|2|502454075|31|0|2|500554127|2||-2||4|1|500000294|500005291|-2||-2|0|5|||7461|12|||1|254548|-1|4|3|44
502230729|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-09|2012-08-27|Followup|2012-03-09|2012-03-20|Complete|Done|4|4|4|4|4|4|4|4|2|3|2|3|4|3|33.33|2|3|3|2|3|2|2.5|2|4|3|3|3|3|3|-16.67|3|2|2|2.33|3|3|2|2.67|-12.73|1|1|1|1|1|2|3|3|3|2.75|-63.64|4|4|4|4|3|3|4|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|4|4|4|4|4|4|0|2|3|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Volunteer: Moved|17.6||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||36|28277|Bachelors Degree|Single|Student: College|28205|0|4|Recruitment Event|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|277|60|598|500000170|500012459|502231160|1|0|1|502483362|1|0|1|500518850|2||-2||4|2|500005291|500005291|-2|500000294, 500005291|-2|34|2|||7459|10|||1|254870|181484|4|3|45
502421671|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2011-05-13|Baseline|2011-03-09|2011-03-31|Complete|Done|3|3|2|2|2|3|2.5|||||||||3|4|4|2|3|3|3.17|||||||||3|3|3|3||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|1.4||1|1|1|1|F|Hispanic|Other Central American|16|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||31|28202|Some College|Single|Business: Marketing||3|0|Self|Self|Big|General Community|Project Big|Enrollment|277|60|598|500000170|500010765|502422110|3|14|2|502272620|1|0|2|500524198|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||7464|9|||1|254952|-1|4|3|44
502495123|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2013-01-08|Baseline|2011-03-09|2011-03-31|Complete|Done|3|4|4|2|1|4|3|||||||||2|4|4|4|4|4|3.67|||||||||4|3|4|3.67||||||5|3|3|4|3.75|||||||4|4|4|4|4|||||||||||||4|4|4|4||||||||||||||||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|21.3||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28207|Bachelors Degree|Single|Finance: Economist|28255|5|0||Relative|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502495572|31|0|2|502473441|1|0|2|500524205|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||0|11|||1|254961|-1|4|3|44
502421176|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-10|2013-03-21|Followup|2012-03-10|2012-04-20|Blank|Done||||||||3|3|3|2|3|2|2.67|||||||||2|2|4|2|4|4|3||||||4|4|4|4|||||||4|5|5|5|4.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|4|4||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|24.4||2|2|1|1|F|Black||18|No|GrandMother|28214|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||33|28273|Bachelors Degree|Single|Insurance||0|0|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500004169|502421614|31|0|2|502419727|31|0|2|500517478|2||-2||4|3|500005291||-2|500000294, 500004640|-2|0|4|||46|2|||1|255236|244394|4|3|45
502030263|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2012-03-31|2012-04-02|Complete|Done|3|4|4|4|3|3|3.5|||||||||3|3|1|4|2|3|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|4|3.67||||||2|4|3|||||2|2||||4|4||||Green|||83.5||1|1|1|1|M|White||15|No|Mother|29710|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community||Match Support|M|White||38|28210|||Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502030662|1|0|1|501923553|1|0|1|500438867|2||-2||2|1|||-2||-2|6855|8|||7464|9|||1|255433||4|3|45
500392419|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-06|2013-08-29|Followup|2012-03-06|2012-04-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Moved|77.8||2|2|1|1|F|Black||21||Father|28105|One Parent: Male|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||32|28277||Single|Business: Sales||0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500392669|31|0|2|500746900|1|0|2|500162012|2||-2||4|2|||-2||-2|6855|8|||7464|9|||1|255590||4|1|45
500765381|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-26|2015-10-20|Followup|2012-02-26|2012-04-20|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|79.7||1|1|1|1|M|Black||16|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|10019|Bachelors Degree|Single|Business: Marketing|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500739190|31|0|1|501579025|1|0|1|500342803|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|255760||4|1|45
501575257|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-18|2013-09-24|Followup|2012-03-18|2012-05-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|54.2||1|1|1|1|M|Black||15|No|Mother|28079|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||38|28079||Married|Law: Police Officer|28211|5|0|Recruitment Event|Self|Big|General Community||Enrollment|277|60|598|500000170|500004169|501575553|31|0|1|501234758|1|0|1|500348757|2||-2||4|3|||-2||-2|0|10|||7458|9|||1|255768||4|1|45
501015962|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-12|2012-05-31|Followup|2012-02-12|2012-01-25|Complete|Early|3|2|4|1|3|2|2.5|||||||||1|2|2|4|2|1|2|||||||||3|3|4|3.33||||||3|2|3|3|2.75|||||||4|4|4|3|3|4|3|3.57||||||||||2|2|2|2||||||3|2|2.5|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Time constraint|51.6||1|1|1|1|F|Black||18|Yes|GrandMother|28208|One Parent: Female|Less than $10,000||Yes||Self|General Community|Amachi|Enrollment|F|White||33|28202|Bachelors Degree|Single|Education: Teacher|28025|1|4|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|501065096|1|0|2|500241396|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||2238|7|||1|255999||4|3|45
502426852|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-22|2012-03-29|Baseline|2011-03-14|2011-03-22|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|2|3|2|3|3|2.67|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4||3|||||||3|3|3|||||2|2|||||||||Yellow||Child/Family: Time constraints|12.3||1|1|1|1|F|Black||19|No|Mother|28278|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||61|28215|Bachelors Degree|Divorced|Self-Employed, Entrepreneur||0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500012459|502427295|31|0|2|502437756|31|0|2|500525086|2||-2||4|2||500000294|-2||-2|0|10|||130|1|||1|256292|-1|4|3|44
501522348|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-17|2013-02-28|Followup|2012-03-17|2012-03-14|Complete|Done|3|4|3|3|4|3|3.33|||||||||3|3|4|2|3|4|3.17|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|3|4|4|4|4|4|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|47.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28031|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Single|Retail: Sales|28117|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|501522640|36|0|1|501223351|1|0|1|500349995|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|256392||4|3|45
500186206|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-24|2013-09-30|Followup|2012-02-24|2012-03-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Moved|103.2||1|1|1|1|M|Black||20||GrandMother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||44|28214|PHD|Married|Medical: Doctor, Provider||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187812|31|0|1|500189157|31|0|1|500037157|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|256724||4|1|45
500796261|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-15|2013-01-31|Followup|2012-03-15|2012-05-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|22.6||4|4|1|1|M|White||15|No|Mother|28031|One Parent: Female|$20,000 to $24,999|Y|No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||36|28078|Bachelors Degree|Single|Real Estate: Realtor|28269|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500796529|1|0|1|502492476|1|0|1|500523882|2||-2||4|1|500005291|500005291|-2||-2|34|2|||7464|9|||1|256907||4|1|45
501376745|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-01|2016-01-11|Followup|2012-04-01|2012-04-12|Complete|Done|3|4|4|4|3|3|3.5|||||||||2|3|2|2|2|3|2.33|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Time constraint|81.3||1|1|3|4|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28269|||Business: Marketing||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|501377024|31|0|2|500725077|31|0|2|500350905|2||-2||4|1|||-2||-2|6854|8|||46|2|||1|256948||4|3|45
501621811|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-16|2017-03-09|Followup|2012-03-16|2012-05-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Project Big|Child/Family: Lost contact with volunteer/agency|95.8||1|1|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||36|28269||Married|Self-Employed, Entrepreneur|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501622131|31|0|2|501621016|31|0|2|500344465|2||-2||4|2|500004640||-2||-2|0|10|||7464|9|||1|257434||4|1|45
502505252|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-21|2012-09-27|Baseline|2011-03-16|2011-03-21|Complete|Done|4|1|4|1|3|3|2.67|||||||||3|4|3|2|1|3|2.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Moved|18.3||2|2|1|1|F|Black||16|No|Mother|28209|One Parent: Female|Less than $10,000|Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28202|Bachelors Degree|Single|Finance: Accountant|28203|2|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500011746|502505701|31|0|2|502350629|1|0|2|500525884|2||-2||4|2|500005291|500005291|-2|500005291|-2|0|10|||7464|9|||1|257458|-1|4|3|44
501989028|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-16|2012-03-27|Followup|2012-03-16|2012-03-09|Declined|Done||||||||4|1|4|1|4|4|3|||||||||2|3|4|3|4|4|3.33||||||4|3|4|3.67|||||||5|4|4|4|4.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|3|2.5||||2|2||||4|4||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|12.4||2|2|1|1|M|Black||15|No|Mother|28273|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black|Other African|44|28212|Bachelors Degree|Married|Business: Marketing||12|0|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|502425720|31|0|1|502346780|31|31|1|500521737|2||-2||4|3|500005291|500005291|-2|500000294|-2|6855|8|||7671|13|||1|257555|251884|4|1|45
502462646|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-18|2013-02-28|Followup|2012-03-18|2012-05-04|Declined|Late||||||||3|3|3|2|4|4|3.17|||||||||3|4|4|2|2|4|3.17||||||4|4|4|4|||||||4|5|3|3|3.75||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||2|3|2.5||||2|2||||4|4||Red|2010-2012 OJJDP JJI|Child: Lost interest|23.4||1|1|1|1|F|Black||19|No|Mother|28262|One Parent: Female|$25,000 to $29,999||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||36|28269|PHD|Living w/ Significant Other|Medical: Pharmacist|28217|4|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|502463093|31|0|2|502431913|31|0|2|500520035|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|258047|248602|4|1|45
501434147|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2012-03-31|2012-05-10|Declined|Done||||||||3|1|4|3|1|3|2.5|||||||||2|4|4|4|4|4|3.67||||||4|4|4|4|||||||4|5|2|5|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Green|||83.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||26|28215|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501434432|31|0|1|501926474|31|0|1|500441566|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|258060|29966|4|1|45
501560189|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-11|2012-05-25|Followup|2012-03-11|2012-04-20|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|26.5||2|2|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||39|28273||Single|Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501560485|31|0|2|501621478|31|0|2|500439156|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|258061||4|1|45
500186385|BBBS of Greater Charlotte|Main Office|C|Completed|2003-02-11|2013-01-09|Followup|2012-02-11|2012-03-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|118.9||1|1|1|1|M|Black||22||Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||43|28269|Bachelors Degree|Single|Finance: Accountant|28262|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|500187967|31|0|1|500189269|31|0|1|500037278|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|258070||4|1|45
501506214|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-28|2016-06-23|Followup|2012-03-28|2012-05-11|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|4|5|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|86.9||1|1|1|1|M|Black||19|No|Mother|28105|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||55|28173|||Unknown|28203|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501506506|31|0|1|501588885|31|0|1|500351462|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|258114||4|3|45
500185863|BBBS of Greater Charlotte|Main Office|C|Completed|2005-03-12|2014-05-15|Followup|2012-03-12|2012-03-30|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|110.1||1|1|1|1|F|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||43|28202|Bachelors Degree|Married|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187435|31|0|2|500188915|1|0|2|500036915|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|258116||4|3|45
501626218|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-24|2014-12-18|Followup|2012-03-24|2012-05-14|Complete|Late|3|4|4|4|3|3|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|68.8||1|1|1|1|F|Black||20|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||30|11215|Bachelors Degree|Single|Consultant|11215|0|5|other|College Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501622822|31|0|2|501587214|31|0|2|500350222|2||-2||4|1|||-2|500000294|-2|0|10|||7670|5|||1|258117||4|3|45
501626199|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-26|2013-09-30|Followup|2012-03-26|2012-05-14|Complete|Late|4|3|2|2|3|3|2.83|||||||||2|3|3|4|2|4|3|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|54.2||1|1|1|1|F|Black||21|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||33|28203|Masters Degree|Single|Finance: Accountant|28211|1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|501622822|31|0|2|501293622|1|0|2|500351814|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|258125||4|3|45
501599416|BBBS of Greater Charlotte|Main Office|C|Active|2009-04-28|NaT|Followup|2011-04-28|2011-06-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||94.6||1|1|1|1|M|White||14|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||46|28078|Masters Degree|Single|Retail: Mgt|28207|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501599736|1|0|1|500188567|1|0|1|500357914|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|258325||4|1|45
500342076|BBBS of Greater Charlotte|Main Office|C|Completed|2006-02-14|2012-02-28|Followup|2012-02-14|2012-02-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|72.4||1|1|1|1|M|Black||23||Mother|28216|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||35|28207|Bachelors Degree|Single|Business: Marketing||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|500342211|31|0|1|500188562|1|0|1|500080816|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|258389||4|1|45
501561529|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-11|2012-08-29|Followup|2011-05-11|2011-06-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|39.6||1|1|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||36|28202|Masters Degree|Single|Business: Sales|28202|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501561821|31|0|1|501333443|1|0|1|500359635|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|258420||4|1|45
502275241|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-21|2015-10-15|Followup|2012-03-21|2012-03-15|Complete|Done|3|3|3|2|3|3|2.83|4|3|3|3|4|3|3.33|-15.02|2|4|3|2|3|3|2.83|3|3|4|3|3|2|3|-5.67|4|4|4|4|4|4|4|4|0|5|4|4|4|4.25|2|3|3|3|2.75|54.55|4|4|4|4|3|4|3|3.71|4|4|4|4|4|||||3|3|2|2.67|3|3|3|3|-11|2|1|1.5|3|3|3|-50|2|2|2|2|0|4|4||||Green|Amachi|Child: Lost interest|54.8||1|1|1|1|F|Black||17|No|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||26|28031|Bachelors Degree|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|502275673|31|0|2|502394690|1|0|2|500521625|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7496|10|||1|258543|235273|4|3|45
502505252|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-21|2012-09-27|Followup|2012-03-21|2012-03-09|Complete|Done|3|4|3|4|3|4|3.5|4|1|4|1|3|3|2.67|31.09|2|3|3|3|2|3|2.67|3|4|3|2|1|3|2.67|0|4|4|4|4|4|4|4|4|0|3|4|4|4|3.75|4|5|4|4|4.25|-11.76|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|3|3.67|4|4|3|3.67|0|4|2|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Volunteer: Moved|18.3||2|2|1|1|F|Black||16|No|Mother|28209|One Parent: Female|Less than $10,000|Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28202|Bachelors Degree|Single|Finance: Accountant|28203|2|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500011746|502505701|31|0|2|502350629|1|0|2|500525884|2||-2||4|2|500005291|500005291|-2|500005291|-2|0|10|||7464|9|||1|258558|257458|4|3|45
502307585|BBBS of Greater Charlotte|Main Office|C|Active|2011-03-21|NaT|Followup|2012-03-21|2012-05-01|Complete|Done|3|2|2|2|2|3|2.33|4|1|2|1|1|1|1.67|39.52|2|4|3|1|2|4|2.67|2|2|4|1|2|3|2.33|14.59|3|4|3|3.33|4|4|4|4|-16.75|5|4|5|4|4.5|4|5|5|5|4.75|-5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|2|2.5|3|3|3|-16.67|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi||71.9||1|1|1|1|F|Black||17|Yes|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||53|28031||Divorced|Medical: Admin|28207|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500020910|502308017|31|0|2|501519450|1|0|2|500521250|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|4|||7446|3|||1|258648|251051|4|3|45
502426852|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-22|2012-03-29|Followup|2012-03-22|2012-03-13|Complete|Done|4|3|3|3|4|4|3.5|4|3|3|3|4|4|3.5|0|3|2|3|2|3|3|2.67|3|2|3|2|3|3|2.67|0|4|4|4|4|4|4|4|4|0|2|3|3|2|2.5|2|3|3|3|2.75|-9.09|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4||3|||3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Yellow||Child/Family: Time constraints|12.3||1|1|1|1|F|Black||19|No|Mother|28278|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||61|28215|Bachelors Degree|Divorced|Self-Employed, Entrepreneur||0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500012459|502427295|31|0|2|502437756|31|0|2|500525086|2||-2||4|2||500000294|-2||-2|0|10|||130|1|||1|259039|256292|4|3|45
500577150|BBBS of Greater Charlotte|Main Office|C|Active|2011-03-22|NaT|Followup|2012-03-22|2012-03-13|Complete|Done|2|2|2|2|2|3|2.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI||71.8||4|5|1|2|F|Black||15||Aunt|28213|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||40|29715|||Customer Service||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500214349|31|0|2|501734288|1|0|2|500526894|2||500004641||2|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|259165||4|3|45
500570756|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-22|2013-02-19|Followup|2012-03-22|2012-03-13|Complete|Done|3|3|3|4|4|3|3.33|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Moved|23||4|5|1|2|F|Black||15||Aunt|28213|Two Parent|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||25|28202|||Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500214349|31|0|2|501865290|1|0|2|500526958|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|259245||4|3|45
501536365|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-03|2014-07-17|Followup|2012-02-03|2012-01-29|Complete|Done|4|4|4|4|4|4|4|||||||||1|4|4|1|2|3|2.5|||||||||4|4|4|4||||||5|5|3|3|4|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||2|2|2|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|65.4||1|1|1|1|M|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Enrollment|M|Black||57|28105|Some College|Married|Retail: Sales|28105|10|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501536657|31|0|1|501443152|31|0|1|500336020|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|259455||4|3|45
500764138|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-07|2013-02-21|Followup|2012-02-07|2012-02-07|Complete|Done|1|2|4|1|4|4|2.67|||||||||2|4|3|1|2|3|2.5|||||||||4|4|4|4||||||5|5|5|3|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||4|2|3|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|72.5||2|2|1|1|M|Black||17|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community|Amachi|Match Support|M|Black||33|28214||Single|Tech: Research/Design||1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500764404|31|0|1|500696779|31|0|1|500154924|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|259457||4|3|45
500938154|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-12|NaT|Followup|2012-01-12|2012-03-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||98.1||2|2|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||32|28208|Associate Degree|Single|Service: Restaurant|28211|4|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500938424|31|0|1|501446421|1|0|1|500323753|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|259488||4|1|45
501811385|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-23|2016-08-19|Followup|2012-03-23|2012-05-02|Complete|Done|4|3|4|4|4|4|3.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI, Cabarrus County|Child: Graduated|64.9||2|2|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||43|28075|Bachelors Degree|Married|Business: Mgt, Admin||7|0|Recruitment Event|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501811730|31|0|2|502460013|31|0|2|500524684|2||-2||4|3|500005291, 500016374|500016374|-2|500016374|-2|6854|8|||7459|10|||1|259753||4|3|45
502102857|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-25|2013-06-18|Followup|2012-03-25|2012-06-09|Expired|Late||||||||4|4|3|1|4|4|3.33|||||||||3|4|3|3|1|4|3||||||4|4|2|3.33|||||||4|4|5|1|3.5||||||||||4|4|4|4|2|4|3|3.57||||||4|4|4|4|||||3|2|2.5||||2|2|||||||Red|2010-2012 OJJDP JJI|Volunteer: Moved|26.8||2|2|1|1|M|Black||18|No|Mother|28278|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||38|28273|Bachelors Degree|Married|Insurance|28202|2|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502103284|31|0|1|502464465|31|0|1|500526162|2||-2||4|3|500005291|500005291|-2|500000294, 500004640|-2|0|4|||7446|3|||1|260346|40474|4|0|45
500186990|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-17|2014-02-28|Followup|2012-02-17|2012-02-17|Complete|Done|4|4|4|2|4|4|3.67|||||||||2|2|3|2|2|3|2.33|||||||||4|4|4|4||||||5|4|2|3|3.5|||||||4|4|4|4|2|4|3|3.57||||||||||3|4|4|3.67||||||2|1|1.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|60.4||2|2|3|3|M|Black||19|Yes|Mother|28269|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||51|28269|Bachelors Degree|Married|Unknown|28202|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500188170|31|0|1|500189496|31|0|1|500339895|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|260439||4|3|45
502418103|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-08|2011-09-07|Baseline|2011-03-29|2011-04-08|Complete|Done|3|2|3|2|3|3|2.67|||||||||1|2|2|3|2|4|2.33|||||||||4|3|4|3.67||||||2|4|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Yellow|2010-2012 OJJDP JJI|Child/Family: Moved|5||1|1|1|1|M|Black||20|No|Mother|28027|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28027|Bachelors Degree|Married|Business: Mgt, Admin|28273|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500002335|502418541|31|0|1|502430938|31|0|1|500528075|2||-2||4|2|500005291|500005291|-2||-2|34|2|||7496|10|||1|261368|-1|4|3|44
500859789|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-29|2013-02-28|Followup|2012-03-29|2012-06-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|71.1||1|1|1|1|F|Black||18|Yes|Mother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||65|28078|||Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500860058|31|0|2|500856753|31|0|2|500169338|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|262144||4|0|45
500896361|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-14|2014-02-27|Followup|2012-01-14|2012-03-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|61.4||2|2|1|1|F|Black||20|Yes|Mother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28075||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500012459|500896631|31|0|2|501276501|31|0|2|500291021|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|262365||4|0|45
500764136|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-10|2012-08-23|Followup|2012-02-10|2012-02-02|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|3|4|4|3.83|||||||||4|3|4|3.67||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|4|2.5|||||1|1||||4|4||||Green|Amachi|Volunteer: Lost contact with child/agency|30.4||3|3|1|1|M|Black||22|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community|Amachi|Match Support|M|White||32|28210|Some College|Single|Business: Mgt, Admin|28206|8|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500764404|31|0|1|501915488|1|0|1|500428501|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|262604||4|3|45
500186905|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-10|2015-11-04|Followup|2012-02-10|2012-02-15|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|4|4|1|4|3|||||||||4|4|4|4||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|1|2.5|||||2|2||||4|4||||Red|Amachi|Child: Graduated|128.8||1|1|1|1|F|Black||19|Yes|Mother|28205|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|F|Black||50|28215|Some College|Single|Finance: Banking||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188151|31|0|2|500189677|31|0|2|500037790|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|262605||4|3|45
501130354|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-15|2012-11-29|Followup|2012-02-15|2012-03-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|57.5||1|1|1|1|M|Black||21|Yes|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||BBBS Board/Staff|General Community|Amachi|Match Support|M|White||43|28205|Bachelors Degree|Married|Finance: Banking||7|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501130628|31|0|1|501124346|1|0|1|500245525|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|13|||46|2|||1|262610||4|1|45
500892914|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-16|2014-09-11|Followup|2012-02-16|2012-03-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Graduated|54.8||2|2|1|1|M|Black||20|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Sales|28269|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500893173|31|0|1|501964388|1|0|1|500429157|2||500003586||4|3|500000294|500000294|-2||-2|0|5|||7464|9|||1|262612||4|1|45
500843863|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-21|2016-06-17|Followup|2012-02-21|2012-03-29|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|4|2|3|3|||||||||4|4|4|4||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|Amachi|Volunteer: Changed workplace/school partnership|99.8||2|2|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|No|TV|Media|General Community|Amachi|Match Support|F|Black||32|28269|Bachelors Degree|Single|Business: Marketing|28273|0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500844129|31|0|2|501078655|31|0|2|500241388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|56|1|||2238|7|||1|262613||4|3|45
500544921|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2013-08-29|Followup|2012-03-31|2012-05-15|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi, Project Big, Project Big AND Amachi|Child: Lost interest|29||2|2|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$15,000 to $19,999|Y|No|TV|Media|General Community|Project Big AND Amachi|Match Support|M|White||31|28211|Bachelors Degree|Married|Finance: Banking|28202|0|2|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011746|500545173|31|0|1|502079132|1|0|1|500523387|2||500004772||4|3|500000294, 500004640, 500004901|500004901|-2||-2|56|1|||7464|9|||1|262640||4|1|45
502495123|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2013-01-08|Followup|2012-03-31|2012-03-05|Complete|Early|4|4|2|4|1|4|3.17|3|4|4|2|1|4|3|5.67|4|1|3|4|1|4|2.83|2|4|4|4|4|4|3.67|-22.89|4|3|4|3.67|4|3|4|3.67|0|5|4|5|4|4.5|5|3|3|4|3.75|20|4|4|4|4|4|4|3|3.86|4|4|4|4|4|||||4|3|3|3.33|4|4|4|4|-16.75|3|1|2|||||2|2||||4|4|4|4|0|Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|21.3||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28207|Bachelors Degree|Single|Finance: Economist|28255|5|0||Relative|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502495572|31|0|2|502473441|1|0|2|500524205|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||0|11|||1|262685|254961|4|3|45
501631547|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2016-07-29|Followup|2012-03-31|2012-05-02|Complete|Done|3|2|2|2|3|3|2.5|||||||||4|4|3|3|3|4|3.5|||||||||4|4|4|4||||||3|2|3|4|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child: Graduated|64||2|2|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||38|28277|Bachelors Degree|Single|Arts, Entertainment, Sports|28203|3|6|UnitedMethodistChrch|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|501631870|31|0|1|502170945|1|0|1|500528464|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||8529|7|||1|262703||4|3|45
501868921|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2016-07-29|Followup|2012-03-31|2012-05-02|Complete|Done|3|4|4|4|3|3|3.5|3|1|1|1|1|2|1.5|133.33|2|3|3|1|2|4|2.5|3|2|4|4|4|4|3.5|-28.57|4|4|3|3.67|4|3|3|3.33|10.21|3|5|4|3|3.75|4|5|5|4|4.5|-16.67|4|4|4|4|3|3|3|3.57|4|4|4|4|3|3|3|3.57|0|3|3|3|3|2|4|3|3|0|3|3|3|2|1|1.5|100|2|2|1|1|100|4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Moved|64||2|2|2|2|F|Black||19|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28211||Married|Finance: Banking|28255|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501869291|31|0|2|501382633|1|0|2|500524206|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|262708|4527|4|3|45
501628854|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2012-11-29|Followup|2012-03-31|2012-04-02|Complete|Done|4|1|2|1|2|3|2.17|||||||||2|2|3|2|2|3|2.33|||||||||4|4|4|4||||||2|3|2|2|2.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|4|3|||||2|2||||4|4||||Green||Volunteer: Moved|20||3|3|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||33|28277|Bachelors Degree|Married|Finance|28209|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|501629177|31|0|2|502091655|1|0|2|500521158|2||500003586||4|1||500000294|-2||-2|0|10|||7496|10|||1|262943||4|3|45
501588821|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-10|2012-05-23|Followup|2012-02-10|2012-04-26|Expired|Late||||||||4|1|2|1|3|3|2.33|||||||||1|4|3|1|1|4|2.33||||||4|4|4|4|||||||5|1|1|2|2.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|4|3||||2|2|||||||Green||Volunteer: Lost contact with child/agency|27.4||1|1|2|2|F|Black||16||Mother|28208|Two Mothers|Unknown||Yes||Self|General Community||Match Support|F|Black||34|28273|Masters Degree|Living w/ Significant Other|Consultant|28273|1|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501589141|31|0|2|501359582|31|0|2|500429105|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|263163|28524|4|0|45
500417525|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-17|2012-11-30|Followup|2012-01-17|2012-02-26|Complete|Done|4|3|4|3|4|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Project Big|Volunteer: Time constraint|70.4||1|1|1|1|M|Black||18||Mother|28208|One Parent: Female|Unknown||No|TV|Media|General Community|Project Big|Match Support|M|White||37|28202|||Medical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500417775|31|0|1|500755435|1|0|1|500151964|2||500004641||4|1|500004640|500004640|-2||-2|56|1|||46|2|||1|263425||4|3|45
502494753|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-14|2013-10-22|Baseline|2011-04-04|2011-04-14|Complete|Done|4|3|3|1|4|3|3|||||||||2|3|2|3|1|4|2.5|||||||||4|4|4|4||||||1|4|3|5|3.25|||||||4|4|4|4|4|4|4|4||||||||||1|4|4|3||||||4|2|3|||||1|1|||||||||Yellow|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|30.3||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28212|Masters Degree|Single|Business|28105|5|8|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500011746|502495202|31|0|2|502481799|31|0|2|500529173|2||500004772||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|4|||7438|1|||1|263617|-1|4|3|44
501777213|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-04|2012-05-22|Followup|2012-04-04|2012-03-05|Complete|Early|4|3|3|3|4|4|3.5|4|1|3|1|2|4|2.5|40|3|4|4|3|3|4|3.5|2|4|3|3|3|3|3|16.67|4|4|4|4|4|4|4|4|0|5|4|3|5|4.25|5|1|2|4|3|41.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|4|4|2|3.33|0|4|3|3.5|2|2|2|75|2|2|2|2|0|4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Moved|13.6||2|2|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||33|28202|Bachelors Degree|Single|Finance: Banking|28255|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500011746|501777568|31|0|1|502475369|31|0|1|500527844|2||-2||4|1|500005291|500005291|-2|500005291|-2|0|10|||7496|10|1202|1|1|263749|21893|4|3|45
501553185|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-23|2012-06-29|Followup|2012-02-23|2012-03-05|Complete|Done|4|4|2|3|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|40.1||1|1|1|1|M|Black||14|No|Mother|28277|One Parent: Female|Unknown||No|Brochure|Media|General Community||Match Support|M|Black||47|28262|Juris Doctorate (JD)|Married|Law: Lawyer|28262|10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501553481|31|0|1|501556179|31|0|1|500342698|2||-2||4|1|||-2||-2|51|1|||7464|9|||1|263866||4|3|45
500186798|BBBS of Greater Charlotte|Main Office|C|Completed|2005-03-30|2015-10-20|Followup|2012-03-30|2012-05-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Time constraints|126.7||1|2|1|2|F|Multi-Race (None of the above)||19|No|Father|28208|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||45|28226|Bachelors Degree||Business: Human Resources||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500187961|7|0|2|500189825|1|0|2|500038158|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|264100||4|1|45
500850236|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-04|2013-09-16|Followup|2012-04-04|2012-05-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|77.4||1|1|2|2|M|Black||21|No|Mother|28205|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|Black||37|28262|Bachelors Degree|Single|Real Estate: Realtor||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500850505|31|0|1|500189198|31|0|1|500169235|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|264121||4|1|45
500868942|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-20|NaT|Followup|2011-09-20|2011-11-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||113.8|Y|1|1|1|1|M|Black||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|M|White||54|28207||Married|Business: Sales||0|0|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500869211|31|0|1|500947018|1|0|1|500195082|2||-2||2|1|||-2||-2|0|10|||7458|9|||1|264269||4|1|45
500185781|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-13|2012-04-30|Followup|2012-02-13|2012-02-13|Complete|Done|3|2|4|3|4|2|3|||||||||3|4|4|2|3|3|3.17|||||||||4|4|4|4||||||4|3|5|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||2|2|1|1.67||||||4|4|4|||||1|1||||4|4||||Red||Child: Graduated|50.5||2|2|2|2|M|Black||23||Mother|28262|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||34|28105||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013709|500187370|31|0|1|500188751|1|0|1|500244796|2||||4|3|||-2||-2|6854|8|||7464|9|||1|264508||4|3|45
502539860|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-15|2014-02-10|Baseline|2011-04-06|2011-04-15|Complete|Done|3|2|1|1|1|4|2|||||||||2|3|3|3|2|3|2.67|||||||||2|2|2|2||||||3|2|1|1|1.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33|||||||||||||1|1||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|33.9||1|1|1|1|M|Hispanic||17|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Hispanic||33|28270|Associate Degree|Married|Business: Sales||9|0|Other|BBBS Board/Staff|Big|General Community|Project Big|Match Support|277|60|598|500000170|500017777|502540313|3|0|1|502498837|3|0|1|500529729|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||7671|13|||1|264531|-1|4|3|44
500997880|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-19|2016-07-29|Followup|2012-02-19|2012-04-13|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|101.3||1|1|1|1|M|Black||18|No|Mother|28204|Two Parent|$40,000 to $44,999||Yes||Self|General Community||Match Support|M|White||33|28202|Bachelors Degree|Married|Business: Marketing||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500998153|31|0|1|500990660|1|0|1|500237316|2||-2||4|1|||-2||-2|0|10|||46|2|||1|264538||4|1|45
502501319|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2011-10-25|Baseline|2011-04-08|2011-04-26|Complete|Done|3|2|3|3|2|3|2.67|||||||||2|4|3|2|1|3|2.5|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|1|1.5|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|5.9||2|2|1|1|F|Black||18|No|Mother|28269|One Parent: Female|$45,000 to $49,999||No||Relative|General Community|2010-2012 OJJDP JJI|Match Support|F|White||57|28269|Associate Degree|Single|Business: Sales|10580|14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011184|502501768|31|0|2|502507619|1|0|2|500530032|2||-2||4|1|500005291|500005291|-2||-2|0|3|||7464|9|||1|265141|-1|4|3|44
500566159|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-23|2012-03-12|Followup|2012-01-23|2012-01-23|Complete|Done|4|3|4|3|4|4|3.67|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|49.6||2|2|1|1|F|Black||16||Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Enrollment|F|White||35|28207|||Business: Clerical||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|500565754|31|0|2|500966678|1|0|2|500230690|2||-2||4|2|||-2||-2|34|2|||46|2|||1|265413||4|3|45
501361902|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-23|NaT|Followup|2012-01-23|2012-01-13|Complete|Done|3|3|4|3|4|4|3.5|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green|Amachi||97.7||1|1|1|1|M|White||17|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28227|Bachelors Degree|Divorced|Business: Sales|28273|9|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501249611|1|0|1|501307192|1|0|1|500328424|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|265427||4|3|45
502229042|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-30|2013-02-22|Followup|2011-09-30|2011-09-15|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|28.8||3|3|1|1|F|Black||14|No|Mother|28269|Two Parent|Unknown||Yes||Relative|General Community||Match Support|F|White||35|28211||Single|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502172965|31|0|2|502272069|1|0|2|500470500|2||-2||4|2|||-2|500000294|-2|0|3|||7496|10|||1|265615||4|1|45
501011735|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-11|2015-03-05|Followup|2012-04-11|2012-04-09|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|2010-2012 OJJDP JJI|Child: Lost interest|46.8||3|3|1|1|F|Black||17||Mother|28215|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28215|High School Graduate|Married|Finance: Banking|28255|13|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500012459|500417756|31|0|2|502473442|31|0|2|500528270|2||-2||4|2|500005291|500005291|-2||-2|0|10|||7446|3|||1|265863||4|3|45
500887862|BBBS of Greater Charlotte|Main Office|C|Active|2011-04-13|NaT|Followup|2012-04-13|2012-04-11|Complete|Done|4|4|4|4|3|4|3.83|||||||||2|3|4|2|2|3|2.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Cabarrus County||71.1||2|2|2|2|F|Black||18|Yes|Mother|28025|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|F|Black||43|28027||Divorced|Finance: Banking||0|7|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500888132|31|0|2|500923430|31|0|2|500530980|2||500016307||2|1|500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|266741||4|3|45
502494753|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-14|2013-10-22|Followup|2012-04-14|2012-05-16|Declined|Done||||||||4|3|3|1|4|3|3|||||||||2|3|2|3|1|4|2.5||||||4|4|4|4|||||||1|4|3|5|3.25||||||||||4|4|4|4|4|4|4|4||||||1|4|4|3|||||4|2|3||||1|1|||||||Yellow|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|30.3||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28212|Masters Degree|Single|Business|28105|5|8|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500011746|502495202|31|0|2|502481799|31|0|2|500529173|2||500004772||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|4|||7438|1|||1|267188|263617|4|1|45
502548212|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2012-12-19|Baseline|2011-04-14|2011-04-29|Complete|Done|4|3|3|2|4|3|3.17|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Moved|19.7||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||28|28210|Bachelors Degree|Single|Business: Marketing||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502548665|31|0|2|502469646|31|0|2|500531329|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|267347|-1|4|3|44
502539860|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-15|2014-02-10|Followup|2012-04-15|2012-04-11|Complete|Done|2|1|1|1|3|4|2|3|2|1|1|1|4|2|0|1|2|3|1|1|3|1.83|2|3|3|3|2|3|2.67|-31.46|4|4|4|4|2|2|2|2|100|3|3|3|3|3|3|2|1|1|1.75|71.43|4|3|4|4|4|4|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|3|4|3|3.33|20.12|4|4|4|||||2|2|1|1|100|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|33.9||1|1|1|1|M|Hispanic||17|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Hispanic||33|28270|Associate Degree|Married|Business: Sales||9|0|Other|BBBS Board/Staff|Big|General Community|Project Big|Match Support|277|60|598|500000170|500017777|502540313|3|0|1|502498837|3|0|1|500529729|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||7671|13|||1|267762|264531|4|3|45
500791567|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-31|2013-04-11|Followup|2012-01-31|2012-01-24|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|4|3|3|3|4|3.17|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|74.3||1|1|2|2|M|Multi-Race (None of the above)||18|No|Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|M|Black||32|28215||Married|Finance: Banking||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|500187654|7|0|1|500578720|31|0|1|500155823|2||-2||4|2|||-2||-2|0|10|||7447|3|||1|268058||4|3|45
500185678|BBBS of Greater Charlotte|Main Office|C|Completed|2003-02-23|2012-07-31|Followup|2012-02-23|2012-05-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|113.2||1|1|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28277|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|500187309|31|0|1|500188619|31|0|1|500036619|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|268399||4|0|45
502482929|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-16|2011-12-13|Baseline|2011-04-19|2011-05-16|Complete|Done|4|2|4|4|4|4|3.67|||||||||2|3|1|2|4|2|2.33|||||||||4|4|4|4||||||1|5|4|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|6.9||1|1|1|1|M|Black||18|No|Mother|28078|One Parent: Female|Less than $10,000|Y|Yes|Billboard|Media|General Community|2010-2012 OJJDP JJI|RTBM|M|Black||31|28227||Single|Retail: Mgt|28104|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502483376|31|0|1|502489447|31|0|1|500531863|2||-2||4|3|500005291|500005291|-2||-2|50|1|||7496|10|||1|268803|-1|4|3|44
502495501|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-20|NaT|Baseline|2011-04-19|2011-05-20|Complete|Done|3|1|4|2|2|2|2.33|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||5|3|2|3|3.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||2|1|1.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI||69.9||1|1|1|1|M|White||15|No|Mother|28226|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||55|28210|Bachelors Degree|Married|Finance|28203|1|6|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500018851|502495950|1|0|1|502508181|1|0|1|500531873|2||-2||2|1|500005291|500005291|-2|500005291|-2|0|10|||7464|9|||1|268809|-1|4|3|44
502530227|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2014-10-20|Baseline|2011-04-19|2011-05-04|Complete|Done|4|1|1|2|4|4|2.67|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|3|4|3|4|3.71||||||||||3|4|3|3.33||||||2|4|3|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|41.6||1|1|1|1|F|Hispanic||15|No|Mother|28213|One Parent: Female|$10,000 to $14,999||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||30|28210|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502530676|3|0|2|502531485|3|0|2|500532078|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|268895|-1|4|3|44
501765404|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-20|2013-08-29|Followup|2012-04-20|2012-06-08|Declined|Late||||||||3|3|3|1|4|3|2.83|||||||||2|3|3|2|3|3|2.67||||||4|4|4|4|||||||3|5|5|4|4.25||||||||||4|4|4|3|2|3|1|3||||||4|3|4|3.67|||||4|3|3.5||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|40.3||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Multi-race (Black & White)||28|28262||Single|Student: College|28262|3|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501765751|31|0|1|501958658|36|0|1|500443642|2||-2||4|2|||-2||-2|0|10|||9221|5|||1|268962|36416|4|1|45
501160887|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2013-05-14|Followup|2011-04-30|2011-06-08|Complete|Done|3|2|4|4|4|4|3.5|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|2|3|||||2|2|||||||||Green|Amachi|Volunteer: Time constraint|36.5||2|2|1|1|F|Black||14|Yes|Mother|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Enrollment|F|White||58|28226|||Education: Teacher Asst/Aid|28203|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|501615415|1|0|2|500447312|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|269146||4|3|45
502530223|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2013-05-21|Baseline|2011-04-20|2011-04-29|Complete|Done|3|2|1|1|2|2|1.83|||||||||1|3|2|1|2|2|1.83|||||||||3|4|4|3.67||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|24.7||1|1|1|1|M|Hispanic||16||Mother|28213|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||44|28078|Masters Degree|Married|Business|28036|8|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502530676|3|0|1|502501248|3|0|1|500533054|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|269200|-1|4|3|44
501868918|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-27|2014-05-22|Followup|2012-05-27|2012-05-02|Complete|Early|3|4|4|4|3|3|3.5|3|3|3|4|3|3|3.17|10.41|2|3|3|4|2|4|3|3|4|4|2|3|3|3.17|-5.36|4|4|3|3.67|4|4|3|3.67|0|3|5|4|3|3.75|3|3|5|5|4|-6.25|4|4|4|4|3|3|3|3.57|3|4|3|3|4|3|2|3.14|13.69|3|3|3|3|3|4|3|3.33|-9.91|3|2|2.5|2|3|2.5|0|2|2|1|1|100|4|4||||Green||Child: Graduated|47.8||1|1|1|1|M|Black||20|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||35|27612|Juris Doctorate (JD)|Living w/ Significant Other|Law|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|501869291|31|0|1|501921115|1|0|1|500454496|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|269399|128915|4|3|45
500186702|BBBS of Greater Charlotte|Main Office|C|Completed|2004-04-28|2014-11-25|Followup|2012-04-28|2012-06-12|Complete|Done|4|4|4|4|4|4|4|||||||||3|2|3|3|3|3|2.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|126.9||1|2|1|2|F|Black||20|Yes|GrandMother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||57|28212|Some College|Married|Unknown||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|RTBM|277|60|598|500000170|500017732|500188150|31|0|2|500189528|31|0|2|500038225|2||500003586||4|1|500000294|500000294|-2|500015184|-1|0|10|||7462|13|||1|269438||4|3|45
502106926|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-25|2012-06-28|Followup|2012-05-25|2012-06-28|Blank|Done||||||||4|4|4|1|2|4|3.17|||||||||1|2|4|3|3|3|2.67||||||4|4|4|4|||||||5|1|5|1|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Red||Volunteer: Time constraint|25.1||2|2|1|1|M|Black||17|No|Mother|28031|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28031||Single|Govt||0|0|AA Task Force|Special Event|Big|General Community||Match Support|277|60|598|500000170|500011746|502107353|31|0|1|502072628|1|0|1|500453665|2||-2||4|3|||-2||-2|0|10|||11098|8|||1|269485|40460|4|3|45
502478428|BBBS of Greater Charlotte|Main Office|C|Active|2011-04-28|NaT|Baseline|2011-04-21|2011-04-28|Complete|Done|4|4|1|4|4|4|3.5|||||||||4|2|4|2|4|4|3.33|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI||70.6||1|1|1|1|M|White||16|No|Mother|28277|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||54|28205|Some College|Separated|Self-Employed, Entrepreneur|28214|29|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502478875|1|0|1|502555822|1|0|1|500533009|2||-2||2|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|270021|-1|4|3|44
502173445|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-23|2013-09-26|Baseline|2011-04-21|2011-05-23|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|4|3|3|4|3|3.17|||||||||4|3|4|3.67||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2|||||||||Red|Amachi|Volunteer: Lost contact with child/agency|28.2||1|1|1|1|F|Black||19|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Service Organization|General Community|Amachi|Match Support|F|White||28|28206|Bachelors Degree|Single|Education: Teacher||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502173869|31|0|2|502266833|1|0|2|500532710|2||500003586||4|3|500000294|500000294|-2||-2|0|11|||7464|9|||1|270032|-1|4|3|44
501389722|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-06|2014-04-24|Followup|2012-02-06|2012-02-07|Complete|Done|3|4|4|1|3|3|3|||||||||3|3|4|2|3|4|3.17|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Graduated|62.5||1|1|1|1|F|White||21|No|Mother|28027|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||56|28027||Divorced|Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500012459|501390003|1|0|2|500787778|1|0|2|500337267|2||-2||4|1|||-2||-2|0|10|||46|2|||1|270704||4|3|45
502540400|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-25|2012-01-26|Baseline|2011-04-23|2011-04-25|Complete|Done|4|1|3|1|4|3|2.67|||||||||1|1|1|2|1|1|1.17|||||||||4|4|4|4||||||3|2|3|2|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||1|1||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Agency: Challenges with program/partnership|9.1||1|1|1|1|M|Black||16|No|GrandMother|28208|Grandparents|Unknown|Y|Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||68|28025||Widowed|Education|28212|5|0|A Child's Place|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500012459|502540853|31|0|1|502540283|1|0|1|500533007|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|7016|11|||11610|6|1210|1|1|270759|-1|4|3|44
502537639|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-26|2012-05-31|Baseline|2011-04-23|2011-04-26|Complete|Done|3|1|1|2|4|4|2.5|||||||||2|3|1|1|3|4|2.33|||||||||4|4|4|4||||||2|3|5|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|13.2||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|White||39|28209|Bachelors Degree|Single|Finance: Banking|28202|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013709|502538092|31|0|2|502387375|1|0|2|500533008|2||-2||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||46|2|||1|270760|-1|4|3|44
502570188|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Baseline|2011-04-26|2011-04-30|Complete|Done|4|3|3|2|4|4|3.33|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|69.8||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||56|28226|Masters Degree|Married|Medical: Nurse|28217|34|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570642|31|0|2|502366830|1|0|2|500533448|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||10326|3|||1|271777|-1|4|3|44
502568883|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-13|2012-05-31|Baseline|2011-04-26|2011-05-13|Complete|Done|2|3|4|1|1|4|2.5|||||||||2|2|4|2|1|4|2.5|||||||||4|4|4|4||||||5|2|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|12.6||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|$15,000 to $19,999||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||30|28262|Masters Degree|Single|Customer Service|28262|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502569337|31|0|2|502501016|31|0|2|500533467|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|271809|-1|4|3|44
502162474|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2013-02-28|Baseline|2011-04-26|2011-05-04|Complete|Done|3|4|4|3|3|4|3.5|||||||||3|3|2|3|4|4|3.17|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|21.9||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||35|28205|Associate Degree|Single|Student: College|28213|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502162903|31|0|1|502536516|1|0|1|500533468|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7496|10|||1|271811|-1|4|3|44
501938282|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-17|NaT|Followup|2011-11-17|2011-11-02|Complete|Done|3|3|3|3|3|3|3|||||||||1|2|2|2|2|2|1.83|||||||||4|4|4|4||||||1|3|1|3|2|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi, Cabarrus County||75.9||1|1|1|1|F|White||14|Yes|Mother|28025|Two Parent|Unknown|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||63|28027|High School Graduate|Married|Self-Employed, Entrepreneur|28027|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501938680|1|0|2|502356100|1|0|2|500493871|2||500016307||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|271939||4|3|45
502431187|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-21|2012-04-20|Baseline|2011-04-27|2011-07-21|Complete|Done|3|2|4|1|3|4|2.83|||||||||2|3|3|2|3|3|2.67|||||||||2|4|4|3.33||||||4|3|5|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|2|3|2.67||||||2|3|2.5|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|9||2|2|1|1|F|Black||17|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|RTBM|F|Black||27|28262|Some College|Single|Retail: Sales||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502431630|31|0|2|502616530|31|0|2|500545377|2||-2||4|3|500005291|500005291|-2||-2|0|5|||7464|9|||1|272216|-1|4|3|44
500968246|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-29|2015-04-30|Followup|2012-04-29|2012-06-10|Complete|Done|3|3|2|2|3|3|2.67|||||||||2|3|2|3|3|4|2.83|||||||||4|3|3|3.33||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|84||1|1|1|1|M|Black||19|No|Aunt|28269|One Parent: Female|$10,000 to $14,999|Y|No||Therapist/Counselor|General Community||Match Support|M|Black||35|28213|Bachelors Degree|Single|Business: Sales||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500968516|31|0|1|501179573|31|0|1|500251681|2||-2||4|1|||-2||-2|0|5|||46|2|||1|272381||4|3|45
501015965|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-29|2013-10-09|Followup|2012-04-29|2012-04-23|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|3|4|3|3|3|3.17|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2||||4|4||||Yellow|Amachi|Child: Lost interest|41.4||2|2|2|2|F|Black||17|Yes|Mother|28208|One Parent: Female|Less than $10,000||Yes||Self|General Community|Amachi|Match Support|F|Black||60|28269|Bachelors Degree|Married|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|500189376|31|0|2|500447721|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|272383||4|3|45
502478428|BBBS of Greater Charlotte|Main Office|C|Active|2011-04-28|NaT|Followup|2012-04-28|2012-04-19|Complete|Done|3|4|4|4|3|4|3.67|4|4|1|4|4|4|3.5|4.86|2|4|3|1|4|3|2.83|4|2|4|2|4|4|3.33|-15.02|4|4|4|4|4|4|4|4|0|4|4|4|5|4.25|4|5|5|5|4.75|-10.53|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|4|4|-8.25|2|4|3|2|4|3|0|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||70.6||1|1|1|1|M|White||16|No|Mother|28277|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||54|28205|Some College|Separated|Self-Employed, Entrepreneur|28214|29|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502478875|1|0|1|502555822|1|0|1|500533009|2||-2||2|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|272553|270021|4|3|45
500791645|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-28|2012-09-27|Followup|2012-04-28|2012-04-23|Complete|Done|3|4|2|2|1|3|2.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Child/Family: Feels incompatible with volunteer|17||4|4|1|1|F|Multi-Race (None of the above)||15||Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||27|28213|Some College|Single|Education|28235|0|6||Relative|Big|General Community||RTBM|277|60|598|500000170|500012459|500187654|7|0|2|502524278|31|0|2|500529175|2||-2||4|3|500005291|500005291|-2||-2|0|10|||0|11|||1|272599||4|3|45
502530223|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2013-05-21|Followup|2012-04-29|2012-05-22|Complete|Done|3|2|2|1|4|3|2.5|3|2|1|1|2|2|1.83|36.61|1|3|3|1|2|2|2|1|3|2|1|2|2|1.83|9.29|2|3|3|2.67|3|4|4|3.67|-27.25|2|3|3|2|2.5|3|2|4|4|3.25|-23.08|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|24.7||1|1|1|1|M|Hispanic||16||Mother|28213|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||44|28078|Masters Degree|Married|Business|28036|8|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502530676|3|0|1|502501248|3|0|1|500533054|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|273218|269200|4|3|45
502548212|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2012-12-19|Followup|2012-04-29|2012-04-19|Complete|Done|4|4|4|1|4|4|3.5|4|3|3|2|4|3|3.17|10.41|2|4|3|4|4|3|3.33|2|4|3|3|2|3|2.83|17.67|4|4|4|4|4|4|4|4|0|3|1|1|1|1.5|2|3|3|3|2.75|-45.45|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3|3|3|33.33|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Moved|19.7||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||28|28210|Bachelors Degree|Single|Business: Marketing||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502548665|31|0|2|502469646|31|0|2|500531329|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|273252|267347|4|3|45
502224918|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-10|2011-10-12|Baseline|2011-04-29|2011-05-10|Complete|Done|3|3|4|1|3|4|3|||||||||4|4|3|3|2|4|3.33|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|5.1||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|M|Asian||31|28202||Single|Law: Lawyer|28202|2|4|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014, Project Big|RTBM|277|60|598|500000170|500011639|502225349|31|0|1|502448424|4|0|1|500533984|2||-2||4|3|500005291|500005291|-2|500004640, 500014506|-1|0|10|||7671|13|||1|273352|-1|4|3|44
502137546|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2015-10-20|Followup|2012-04-29|2012-06-27|Comprehension|Late||||||||4|4|2|2|4|4|3.33|||||||||2|4|3|2|2|3|2.67||||||4|4|4|4|||||||4|3|5|4|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|4|3.5||||2|2|||||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|53.7||1|2|1|2|F|Black||16||Mother|28213|Other/Unknown|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28262|||Business: Mgt, Admin|75234|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502137975|31|0|2|501641708|31|0|2|500520728|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|273564|36419|4|2|45
502570183|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Baseline|2011-04-30|2011-04-30|Complete|Done|3|3|4|3|4|3|3.33|||||||||4|4|4|4|4|3|3.83|||||||||4|4|3|3.67||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Amachi, Project Big, Project Big AND Amachi|Agency: Challenges with program/partnership|69.8||1|1|1|1|F|Black||17|Yes|Mother|28206|Other/Unknown|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||61|28134|Bachelors Degree|Married|Medical: Admin||33|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570637|31|0|2|502570153|31|0|2|500534090|2||500004772||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|273709|-1|4|3|44
502570183|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Followup|2012-04-30|2012-05-22|Complete|Done|4|3|3|4|4|4|3.67|3|3|4|3|4|3|3.33|10.21|2|2|3|2|3|4|2.67|4|4|4|4|4|3|3.83|-30.29|4|4|4|4|4|4|3|3.67|8.99|2|2|2|2|2|3|3|4|3|3.25|-38.46|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|3|3.67|4|4|4|4|-8.25|2|4|3|3|3|3|0|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Agency: Challenges with program/partnership|69.8||1|1|1|1|F|Black||17|Yes|Mother|28206|Other/Unknown|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||61|28134|Bachelors Degree|Married|Medical: Admin||33|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570637|31|0|2|502570153|31|0|2|500534090|2||500004772||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|273711|273709|4|3|45
502570188|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Followup|2012-04-30|2012-04-23|Complete|Done|3|4|4|4|4|2|3.5|4|3|3|2|4|4|3.33|5.11|4|3|4|4|4|4|3.83|2|4|4|2|3|4|3.17|20.82|4|4|4|4|4|4|4|4|0|4|4|2|3|3.25|5|5|5|4|4.75|-31.58|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|3|2|2.5|2|2|2|25|1|1|2|2|-50|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|69.8||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||56|28226|Masters Degree|Married|Medical: Nurse|28217|34|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570642|31|0|2|502366830|1|0|2|500533448|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||10326|3|||1|273717|271777|4|3|45
501365904|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-20|2012-09-05|Followup|2012-04-20|2012-06-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Moved|40.5||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown|Y|No||Self|General Community||Enrollment|M|Black||48|28269|Some College|Married|Business: Engineer|28262|20|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501366183|31|0|1|501459709|31|0|1|500353421|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|274310||4|1|45
502537469|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2012-08-31|Baseline|2011-05-02|2011-05-04|Complete|Done|4|2|3|4|3|4|3.33|||||||||3|4|3|2|3|3|3|||||||||3|4|3|3.33||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|4|3|||||2|2||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|15.9||3|3|1|1|F|Black||16|No|Mother|28208|One Parent: Female|$15,000 to $19,999||No||School|General Site||Match Support|F|White||38|28205|Bachelors Degree|Divorced|Customer Service||1|3|TV|Media|Big|General Community|Project Big|Match Support|277|60|598|500000170|500001281|502537922|31|0|2|502227984|1|0|2|500534571|2||500004641||4|2|500004640, 500005291||-1|500004640|-2|0|4|||130|1|1204|3|1|274447|-1|4|3|44
500781988|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-16|2013-09-04|Followup|2012-02-16|2012-05-02|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|78.6||1|1|1|1|M|White||21||Mother|28027||Unknown||No||Self|General Community||Match Support|M|White||71|28083|Some College|Married|Business: Mgt, Admin|28027|13|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500002335|500782256|1|0|1|500773716|1|0|1|500160560|2||-2||4|1|||-2||-2|0|10|||46|2|||1|274758||4|0|45
502287066|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-03|2014-09-04|Followup|2012-05-03|2012-05-22|Complete|Done|4|4|4|4|4|3|3.83|||||||||2|3|3|2|2|4|2.67|||||||||4|4|3|3.67||||||3|3|3|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|40.1||2|2|1|1|M|Black||15||GrandMother|28227|One Parent: Female|Unknown|Y|Yes|AARTF|BBBS Board/Staff|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28215|Associate Degree|Married|Medical: Nurse||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502287498|31|0|1|502501212|1|0|1|500532817|2||-2||4|1|500005291|500005291|-2||-2|7294|13|||7464|9|||1|274962||4|3|45
502566369|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-18|2012-04-30|Baseline|2011-05-03|2011-05-18|Complete|Done|3|1|4|2|4|4|3|||||||||4|4|4|1|3|4|3.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|11.4||2|2|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||31|28105|Bachelors Degree|Single|Tech: Production Line|28203|3|8|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500011746|502566823|31|0|2|502484867|31|0|2|500534744|2||-2||4|2|500005291||-2|500005291|-2|0|10|||7464|9|||1|275023|-1|4|3|44
502567548|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-27|2012-10-31|Baseline|2011-05-03|2011-05-27|Complete|Done|3|4|3|4|4|4|3.67|||||||||4|4||4|4|4||||||||||4|4|4|4||||||5|2|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Red|Amachi, Project Big AND Amachi|Child/Family: Moved|17.2||1|1|2|2|F|Hispanic||16|Yes|Mother|28227|One Parent: Female|Unknown||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502568002|3|0|2|502564910|31|0|2|500534824|2||500003586||4|3|500000294, 500004901|500004640, 500004901|-2||-2|0|4|||17161|11|||1|275240|-1|4|3|44
502162474|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2013-02-28|Followup|2012-05-04|2012-06-29|Declined|Late||||||||3|4|4|3|3|4|3.5|||||||||3|3|2|3|4|4|3.17||||||4|4|4|4|||||||5|4|4|5|4.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|21.9||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||35|28205|Associate Degree|Single|Student: College|28213|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502162903|31|0|1|502536516|1|0|1|500533468|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7496|10|||1|275652|271811|4|1|45
502530227|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2014-10-20|Followup|2012-05-04|2012-05-03|Complete|Done|1|4|1|1|2|4|2.17|4|1|1|2|4|4|2.67|-18.73|4|3|4|2|4|4|3.5|2|4|4|2|3|4|3.17|10.41|2|2|2|2|4|4|4|4|-50|3|4|3|3|3.25|5|5|4|5|4.75|-31.58|4|4|4|3|4|4|4|3.86|4|4|4|3|4|3|4|3.71|4.04|4|4|2|3.33|3|4|3|3.33|0|4|4|4|2|4|3|33.33|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|41.6||1|1|1|1|F|Hispanic||15|No|Mother|28213|One Parent: Female|$10,000 to $14,999||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||30|28210|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502530676|3|0|2|502531485|3|0|2|500532078|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|275956|268895|4|3|45
502537469|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2012-08-31|Followup|2012-05-04|2012-05-25|Declined|Done||||||||4|2|3|4|3|4|3.33|||||||||3|4|3|2|3|3|3||||||3|4|3|3.33|||||||3|3|4|5|3.75||||||||||4|4|4|4|4|4|4|4||||||3|4|4|3.67|||||2|4|3||||2|2||||4|4||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|15.9||3|3|1|1|F|Black||16|No|Mother|28208|One Parent: Female|$15,000 to $19,999||No||School|General Site||Match Support|F|White||38|28205|Bachelors Degree|Divorced|Customer Service||1|3|TV|Media|Big|General Community|Project Big|Match Support|277|60|598|500000170|500001281|502537922|31|0|2|502227984|1|0|2|500534571|2||500004641||4|2|500004640, 500005291||-1|500004640|-2|0|4|||130|1|1204|3|1|275960|274447|4|1|45
502402515|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-17|2015-12-28|Baseline|2011-05-05|2011-05-17|Complete|Done|3|1|3|1|1|4|2.17|||||||||1|4|3|1|3|4|2.67|||||||||4|4|4|4||||||3|2|2|2|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|3|3.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|55.4||1|1|1|1|M|Black||16|No|Mother|28215|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28215||Single|Law: Police Officer||14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502402953|31|0|1|502537081|31|0|1|500535130|2||-2||4|1|500005291|500005291|-2||-2|34|2|||7464|9|||1|276236|-1|4|3|44
500546821|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-21|2015-09-15|Followup|2012-02-21|2012-04-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|102.8||1|1|3|3|M|Black||20|No|Mother|28083|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||52|28025||Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500012459|500547073|31|0|1|500790181|31|0|1|500159910|2||-2||4|1|||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|277356||4|1|45
502179818|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-16|2013-02-26|Followup|2011-07-16|2011-07-06|Complete|Done|4|3|4|4|1|4|3.33|||||||||1|4|4|2|4|4|3.17|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Yellow|Amachi|Volunteer: Moved|31.4||1|1|1|1|F|Black||14|Yes|GrandMother|28216|Grandparents|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Enrollment|F|Black||28|28216||Single|Student: College||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502180247|31|0|2|502057930|31|0|2|500460281|2||500003586||4|2|500000294|500000294|-2|500000294|-2|5635|9|||7464|9|||1|277414||4|3|45
502537477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-12|2016-07-14|Baseline|2011-05-09|2011-05-12|Complete|Done|3|2|1|1|3|3|2.17|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||2|3|2|2.33||||||2|4|3|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child: Graduated|62.1||1|1|3|4|F|Black||19||Mother|28208|Two Parent|$15,000 to $19,999||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||48|28214|Bachelors Degree|Single|Tech: Management|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Project Big|Enrollment|277|60|598|500000170|500017732|502537922|31|0|2|500189507|31|0|2|500535475|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2|500000294, 500004640|-2|0|4|||2238|7|||1|277756|-1|4|3|44
502469110|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-11|2014-03-03|Baseline|2011-05-09|2011-05-11|Complete|Done|3|3|3|2|4|3|3|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||2|5|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Moved|33.7||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||35|28269|Associate Degree|Married|Arts, Entertainment, Sports|28262|3|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502469557|31|0|1|502564995|31|0|1|500535534|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7496|10|||1|277903|-1|4|3|44
502206676|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-31|2011-10-25|Baseline|2011-05-10|2011-05-31|Complete|Done|3|2|2|1|3|3|2.33|||||||||3|3|3|3|2|3|2.83|||||||||4|4|4|4||||||3|2|3|2|2.5|||||||4|4|4|4|4|4||||||||||||4|4|4|4||||||3|3|3|||||2|2|||||||||Green|Amachi|Child: Severity of challenges|4.8||1|1|1|1|M|Black||18|Yes|Mother|28216|Other Relative|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|M|White||47|28269|Bachelors Degree|Married|Education: Teacher||7|0|Local Print|Media|Big|General Community|Amachi|RTBM|277|60|598|500000170|500011184|502207102|31|0|1|502562455|1|0|1|500535587|2||500003586||4|1|500000294|500000294, 500004640, 500004901|-2|500000294|-2|7016|11|||7439|1|||1|278234|-1|4|3|44
502469110|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-11|2014-03-03|Followup|2012-05-11|2012-05-07|Complete|Done|2|1|1|1|2|2|1.5|3|3|3|2|4|3|3|-50|3|4|2|1|3|2|2.5|2|4|3|2|2|3|2.67|-6.37|4|4|4|4|4|4|4|4|0|3|3|3|3|3|2|5|3|4|3.5|-14.29|4|4|4|3|4|4|4|3.86|4|4|4|4|4|4|3|3.86|0|3|4|4|3.67|4|4|4|4|-8.25|2|2|2|4|3|3.5|-42.86|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Moved|33.7||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||35|28269|Associate Degree|Married|Arts, Entertainment, Sports|28262|3|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502469557|31|0|1|502564995|31|0|1|500535534|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7496|10|||1|278955|277903|4|3|45
501919423|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-24|NaT|Followup|2012-03-24|2012-05-16|Declined|Late||||||||4|4|4|4|4|4|4|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||4|5|4|3|4||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|3|3.5||||1|1|||||||Green|Project Big||83.7||1|1|1|1|M|Multi-race (Black & Hispanic)||17|No|Mother|28214|One Parent: Female|Unknown||No|TV|Media|General Community|Project Big|Match Support|M|White||34|28164|Masters Degree||Finance|28210|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501919819|38|0|1|502034798|1|0|1|500442066|2||500004641||2|1|500004640|500004640|-2||-2|56|1|||7464|9|||1|278992|36152|4|1|45
502530688|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-16|2012-05-10|Baseline|2011-05-11|2011-11-16|Complete|Done|4|3|2|2|4|4|3.17|||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||3|2|4|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|2|2|||||1|1||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|5.8||2|2|3|3|M|Black||17||Mother|28210|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28277|Bachelors Degree|Married|Business||0|0|Michael Baisden|Media|Big|General Community||Match Support|277|60|598|500000170|500011746|502531141|31|0|1|502166996|31|0|1|500571794|2||-2||4|3||500005291|-2||-2|0|3|||11272|1|||1|279295|-1|4|3|44
502566108|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-24|2014-09-08|Baseline|2011-05-11|2011-05-24|Complete|Done|3|2|4|1|3|4|2.83|||||||||2|3|3|2|2|3|2.5|||||||||4|3|4|3.67||||||4|1|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|4|3.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|39.5||1|1|1|1|F|Hispanic||17|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||33|28209||Single|Student: College||0|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502566562|3|0|2|502562271|1|0|2|500535933|2||-2||4|1|500005291|500005291|-2|500005291|-2|0|4|||7464|9|||1|279328|-1|4|3|44
500783100|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-08-29|Followup|2012-04-30|2012-06-25|Complete|Late|4|4|4|4|4|4|4|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|3|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|||||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|112||1|1|1|1|M|Black||16||Mother|28206|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||36|28203|||Retail: Sales|28226|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|500783368|31|0|1|500777047|1|0|1|500174449|2||-2||4|2|||-2||-2|0|10|||46|2|||1|279659||4|3|45
500378354|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-01|NaT|Followup|2012-05-01|2012-06-19|Blank|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||106.5||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$40,000 to $44,999||No|Big|Neighbor/Friend|General Community||Match Support|M|White||36|28270|Juris Doctorate (JD)|Married|Law: Lawyer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500378596|31|0|1|501181060|1|0|1|500264206|2||-2||2|1|||-2||-2|6854|8|||46|2|||1|279661||4|3|45
501092911|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-01|2015-08-18|Followup|2013-05-01|2013-05-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|87.6||1|1|1|1|M|Black||19||Mother|28226|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|M|White||37|28210|Some College|Single|Business: Mgt, Admin||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|501064244|31|0|1|501176101|1|0|1|500261235|2||-2||4|3|||-2||-2|0|4|||46|2|||1|279662||4|1|45
501526673|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-25|2013-10-09|Followup|2013-02-25|2013-02-19|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|3|3|4|3|4|3.33|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|3|4|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|Amachi|Child: Lost interest|55.4||1|1|1|1|F|White||18|Yes||28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||34|28213|Bachelors Degree|Single|Real Estate: Realtor|28215|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500012459|501526965|1|0|2|501361484|1|0|2|500332705|2||500003586||4|2|500000294||-2||-2|0|10|||7496|10|||1|279776||4|3|45
501526664|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-25|2013-02-19|Followup|2012-02-25|2012-04-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Moved|47.8||1|1|1|1|F|White||15|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|F|White||35|28269|Bachelors Degree|Single|Business: Sales|33609|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|501526956|1|0|2|501233757|1|0|2|500332719|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7496|10|||1|279778||4|1|45
502490193|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-24|2013-01-09|Baseline|2011-05-12|2011-05-24|Complete|Done|3|3|2|3|3|3|2.83|||||||||3|3|3|3|3|3|3|||||||||4|3|3|3.33||||||3|3|4|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|19.6||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||40|28277|Masters Degree|Single|Medical: Pharmacist||0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500004169|502490640|31|0|1|502547160|1|0|1|500536146|2||-2||4|3|500005291|500005291|-2||-2|6854|8|||7496|10|||1|280209|-1|4|3|44
502185074|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-12|2016-08-02|Followup|2012-05-12|2012-06-29|Declined|Late||||||||1|2|1|4|1|1|1.67|||||||||3|1|3|1|1|1|1.67||||||4|4|4|4|||||||3|2|4|5|3.5||||||||||4|4|4|4|4|4|4|4||||||2|3|2|2.33|||||2|2|2||||2|2|||||||Green|2010-2012 OJJDP JJI|Child: Graduated|62.7||2|2|1|1|F|Black||18|No|GrandMother|28208|Grandparents|Unknown||Yes|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||68|28262|Bachelors Degree|Living w/ Significant Other|Business: Clerical||2|0|Relative|Relative|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017732|502185503|31|0|2|502490418|31|0|2|500533846|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|5635|9|||17161|11|||1|280250|159621|4|1|45
502551092|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-20|2015-10-29|Baseline|2011-05-12|2011-05-20|Complete|Done|3|3|4|1|4|4|3.17|||||||||2|4|3|1|2|4|2.67|||||||||4|4|4|4||||||3|4|5|3|3.75|||||||4|4|4|4|4|4|2|3.71||||||||||3|4|4|3.67||||||4|2|3|||||1|1||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|53.3||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||42|28210||Single|Business: Human Resources||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|502551545|31|0|2|502366844|1|0|2|500536172|2||-2||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||10326|3|460|3|1|280274|-1|4|3|44
500727291|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-17|2016-07-29|Followup|2012-05-17|2012-05-07|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|110.4||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|Black||46|28269|||Human Services: Non-Profit||0|0|BBBS National Site|Web Link|Big|General Community|VOL - Adjudicated, VOL - Cultural Comp, VOL - PreMatch|Match Support|277|60|598|500000170|500008321|500727558|31|0|1|500857838|31|0|1|500176403|2||-2||4|1|||-2|500007913, 500007920, 500011311|-2|0|10|||46|2|||1|280390||4|3|45
502537477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-12|2016-07-14|Followup|2012-05-12|2012-06-29|Declined|Late||||||||3|2|1|1|3|3|2.17|||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||3|5|4|4|4||||||||||4|4|4|4|3|4|3|3.71||||||2|3|2|2.33|||||2|4|3||||2|2||||4|4||Green|Project Big, 2010-2012 OJJDP JJI|Child: Graduated|62.1||1|1|3|4|F|Black||19||Mother|28208|Two Parent|$15,000 to $19,999||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||48|28214|Bachelors Degree|Single|Tech: Management|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Project Big|Enrollment|277|60|598|500000170|500017732|502537922|31|0|2|500189507|31|0|2|500535475|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2|500000294, 500004640|-2|0|4|||2238|7|||1|280463|277756|4|1|45
501390344|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-26|NaT|Followup|2012-02-26|2012-02-13|Complete|Done|4|2|2|2|2|3|2.5|||||||||1|3|4|1|2|3|2.33|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Amachi||96.6||1|1|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Single|Tech: Computer/Programmer||0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|501390617|31|0|1|501380163|1|0|1|500342682|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|280656||4|3|45
500185571|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-02|2015-07-14|Followup|2013-05-02|2013-05-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|110.4||1|1|1|1|M|Black||19||Mother|28215|Other/Unknown|Unknown||No|Other|Faith Organization|General Community||Match Support|M|Black||49|28213|Bachelors Degree|Married|Finance: Banking|28288|4|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187198|31|0|1|500188438|31|0|1|500089543|2||-2||4|3|||-2||-2|5635|9|||7464|9|||1|282556||4|1|45
500186141|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-02|2014-04-30|Followup|2012-04-02|2012-05-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|72.9||3|3|1|1|F|Black||20|No|Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||45|28269|Bachelors Degree|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|500187731|31|0|2|501046739|31|0|2|500254296|2||-2||4|1|||-2|500000294|-2|0|10|||46|2|||1|282588||4|1|45
502000252|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-22|NaT|Followup|2011-08-22|2011-08-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||78.8||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020910|502000651|31|0|1|502127058|1|0|1|500465318|2||-2||2|1|||-2||-2|0|10|||130|1|||1|282653||4|1|45
501716720|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-02|2017-02-06|Followup|2012-03-02|2012-05-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Cabarrus County|Child/Family: Lost contact with volunteer/agency|83.2||1|1|1|1|M|Black||15|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||52|28075||Married|Medical: Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501716992|31|0|1|501878786|31|0|1|500435676|2||500016307||4|3|500016374|500016374|-2|500016374|-2|6854|8|||7464|9|||1|282685||4|0|45
502242649|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-27|2012-05-09|Baseline|2011-05-17|2011-05-27|Complete|Done|4|1|2|1|2|3|2.17|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|4|2.5|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Moved|11.4||1|1|1|1|M|Hispanic|Dominican|17|No|Mother|28212|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|M|Hispanic||44|28211|Masters Degree|Married|Finance: Banking|28277|2|10|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502243080|3|13|1|502576783|3|0|1|500536543|2||-2||4|3|500005291|500005291|-2||-2|6854|8|||7462|13|||1|282768|-1|4|3|44
502402515|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-17|2015-12-28|Followup|2012-05-17|2012-07-02|Complete|Late|4|4|4|4|4|4|4|3|1|3|1|1|4|2.17|84.33|2|3|3|3|3|3|2.83|1|4|3|1|3|4|2.67|5.99|4|4|4|4|4|4|4|4|0|5|3|2|2|3|3|2|2|2|2.25|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|3|3|3|4|3|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|55.4||1|1|1|1|M|Black||16|No|Mother|28215|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28215||Single|Law: Police Officer||14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502402953|31|0|1|502537081|31|0|1|500535130|2||-2||4|1|500005291|500005291|-2||-2|34|2|||7464|9|||1|282908|276236|4|3|45
502549829|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-30|NaT|Baseline|2011-05-17|2011-06-30|Complete|Done|3|1|2|1|2|2|1.83|||||||||2|3|2|2|2|2|2.17|||||||||3|2|2|2.33||||||3|2|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Green|Amachi, Project Big, Project Big AND Amachi||68.5||1|1|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|Amachi, PERL 2014-2016, Project Big, Project Big AND Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Business: Engineer|30357|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|1|502594393|31|0|1|500541795|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901, 500014681|-1||-2|0|4|||7464|9|||1|283404|-1|4|3|44
501990745|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-14|2012-08-29|Followup|2012-05-14|2012-05-22|Declined|Done||||||||2|2|3|1|1|2|1.83|||||||||3|3|3|3|4|3|3.17||||||3|3|3|3|||||||5|4|3|5|4.25||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||4|4|4||||1|1|||||||Red||Child: Severity of challenges|27.5||1|1|1|1|M|Black||16||Mother|28269|One Parent: Female|Unknown||Yes||BBBS Board/Staff|General Community||Match Support|M|Black||35|28213||Married|Human Services: Youth Worker||0|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500011746|501991144|31|0|1|502098002|31|0|1|500447817|2||-2||4|3|||-2||-2|0|13|||4748|14|||1|283820|38490|4|1|45
502045254|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-08|2015-10-09|Followup|2012-06-08|2012-07-09|Declined|Done||||||||2|4|4|4|3|4|3.5|||||||||2|4|3|2|2|3|2.67||||||4|4|4|4|||||||2|4|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|3|2|3|||||3|3|3||||1|1|||||||Yellow||Child: Graduated|64||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502171015|31|0|2|500454926|2||-2||4|2|||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1|283829|134736|4|1|45
502590656|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2011-11-09|Baseline|2011-05-18|2011-06-30|Complete|Done|4|4|4|4|4|4|4|||||||||4|3|4|4|3|4|3.67|||||||||4|4|4|4||||||5|3|3|5|4|||||||4|2|4|4|4|4|3|3.57||||||||||4|4|4|4||||||4|3|3.5|||||1|1||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|4.3||1|1|1|1|F|Black||19|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|RTBM|F|Black||34|28262|Bachelors Degree|Single|Medical: Nurse|28262|1|6|TV|Media|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502591168|31|0|2|502578640|31|0|2|500538729|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||130|1|||1|284189|-1|4|3|44
502596391|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-12|2013-08-20|Baseline|2011-05-18|2011-06-12|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|4|3|4|4|3|3.5|||||||||4|2|2|2.67||||||2|3|5|3|3.25|||||||4|4|4|3|1|3|2|3||||||||||3|4|2|3||||||1|4|2.5|||||2|2||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|26.3||1|1|2|2|F|Black||16|No|Mother|28208|Two Mothers|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502596909|31|0|2|502485670|31|0|2|500540403|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7462|13|1204|3|1|284319|-1|4|3|44
500948129|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-18|2016-06-30|Followup|2012-03-18|2012-03-29|Complete|Done|4|2|4|2|3|4|3.17|||||||||3|4|4|4|1|4|3.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Child: Graduated|75.4||2|2|1|1|F|Black||18|No|Mother|28217|One Parent: Female|$25,000 to $29,999|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||40|28203|Some College|Living w/ Significant Other|Finance: Banking|28281|1|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501891556|1|0|2|500438403|2||500003586||4|1|500000294|500000294|-2||-2|34|2|||7464|9|||1|284744||4|3|45
501340097|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-23|2016-09-19|Followup|2012-03-23|2012-04-13|Complete|Done|3|4|4|2|4|3|3.33|||||||||2|2|3|3|2|3|2.5|||||||||3|2|4|3||||||2|5|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||2|2|2|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|77.9||2|2|1|1|M|Multi-race (Black & Hispanic)||17|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Hispanic||28|28277|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340376|38|0|1|501934966|3|0|1|500440292|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|284745||4|3|45
502569117|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-31|NaT|Baseline|2011-05-19|2011-05-26|Complete|Done|4|2|4|1|3|4|3|||||||||2|4|4|3|4|4|3.5|||||||||4|4|4|4||||||5|4|5|3|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|2|3||||||2|2|2|||||1|1||||4|4||||Green|Amachi, 2010-2012 OJJDP JJI||69.5||1|1|1|1|F|Black||15|Yes|Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||40|28269|Masters Degree|Single|Tech: Engineer|77058|6|6|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500017732|502569571|31|0|2|502538689|31|0|2|500536957|2||500003586||2|1|500000294, 500005291|500005291|-2||-2|0|10|||17161|11|||1|284793|-1|4|3|44
502495501|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-20|NaT|Followup|2012-05-20|2012-05-17|Complete|Done|3|2|3|1|1|2|2|3|1|4|2|2|2|2.33|-14.16|2|3|3|3|3|3|2.83|2|3|3|1|2|3|2.33|21.46|4|3|4|3.67|4|4|4|4|-8.25|5|3|3|4|3.75|5|3|2|3|3.25|15.38|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|3|3.71|4.04|4|4|3|3.67|4|4|3|3.67|0|3|1|2|2|1|1.5|33.33|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||69.9||1|1|1|1|M|White||15|No|Mother|28226|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||55|28210|Bachelors Degree|Married|Finance|28203|1|6|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500018851|502495950|1|0|1|502508181|1|0|1|500531873|2||-2||2|1|500005291|500005291|-2|500005291|-2|0|10|||7464|9|||1|285685|268809|4|3|45
502549826|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-13|2013-02-27|Baseline|2011-05-20|2011-06-13|Complete|Done|3|2|3|2|3|4|2.83|||||||||2|4|4|3|3|3|3.17|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|20.5||4|4|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||32|28209|Bachelors Degree|Single|Law: Paralegal|28204|1|5||Relative|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011349|502550279|31|0|2|502584664|1|0|2|500537198|2||500004772||4|3|500000294, 500004640, 500004901, 500005291|500014505, 500015184|-1|500004640|-2|0|4|||0|11|||1|285796|-1|4|3|44
502259046|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-25|2013-09-16|Baseline|2011-05-20|2011-05-25|Complete|Done|2|3|4|3|3|4|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1|||||||||Yellow||Volunteer: Time constraint|27.8||1|1|1|1|F|White||17|No|Mother|28025|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Enrollment|F|White||64|28083|High School Graduate|Married|Finance: Banking||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502259478|1|0|2|502502361|1|0|2|500537239|2||||4|2|||-2||-2|6854|8|||7464|9|||1|285946|-1|4|3|44
502551092|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-20|2015-10-29|Followup|2012-05-20|2012-06-11|Complete|Done|3|2|4|2|3|3|2.83|3|3|4|1|4|4|3.17|-10.73|2|3|3|3|2|3|2.67|2|4|3|1|2|4|2.67|0|4|4|4|4|4|4|4|4|0|3|3|2|4|3|3|4|5|3|3.75|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|||3|4|4|3.67||3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|53.3||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||42|28210||Single|Business: Human Resources||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|502551545|31|0|2|502366844|1|0|2|500536172|2||-2||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||10326|3|460|3|1|285955|280274|4|3|45
502552443|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-08|2014-12-30|Baseline|2011-05-20|2011-06-08|Complete|Done|4|4|4|2|3|4|3.5|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||2|2|2|||||||||||||||Green|Project Big|Child: Graduated|42.7||1|1|1|1|F|Multi-race (Black & Hispanic)||20|No|GrandMother|28208|Grandparents|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28209|Bachelors Degree|Single|Medical|28209|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502552891|38|0|2|502471967|1|0|2|500537261|2||-2||4|1|500004640|500004640, 500005291|-2||-2|0|4|||7496|10|||1|286064|-1|4|3|44
500724632|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-07|NaT|Followup|2012-03-07|2012-05-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||120.3||1|1|1|1|F|Black||17||Mother|28213|One Parent: Female|Less than $10,000|Y|No||School|General Community||Match Support|F|Black||32|28214|Bachelors Degree|Married|Architect|28270|0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|500724899|31|0|2|500803551|31|0|2|500164708|2||-2||2|1|||-2||-2|0|4|||46|2|||1|286396||4|0|45
502173445|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-23|2013-09-26|Followup|2012-05-23|2012-06-12|Complete|Done|4|4|4|1|4|4|3.5|4|4|4|3|4|4|3.83|-8.62|2|4|4|4|2|4|3.33|2|4|3|3|4|3|3.17|5.05|3|4|4|3.67|4|3|4|3.67|0|5|3|4|5|4.25|5|4|4|4|4.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|2|2|4|3|3.5|-42.86|2|2|2|2|0|4|4||||Red|Amachi|Volunteer: Lost contact with child/agency|28.2||1|1|1|1|F|Black||19|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Service Organization|General Community|Amachi|Match Support|F|White||28|28206|Bachelors Degree|Single|Education: Teacher||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502173869|31|0|2|502266833|1|0|2|500532710|2||500003586||4|3|500000294|500000294|-2||-2|0|11|||7464|9|||1|286615|270032|4|3|45
502566108|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-24|2014-09-08|Followup|2012-05-24|2012-06-13|Complete|Done|4|2|3|2|3|4|3|3|2|4|1|3|4|2.83|6.01|2|3|4|1|3|4|2.83|2|3|3|2|2|3|2.5|13.2|4|4|4|4|4|3|4|3.67|8.99|5|4|4|5|4.5|4|1|4|4|3.25|38.46|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3.67|8.99|2|3|2.5|3|4|3.5|-28.57|||1|1||4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|39.5||1|1|1|1|F|Hispanic||17|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||33|28209||Single|Student: College||0|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502566562|3|0|2|502562271|1|0|2|500535933|2||-2||4|1|500005291|500005291|-2|500005291|-2|0|4|||7464|9|||1|288039|279328|4|3|45
500903951|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-04|2013-02-26|Followup|2012-04-04|2012-05-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Lost interest|58.8||1|1|1|1|M|Black||21|Yes|Mother|28203|One Parent: Female|Less than $10,000|Y|No||Faith Organization|General Community|Amachi|Match Support|M|White||34|28202|Bachelors Degree|Single|Finance: Banking||3|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|500904221|31|0|1|501167853|1|0|1|500252953|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|288303||4|1|45
500185752|BBBS of Greater Charlotte|Main Office|C|Completed|2004-03-16|2012-10-17|Followup|2012-03-16|2012-05-01|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|103.1||1|2|1|2|M|Black||22|Yes|Mother|28227|One Parent: Female|Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||51|28212|Some College|Single|Clergy||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500012459|500187343|31|0|1|500188744|31|0|1|500038128|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|288306||4|1|45
502490193|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-24|2013-01-09|Followup|2012-05-24|2012-06-13|Complete|Done|3|2|2|2|3|3|2.5|3|3|2|3|3|3|2.83|-11.66|3|3|3|4|4|3|3.33|3|3|3|3|3|3|3|11|4|4|4|4|4|3|3|3.33|20.12|4|3|4|3|3.5|3|3|4|2|3|16.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|2|3|2.5|3|2|2.5|0|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|19.6||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||40|28277|Masters Degree|Single|Medical: Pharmacist||0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500004169|502490640|31|0|1|502547160|1|0|1|500536146|2||-2||4|3|500005291|500005291|-2||-2|6854|8|||7496|10|||1|288719|280209|4|3|45
501811395|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-10|NaT|Followup|2012-03-10|2012-02-07|Complete|Early|4|4|4|4|1|4|3.5|||||||||1|4|4|4|4|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|Cabarrus County||84.2||1|1|1|1|F|Black||15|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||60|28213||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501811730|31|0|2|500876892|31|0|2|500436702|2||500016307||2|1|500016374|500016374|-2|500016374|-2|6854|8|||2238|7|||1|289348||4|3|45
502241113|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-17|2012-06-28|Baseline|2011-05-25|2011-06-17|Complete|Done|3|1|4|4|2|4|3|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||2|4|4|3.33||||||2|2|2|||||1|1|||||||||Red||Child: Lost interest|12.4||1|1|2|2|F|Black||17|No|GrandMother|28025|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||43|28027|Masters Degree||Education: Teacher|28027|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|502241544|31|0|2|502460114|31|0|2|500538414|2||-2||4|3|||-2|500016374|-2|0|10|||7464|9|||1|289617|-1|4|3|44
502270499|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-25|NaT|Followup|2012-05-25|2012-06-06|Complete|Done|4|2|3|2|3|4|3|4|2|1|1|3|4|2.5|20|3|4|3|4|3|4|3.5|2|4|4|2|1|3|2.67|31.09|4|4|4|4|4|4|4|4|0|3|4|5|3|3.75|3|4|3|4|3.5|7.14|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|3|3|3|4|4|4|-25|2|2|2|2|0|4|4||||Green|Amachi||69.7||2|2|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||34|28203|Masters Degree|Single|Business: Mgt, Admin|28273|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502231230|31|0|2|502510107|1|0|2|500536754|2||500003586||2|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|289704|218599|4|3|45
500736177|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-25|2012-11-30|Followup|2012-05-25|2012-07-03|Complete|Done|3|2|3|2|3|3|2.67|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|18.2||2|3|1|1|F|Black||17||Mother|28269|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||38|28206|Bachelors Degree|Single|Finance|28255|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500710887|31|0|2|502513250|1|0|2|500536659|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|290237||4|3|45
502259046|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-25|2013-09-16|Followup|2012-05-25|2012-05-14|Complete|Done|4|4|4|4|4|4|4|2|3|4|3|3|4|3.17|26.18|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|5|5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|3|3|3|16.67|2|2|1|1|100|4|4||||Yellow||Volunteer: Time constraint|27.8||1|1|1|1|F|White||17|No|Mother|28025|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Enrollment|F|White||64|28083|High School Graduate|Married|Finance: Banking||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502259478|1|0|2|502502361|1|0|2|500537239|2||||4|2|||-2||-2|6854|8|||7464|9|||1|290397|285946|4|3|45
502589869|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2011-10-10|Baseline|2011-05-26|2011-06-30|Complete|Done|4|2|2|3|1|1|2.17|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|3|4|4|4|4|3|3.71||||||||||4|3|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|3.4||2|2|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||43|28262||Married|Medical: Nurse|28208|0|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502590381|31|0|2|501833131|31|0|2|500538612|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|290937|-1|4|3|44
502508499|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-06|2012-08-29|Baseline|2011-05-26|2011-06-06|Complete|Done|4|2|3|2|4|4|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|14.8||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|White||33|28209|Bachelors Degree|Single|Consultant||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502508948|31|0|2|502079235|1|0|2|500538672|2||-2||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||7496|10|||1|291168|-1|4|3|44
502551116|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2013-08-01|Baseline|2011-05-26|2011-06-30|Complete|Done|2|2|2|2|1|2|1.83|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||3|4|3.5|||||2|2||||4|4||||Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Moved|25.1||1|1|2|2|F|Hispanic||17|Yes|GrandFather|28216|One Parent: Male|$15,000 to $19,999||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black|Other African|36|28105||Single|Consultant|28244|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|502551569|3|0|2|500892262|31|31|2|500541956|2||500004772||4|2|500000294, 500004640, 500004901, 500005291|500004640, 500005291|-2||-2|0|4|||46|2|||1|291380|-1|4|3|44
502589865|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-29|Baseline|2011-05-26|2011-06-30|Complete|Done|1|4|2|3|1|1|2|||||||||3|1|3|4|4|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|1|1|||||2|2||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|52||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Black||40|28037|Bachelors Degree|Married|Medical: Doctor, Provider||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502590381|31|0|1|502625828|31|0|1|500544108|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|291589|-1|4|3|44
502567548|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-27|2012-10-31|Followup|2012-05-27|2012-07-11|Complete|Done|3|3|2|2|3|2|2.5|3|4|3|4|4|4|3.67|-31.88|2|4|3|2|3|3|2.83|4|4||4|4|4|||4|4|4|4|4|4|4|4|0|3|3|2|2|2.5|5|2|5|4|4|-37.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|4|4|4|4|-8.25|3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Red|Amachi, Project Big AND Amachi|Child/Family: Moved|17.2||1|1|2|2|F|Hispanic||16|Yes|Mother|28227|One Parent: Female|Unknown||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502568002|3|0|2|502564910|31|0|2|500534824|2||500003586||4|3|500000294, 500004901|500004640, 500004901|-2||-2|0|4|||17161|11|||1|291873|275240|4|3|45
502552438|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-02|2017-02-23|Baseline|2011-05-27|2011-06-02|Complete|Done|4|3|4|1|3|4|3.17|||||||||4|4|4|2|4|3|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|4|3|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|68.8||1|1|1|1|M|Black||16|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||36|28205|Masters Degree|Living w/ Significant Other|Journalist/Media|28202|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502552891|31|0|1|502549491|1|0|1|500538826|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||7464|9|||1|292098|-1|4|3|44
502008563|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-02|2013-07-29|Followup|2011-06-02|2011-06-14|Complete|Done|4|1|4|1|1|4|2.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green||Volunteer: Moved|37.9||2|2|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|28210|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502008962|31|0|1|502053340|1|0|1|500453826|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|292746||4|3|45
500824037|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-15|NaT|Followup|2012-03-15|2012-03-13|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4||4|4|4|||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||120||1|1|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|F|White||34|28210|Bachelors Degree|Single|Education: Teacher|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500824306|31|0|2|500789337|1|0|2|500165956|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|292930||4|3|45
502569117|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-31|NaT|Followup|2012-05-31|2012-06-26|Complete|Done|3|3|3|3|3|3|3|4|2|4|1|3|4|3|0|4|4|4|4|4|4|4|2|4|4|3|4|4|3.5|14.29|4|4|4|4|4|4|4|4|0|5|5|4|5|4.75|5|4|5|3|4.25|11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|3|2|3|33.33|4|4|4|2|2|2|100|2|2|1|1|100|4|4|4|4|0|Green|Amachi, 2010-2012 OJJDP JJI||69.5||1|1|1|1|F|Black||15|Yes|Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||40|28269|Masters Degree|Single|Tech: Engineer|77058|6|6|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500017732|502569571|31|0|2|502538689|31|0|2|500536957|2||500003586||2|1|500000294, 500005291|500005291|-2||-2|0|10|||17161|11|||1|293365|284793|4|3|45
502590651|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2013-08-22|Baseline|2011-05-31|2011-06-30|Complete|Done|4|3|4|2|4|4|3.5|||||||||2|4|3|1|2|4|2.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||4|3|3.5|||||1|1||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|25.8||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||36|28205|Bachelors Degree|Single|Business: Marketing|28117|7|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011746|502591168|31|0|2|502589724|1|0|2|500542166|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|294373|-1|4|3|44
502591898|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-04|2012-05-24|Baseline|2011-05-31|2011-06-04|Complete|Done|3|3|4|2|3|4|3.17|||||||||4|3|4|2|4|4|3.5|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Moved|11.7||2|2|1|1|F|Black||16|No|Mother|28214|Two Parent|$40,000 to $44,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||28|28202|Bachelors Degree|Single|Finance: Banking|28210|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502592415|31|0|2|502476195|1|0|2|500539115|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7496|10|||1|294647|-1|4|3|44
501212047|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-07|NaT|Followup|2012-05-07|2012-06-19|Complete|Done|4|3|3|2|4|4|3.33|||||||||2|4|3|3|4|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green|||106.3||1|1|1|1|F|White||18|No|Father|28207|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||33|28226||Single|Human Services: Non-Profit|28205|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501212321|1|0|2|501242250|1|0|2|500264889|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|294759||4|3|45
502045258|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-25|2016-08-29|Followup|2012-06-25|2012-07-02|Complete|Done|3|4|4|2|4|4|3.5|4|2|4|1|4|4|3.17|10.41|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|5|4|4.75|5|5|5|5|5|-5|4|3|4|4|4|4|3|3.71|4|4|4|4|4|4|3|3.86|-3.89|4|4|4|4|3|4|4|3.67|8.99|3|4|3.5|4|3|3.5|0|2|2|2|2|0|4|4||||Green||Volunteer: Lost contact with child/agency|74.2||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28262|Bachelors Degree|Single|Medical: Nurse|28262|4|9|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502190790|31|0|2|500457916|2||-2||4|1|||-2||-2|0|10|||6247|12|||1|296299|148107|4|3|45
502570396|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-08|Baseline|2011-06-01|2011-06-30|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|3|4|2|3|3.33|||||||||4|4|4|4||||||3|5|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|51.3||1|1|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28078|Bachelors Degree|Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018987|502570850|38|0|2|502545897|31|0|2|500539251|2||-2||4|1|500005291|500005291|-2||-2|34|2|||46|2|||1|296321|-1|4|3|44
502552438|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-02|2017-02-23|Followup|2012-06-02|2012-05-17|Complete|Early|3|3|3|1|3|3|2.67|4|3|4|1|3|4|3.17|-15.77|3|4|4|3|3|3|3.33|4|4|4|2|4|3|3.5|-4.86|4|4|4|4|4|4|4|4|0|5|4|4|5|4.5|5|4|4|5|4.5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|4|3.67|3|4|4|3.67|0|2|2|2|2|4|3|-33.33|2|2|2|2|0|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|68.8||1|1|1|1|M|Black||16|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||36|28205|Masters Degree|Living w/ Significant Other|Journalist/Media|28202|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502552891|31|0|1|502549491|1|0|1|500538826|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||7464|9|||1|297947|292098|4|3|45
502528773|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-16|2012-05-30|Baseline|2011-06-03|2011-06-15|Complete|Done|4|4|3|4|4|4|3.83|||||||||2|4|3|3|3|4|3.17|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|2|2|2.33||||||3|4|3.5|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Moved|11.5||1|1|1|1|F|Hispanic|Mexican|18|No|Mother|28215|One Parent: Female|Unknown||No|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||36|28262|Masters Degree|Single|Finance|28273|3|10|BBBS National Site|Web Link|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500011746|502529226|3|10|2|502552143|3|0|2|500539575|2||-2||4|3|500005291|500005291|-2|500005291|-2|2203|12|||46|2|||1|298818|-1|4|3|44
502591943|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-29|2012-08-30|Baseline|2011-06-03|2012-01-29|Complete|Done|4|2|2|1|3|3|2.5|||||||||2|2|3|1|2|3|2.17|||||||||3|2|2|2.33||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Red||Child: Family structure changed|7||1|1|1|1|F|White||17|No|Mother|28278|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28209|Bachelors Degree|Single|Business: Mgt, Admin|28210|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502592460|1|0|2|502757658|1|0|2|500593218|2||||4|3||500005291|-2||-2|0|4|||7496|10|||1|298866|-1|4|3|44
500361200|BBBS of Greater Charlotte|Main Office|C|Active|2006-03-21|NaT|Followup|2012-03-21|2012-04-23|Complete|Done|2|2|2|3|1|3|2.17|||||||||2|1|3|1|3|3|2.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|4|3|||||2|2||||4|4||||Green|Cabarrus County||131.8||2|2|1|1|F|White||17|No|Mother|28027|Two Parent|Unknown||No||Relative|General Community|Cabarrus County|Match Support|F|White||32|28115|Bachelors Degree|Single|Human Services: Social Worker||0|0|other|College Partner|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500361450|1|0|2|500368628|1|0|2|500085591|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|3|||7670|5|||1|299427||4|3|45
500408135|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-25|2015-01-30|Followup|2012-05-25|2012-07-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|104.2||1|1|4|4|F|Black||19|Yes|Mother|28083|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500008321|500408385|31|0|2|500189709|31|0|2|500099932|2||500003586||4|1|500000294|500000294|-2|500000294, 500016374|-2|6854|8|||2230|7|||1|299538||4|1|45
502508499|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-06|2012-08-29|Followup|2012-06-06|2012-05-03|Complete|Early|3|2|4|4|4|4|3.5|4|2|3|2|4|4|3.17|10.41|3|4|4|3|3|4|3.5|4|4|4|4|4|4|4|-12.5|4|4|4|4|4|4|4|4|0|4|4|5|4|4.25|5|3|5|5|4.5|-5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|4|3.67|4|4|3|3.67|0|2|4|3|1|4|2.5|20|1|1|2|2|-50|4|4|4|4|0|Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|14.8||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|White||33|28209|Bachelors Degree|Single|Consultant||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502508948|31|0|2|502079235|1|0|2|500538672|2||-2||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||7496|10|||1|300199|291168|4|3|45
502597596|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-04-11|Baseline|2011-06-06|2011-06-30|Complete|Done|3|3|3|2|4|3|3|||||||||3|4|3|4|3|4|3.5|||||||||3|3|3|3||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||1|1||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Moved|9.4||1|1|1|1|F|Black||15||Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28273|Bachelors Degree|Single|Medical|28277|2|9|Self|Self|Big|General Site||RTBM|277|60|598|500000170|500013709|502598113|31|0|2|502560341|31|0|2|500540008|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2||-1|0|4|||7464|9|||1|300353|-1|4|3|44
502552443|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-08|2014-12-30|Followup|2012-06-08|2012-06-27|Complete|Done|4|4|4|4|4|4|4|4|4|4|2|3|4|3.5|14.29|2|4|4|4|4|4|3.67|4|4|4|4|2|4|3.67|0|4|4|4|4|4|4|4|4|0|5|4|3|4|4|5|4|4|5|4.5|-11.11|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|3|4|4|3.67|3|4|3|3.33|10.21|4|4|4|2|2|2|100|2|2||||4|4||||Green|Project Big|Child: Graduated|42.7||1|1|1|1|F|Multi-race (Black & Hispanic)||20|No|GrandMother|28208|Grandparents|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28209|Bachelors Degree|Single|Medical|28209|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502552891|38|0|2|502471967|1|0|2|500537261|2||-2||4|1|500004640|500004640, 500005291|-2||-2|0|4|||7496|10|||1|301988|286064|4|3|45
501160887|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2013-05-14|Followup|2012-04-30|2012-04-30|Complete|Done|4|3|3|1|4|4|3.17|||||||||3|3|4|4|3|4|3.5|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|36.5||2|2|1|1|F|Black||14|Yes|Mother|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Enrollment|F|White||58|28226|||Education: Teacher Asst/Aid|28203|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|501615415|1|0|2|500447312|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|302630||4|3|45
500799303|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-27|2016-08-19|Followup|2012-03-27|2012-04-23|Complete|Done|3|1|4|2|2|3|2.5|||||||||2|4|4|4|3|4|3.5|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|4|3.5|||||2|2||||4|4||||Red||Child: Graduated|112.8||1|1|1|1|M|White||19|No|Mother|28081|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||46|28202||Single|Business: Sales||0|4|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500799571|1|0|1|500798390|1|0|1|500167062|2||-2||4|3||500016374|-2|500016374|-2|34|2|||7464|9|||1|304490||4|3|45
501987736|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-29|2014-06-18|Followup|2012-06-29|2012-08-23|Blank|Late||||||||4|4|4|2|4|4|3.67|||||||||2|4|4|2|4|4|3.33||||||4|2|2|2.67|||||||4|3|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|1|1.5||||1|1|||||||Green||Child: Graduated|47.6||1|1|1|1|F|White||20|No|Father|28217|One Parent: Male|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||40|28203|Masters Degree|Single|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501988135|1|0|2|502109789|1|0|2|500456045|2||-2||4|1|||-2||-2|6855|8|||7464|9|||1|304709|142908|4|3|45
502596391|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-12|2013-08-20|Followup|2012-06-12|2012-05-07|Complete|Early|3|4|4|4|3|4|3.67|3|4|4|4|4|4|3.83|-4.18|2|4|4|3|2|3|3|3|4|3|4|4|3|3.5|-14.29|3|2|4|3|4|2|2|2.67|12.36|5|2|1|1|2.25|2|3|5|3|3.25|-30.77|4|4|4|4|4|4|3|3.86|4|4|4|3|1|3|2|3|28.67|3|4|3|3.33|3|4|2|3|11|1|2|1.5|1|4|2.5|-40|2|2|2|2|0|4|4|4|4|0|Yellow|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|26.3||1|1|2|2|F|Black||16|No|Mother|28208|Two Mothers|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502596909|31|0|2|502485670|31|0|2|500540403|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7462|13|1204|3|1|304801|284319|4|3|45
502549826|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-13|2013-02-27|Followup|2012-06-13|2012-07-02|Complete|Done|4|2|1|1|2|4|2.33|3|2|3|2|3|4|2.83|-17.67|1|2|3|3|4|3|2.67|2|4|4|3|3|3|3.17|-15.77|4|4|4|4|4|4|4|4|0|4|4|5|4|4.25|3|3|3|3|3|41.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|4|4|3.67|-9.26|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Red|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|20.5||4|4|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||32|28209|Bachelors Degree|Single|Law: Paralegal|28204|1|5||Relative|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011349|502550279|31|0|2|502584664|1|0|2|500537198|2||500004772||4|3|500000294, 500004640, 500004901, 500005291|500014505, 500015184|-1|500004640|-2|0|4|||0|11|||1|304966|285796|4|3|45
501626226|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-30|2017-03-14|Followup|2012-06-30|2012-06-18|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|3|3|3|4|3|3|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green||Child: Graduated|80.5||2|2|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||33|28203|High School Graduate|Single|Retail: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501622822|31|0|2|502036832|1|0|2|500457771|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|305233||4|3|45
502008563|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-02|2013-07-29|Followup|2012-06-02|2012-06-08|Complete|Done|4|3|2|2|3|3|2.83|||||||||4|3|4|4|3|4|3.67|||||||||3|3|3|3||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|37.9||2|2|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|28210|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502008962|31|0|1|502053340|1|0|1|500453826|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|305837||4|3|45
501631140|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-17|2016-03-03|Followup|2012-06-17|2012-08-10|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|80.5||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Service: Hotel|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501631463|31|0|1|501628976|1|0|1|500367187|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|305859||4|1|45
502581328|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-28|2015-07-27|Baseline|2011-06-14|2013-02-27|Complete|Done|3|2|3|2|1|3|2.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Yellow||Child: Lost interest|28.9||1|1|1|1|F|Black||16|No|GrandMother|28212|One Parent: Female|$20,000 to $24,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||46|28262|PHD|Single|Education: College Professor|28223|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502581832|31|0|2|503144090|31|0|2|500681651|2||-2||4|2|||-2||-2|6854|8|||7464|9|||1|306034|-1|4|3|44
502544191|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-21|2014-01-06|Baseline|2011-06-14|2011-06-19|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||1|1|||||||||Green|Amachi|Volunteer: Lost contact with child/agency|30.6||1|1|2|2|F|Black||20|Yes|Mother|28277|One Parent: Female|$50,000 to $59,999||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||29|28277|Bachelors Degree|Single|Consultant|28204|0|11|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502544644|31|0|2|502231024|1|0|2|500541173|2||-2||4|1|500000294|500000294|-2|500000294|-2|34|2|||46|2|||1|306127|-1|4|3|44
501599416|BBBS of Greater Charlotte|Main Office|C|Active|2009-04-28|NaT|Followup|2012-04-28|2012-05-31|Complete|Done|4|4|4|2|2|4|3.33|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||94.6||1|1|1|1|M|White||14|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||46|28078|Masters Degree|Single|Retail: Mgt|28207|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501599736|1|0|1|500188567|1|0|1|500357914|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|306145||4|3|45
500271303|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-30|2015-08-03|Followup|2012-04-30|2012-06-18|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|75.1||2|2|1|1|F|Black||17|Yes|Mother|28227|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|White||31|28204|Bachelors Degree|Single|Business: Engineer|28269|0|2|TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500271368|31|0|2|501291358|1|0|2|500354049|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||130|1|||1|306147||4|1|45
501074345|BBBS of Greater Charlotte|Main Office|C|Active|2008-03-31|NaT|Followup|2012-03-31|2012-04-23|Complete|Done|3|1|4|1|4|4|2.83|||||||||1|2|1|2|2|3|1.83|||||||||4|4|4|4||||||3|3|2|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Green|Amachi, Cabarrus County||107.5||1|1|1|1|M|White||16|Yes|GrandMother|28025|Grandparents|Unknown||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|White||46|28027|Bachelors Degree|Divorced|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501074618|1|0|1|501158523|1|0|1|500250038|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|5635|9|||46|2|||1|306521||4|3|45
502527850|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-10-04|Baseline|2011-06-15|2011-06-30|Complete|Done|3|3|4|3|3|3|3.17|||||||||2|3|2|2|3|3|2.5|||||||||4|4|4|4||||||3|1|3|4|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|3|3||||||4|4|4|||||2|2||||4|4||||Yellow|2010-2012 OJJDP JJI|Child: Lost interest|15.2||1|1|2|2|F|Black||19|No|Mother|28027|One Parent: Female|Less than $10,000||Yes|Brochure|Media|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||42|28213|Bachelors Degree|Single|Finance: Banking|28202|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|502528298|31|0|2|502598777|31|0|2|500541242|2||-2||4|2|500005291|500005291|-2|500016374|-2|51|1|||7464|9|||1|306634|-1|4|3|44
502482642|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-22|2012-07-31|Baseline|2011-06-15|2011-06-22|Complete|Done|3|3|4|3|3|3|3.17|||||||||3|3|3|4|2|3|3|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|13.3||2|2|1|1|F|Black||16|No|Mother|28052|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28204|Masters Degree|Single|Finance: Auditor|28202|2|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502391834|31|0|2|502601273|1|0|2|500541388|2||-2||4|3|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|10|||7496|10|||1|307140|-1|4|3|44
500185778|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-17|2016-06-23|Followup|2012-06-17|2012-08-10|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|144.2||1|1|1|1|M|Black||18||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||42|27514||Married|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187368|31|0|1|500188776|1|0|1|500036776|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|307582||4|1|45
502489575|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-08-29|Baseline|2011-06-16|2011-06-30|Complete|Done|4|2|3|1|4|4|3|||||||||3|4|3|3|4|3|3.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|14||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||44|28105|Masters Degree|Married|Business: Mgt, Admin|28202|3|6|Ally Financial|Workplace Partner|Big|General Site||RTBM|277|60|598|500000170|500011746|502490022|31|0|1|502432606|31|0|1|500541789|2||-2||4|3|500004640, 500005291|500005291|-2||-1|56|1|||12831|3|1209, 635|1|1|307800|-1|4|3|44
502241113|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-17|2012-06-28|Followup|2012-06-17|2012-06-28|Declined|Done||||||||3|1|4|4|2|4|3|||||||||3|4|4|4|4|4|3.83||||||4|4|4|4|||||||5|4|4|4|4.25||||||||||4|4|4|4|4|4|4|4||||||2|4|4|3.33|||||2|2|2||||1|1|||||||Red||Child: Lost interest|12.4||1|1|2|2|F|Black||17|No|GrandMother|28025|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||43|28027|Masters Degree||Education: Teacher|28027|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|502241544|31|0|2|502460114|31|0|2|500538414|2||-2||4|3|||-2|500016374|-2|0|10|||7464|9|||1|308098|289617|4|1|45
500186645|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-03|2016-01-06|Followup|2012-06-03|2012-06-10|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|139.1||1|1|1|1|M|Black||18|Yes|Mother|28208|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28256|High School Graduate|Married|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500018987|500188043|31|0|1|500189545|31|0|2|500037636|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|308105||4|1|45
502549784|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-29|2013-06-06|Baseline|2011-06-17|2011-06-29|Complete|Done|4|4|4|3|3|3|3.5|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||3|2|4|3|3|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|23.3||1|1|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|$20,000 to $24,999||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||30|28227||Single|Transport: Driver||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500011746|502550237|31|0|1|502558315|31|0|1|500541875|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|10|||7496|10|||1|308122|-1|4|3|44
502142541|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-18|2015-07-23|Followup|2012-06-18|2012-08-07|Declined|Late||||||||3|4|4|3|4|4|3.67|||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||4|4|5|3|4||||||||||4|4|4|4|3|4|3|3.71||||||4|4|4|4|||||2|2|2||||2|2|||||||Green||Child: Graduated|61.1||1|1|2|2|F|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502142970|31|0|2|501905673|31|0|2|500455759|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|308353|141478|4|1|45
502076679|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2012-09-06|Followup|2012-04-30|2012-07-15|Expired|Late||||||||4|2|3|2|3|4|3|||||||||3|3||3|3|3|||||||3|3|3|3|||||||2|4|4|4|3.5||||||||||4|4|4|4||4|4|||||||4|4|4|4|||||3|3|3||||2|2|||||||Red||Volunteer: Time constraint|28.3||1|1|1|1|M|Black||17|No|Mother|28273|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||37|28278|||Finance: Banking||0|0|AA Task Force|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502077103|31|0|1|502003579|1|0|1|500446859|2||-2||4|3|||-2||-2|0|4|||9228|10|||1|308358|38100|4|0|45
500956242|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-14|2013-02-28|Followup|2012-04-14|2012-05-21|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Moved|58.5||1|1|2|2|M|Multi-Race (None of the above)||19|No|Mother|28210|One Parent: Female|$20,000 to $24,999||Yes||Therapist/Counselor|General Community||Match Support|M|White||38|28210|||Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500956512|7|0|1|500189847|1|0|1|500259433|2||-2||4|3|||-2||-2|0|5|||7464|9|||1|308585||4|1|45
502581751|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2014-05-08|Baseline|2011-06-20|2011-06-27|Complete|Done|2|3|4|2|4|4|3.17|||||||||1|3|3|4|2|3|2.67|||||||||4|4|4|4||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Moved|34.4||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Black||38|28206|Masters Degree|Single|Business: Human Resources|28255|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502582259|31|0|1|502587677|31|0|1|500542041|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|308841|-1|4|3|44
502544191|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-21|2014-01-06|Followup|2012-06-21|2012-09-05|Expired|Late||||||||3|3|4|3|3|4|3.33|||||||||3|4|4|3|3|3|3.33||||||4|4|4|4|||||||5|5|4|4|4.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|2|2.5||||1|1|||||||Green|Amachi|Volunteer: Lost contact with child/agency|30.6||1|1|2|2|F|Black||20|Yes|Mother|28277|One Parent: Female|$50,000 to $59,999||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||29|28277|Bachelors Degree|Single|Consultant|28204|0|11|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502544644|31|0|2|502231024|1|0|2|500541173|2||-2||4|1|500000294|500000294|-2|500000294|-2|34|2|||46|2|||1|309330|306127|4|0|45
502545735|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-12|2012-06-22|Baseline|2011-06-21|2011-07-12|Complete|Done|4|2|4|2|1|4|2.83|||||||||2|3|3|3|2|4|2.83|||||||||4|4|4|4||||||2|5|1|5|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||1|3|2|||||2|2|||||||||Red||Volunteer: Health|11.4||1|1|1|1|M|Multi-race (Hispanic & White)||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||No|Big|Neighbor/Friend|General Community||RTBM|M|White||41|28205|Bachelors Degree|Married|Finance|28255|9|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502546188|35|0|1|502388739|1|0|1|500542256|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|309494|-1|4|3|44
502482642|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-22|2012-07-31|Followup|2012-06-22|2012-07-31|Declined|Done||||||||3|3|4|3|3|3|3.17|||||||||3|3|3|4|2|3|3||||||4|4|4|4|||||||3|4|4|4|3.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|2|2.5||||2|2||||4|4||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|13.3||2|2|1|1|F|Black||16|No|Mother|28052|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28204|Masters Degree|Single|Finance: Auditor|28202|2|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502391834|31|0|2|502601273|1|0|2|500541388|2||-2||4|3|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|10|||7496|10|||1|309919|307140|4|1|45
502510347|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-31|2016-08-30|Baseline|2011-06-22|2011-10-28|Complete|Done|4|1|2|1|4|4|2.67|||||||||1|4|2|2|2|2|2.17|||||||||4|4|4|4||||||3|4|2|4|3.25|||||||4|4|4|4|4|4|2|3.71||||||||||3|2|1|2||||||4|2|3|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child: Graduated|58||1|1|1|1|F|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28262|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502510796|31|0|2|502677833|31|0|2|500557844|2||-2||4|1|500005291|500005291|-2||-2|0|5|||7464|9|||1|310349|-1|4|3|44
501174643|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-06|2012-11-08|Followup|2012-05-06|2012-06-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|42.1||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|Black||34|28214||Married|Business: Sales|28210|0|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011349|501174917|31|0|1|501687908|31|0|1|500358149|2||-2||4|3|||-2||-2|0|10|||7446|3|||1|310539||4|1|45
502583109|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-26|2012-09-06|Baseline|2011-06-23|2011-10-26|Complete|Done|3|4|3|2|1|3|2.67|||||||||2|2|2|3|2|2|2.17|||||||||4|4|3|3.67||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||2|3|2|2.33||||||3|3|3|||||1|1||||4|4||||Green|Amachi|Child: Lost interest|10.4||1|1|2|2|F|Black||17|Yes|Mother|28277|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|Amachi|Match Support|F|White||39|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28217|1|7|Radio|Media|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008629|502583617|31|0|2|502236275|1|0|2|500551832|2||-2||4|1|500000294|500000294|-2|500000294|-2|0|10|||131|1|||1|310826|-1|4|3|44
501561529|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-11|2012-08-29|Followup|2012-05-11|2012-06-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|39.6||1|1|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||36|28202|Masters Degree|Single|Business: Sales|28202|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008629|501561821|31|0|1|501333443|1|0|1|500359635|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|311523||4|1|45
500961015|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-11|2014-10-02|Followup|2012-04-11|2012-04-16|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|2|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|77.7||1|1|1|1|M|Black||20|Yes|Mother|28227|Two Parent|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||43|28104||Married|Tech: Computer/Programmer|29607|10|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500013781|500934638|31|0|1|501210561|31|0|1|500257073|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||17161|11|||1|311571||4|3|45
501611456|BBBS of Greater Charlotte|Main Office|C|Active|2010-05-28|NaT|Followup|2012-05-28|2012-07-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||81.6||1|1|1|1|M|Black||15|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black|Other African|32|28262||Married|Law: Police Officer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501611776|31|0|1|501876475|31|31|1|500450969|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|311772||4|1|45
502581751|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2014-05-08|Followup|2013-06-27|2013-09-11|Expired|Late||||||||2|3|4|2|4|4|3.17|||||||||1|3|3|4|2|3|2.67||||||4|4|4|4|||||||3|2|4|4|3.25||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||3|3|3||||2|2|||||||Yellow||Volunteer: Moved|34.4||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Black||38|28206|Masters Degree|Single|Business: Human Resources|28255|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502582259|31|0|1|502587677|31|0|1|500542041|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|311872|308841|4|0|45
501842678|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2015-06-19|Followup|2012-06-27|2012-09-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Feels incompatible with child/family|47.7||2|2|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|White||53|28117|Bachelors Degree|Married|Real Estate: Realtor|28031|0|0|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|277|60|598|500000170|500015820|501843047|31|0|1|502335257|1|0|1|500542227|2||-2||4|2|||-2|500000294, 500004901|-2|0|10|||7464|9|||1|311980||4|0|45
500767208|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-03-24|Followup|2012-07-10|2012-09-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Child: Graduated|68.4||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|Black||32|28216|Masters Degree|Single|Human Services|28215|0|7|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Enrollment|277|60|598|500000170|500017732|500767473|31|0|2|501341042|31|0|2|500276669|2||500004641||4|1|500004640||-2|500014506|-1|0|10|||7671|13|||1|312260||4|1|45
500185534|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-13|2012-12-20|Followup|2012-05-13|2012-06-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Family structure changed|79.3||1|1|3|5|M|Black||18||Mother|28204|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||63|28206|Some College|Married|Self-Employed, Entrepreneur|28206|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187159|31|0|1|500189461|31|0|1|500093294|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|312308||4|1|45
500740293|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2012-06-12|2012-06-06|Complete|Done|1|4|3|3|3|4|3|||||||||1|4|4|1|4|3|2.83|||||||||4|4|4|4||||||5|3|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Yellow||Child: Lost interest|85||1|1|1|1|M|Black||19||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|Black||39|28216||Single|Transport: Pilot||3|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500876177|31|0|1|500179697|2||-2||4|2|||-2||-2|0|5|||6450|12|||1|312853||4|3|45
502646551|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-07-03|Baseline|2011-06-29|2011-06-30|Complete|Done|4|3|4|3|3|3|3.33|||||||||2|3|3|3|3|3|2.83|||||||||4|3|3|3.33||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|2|2.5|||||1|1||||4|4||||Green|Project Big|Child/Family: Moved|12.1||1|1|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|White||34|28210|High School Graduate|Single|Business: Sales|28269|0|8|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502598113|31|0|2|502262622|1|0|2|500543369|2||500004641||4|1|500004640|500004640|-2|500004640|-2|0|10|||7464|9|||1|312938|-1|4|3|44
502646565|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2011-10-04|Baseline|2011-06-29|2011-06-30|Complete|Done|4|3|4|2|4|4|3.5|||||||||2|4|2|2|2|3|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|2|2.5|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|3.2||1|1|2|2|M|Black||20|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|277|60|598|500000170|500008321|502598113|31|0|1|502528355|1|0|1|500543433|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||132|8|||1|313112|-1|4|3|44
502645489|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-07-03|Baseline|2011-06-29|2011-06-30|Complete|Done|4|4|4|3|4|3|3.67|||||||||3|4|3|3|3|3|3.17|||||||||4|3|3|3.33||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Child/Family: Moved|12.1||1|1|1|1|F|Black||20||Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||43|28214|Masters Degree|Married|Arts, Entertainment, Sports|28202|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502508948|31|0|2|502480739|31|0|2|500543463|2||500004641||4|1|500004640|500004640, 500005291|-2||-2|0|4|||7464|9|||1|313195|-1|4|3|44
502549784|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-29|2013-06-06|Followup|2012-06-29|2012-06-28|Complete|Done|4|4|4|1|4|3|3.33|4|4|4|3|3|3|3.5|-4.86|2|4|4|1|3|4|3|2|4|3|2|3|3|2.83|6.01|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|3|2|4|3|3|8.33|3|4|4|4|4|4|4|3.86|4|4|4|4|3|4|4|3.86|0|4|4|4|4|4|4|4|4|0|4|3|3.5|3|2|2.5|40|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|23.3||1|1|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|$20,000 to $24,999||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||30|28227||Single|Transport: Driver||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500011746|502550237|31|0|1|502558315|31|0|1|500541875|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|10|||7496|10|||1|313214|308122|4|3|45
501069450|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-07|2017-02-28|Followup|2011-11-07|2012-01-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|111.7||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||66|28075||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501048131|31|0|1|500887364|31|0|1|500212043|2||-2||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|313558||4|0|45
502589865|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-29|Followup|2012-06-30|2012-06-04|Complete|Early|3|3|3|3|2|4|3|1|4|2|3|1|1|2|50|4|4|4|2|2|4|3.33|3|1|3|4|4|4|3.17|5.05|4|3|3|3.33|4|4|4|4|-16.75|3|3|3|3|3|5|5|5|5|5|-40|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|3|3.33|20.12|3|4|3.5|1|1|1|250|2|2|2|2|0|4|4|4|4|0|Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|52||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Black||40|28037|Bachelors Degree|Married|Medical: Doctor, Provider||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502590381|31|0|1|502625828|31|0|1|500544108|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|313939|291589|4|3|45
500814240|BBBS of Greater Charlotte|Main Office|C|Active|2008-04-24|NaT|Followup|2012-04-24|2012-04-30|Complete|Done|3|3|3|1|4|3|2.83|||||||||2|4|4|3|3|4|3.33|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi||106.7||1|1|1|1|M|Black||18|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||46|28215|Bachelors Degree|Single|Business: Mgt, Admin|28226|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500814509|31|0|1|500981509|31|0|1|500248568|2||500003586||2|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|313998||4|3|45
501402710|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-19|2015-06-17|Followup|2012-06-19|2012-07-23|Complete|Done|3|2|3|2|3|3|2.67|||||||||2|3|3|2|1|2|2.17|||||||||4|4|4|4||||||2|5|5|3|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||3|3|2|2.67||||||3|3|3|||||2|2||||4|4||||Green||Child/Family: Moved|71.9||1|1|1|1|M|Black||18|No|Mother|30058|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28215||Married|Consultant|28285|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501402995|31|0|1|501728845|1|0|1|500368860|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|314002||4|3|45
500545470|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-01-25|Followup|2012-04-30|2012-06-15|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|104.9||1|1|1|1|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||34|29708|Bachelors Degree|Single|Self-Employed, Entrepreneur|29708|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501750989|31|0|1|500815012|1|0|1|500173957|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|3|||2238|7|||1|314086||4|1|45
500418050|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-12|2012-11-28|Followup|2012-05-12|2012-07-19|Complete|Late|4|4|4|1|4|4|3.5|||||||||2|2|3|4|2|3|2.67|||||||||4|4|4|4||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|3|2.5|||||1|1||||4|4||||Green|Amachi|Volunteer: Lost contact with child/agency|78.6||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||34|28273|High School Graduate|Single|Transport: Driver|28216|0|10|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188055|31|0|1|500417272|31|0|1|500093386|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|314096||4|3|45
500186955|BBBS of Greater Charlotte|Main Office|C|Completed|2004-05-21|2014-02-19|Followup|2012-05-21|2012-05-31|Complete|Done|4|4|4|4|4|3|3.83|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Lost contact with child/agency|117||1|1|1|1|F|Black||18|No|Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||55|28226|||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|2|500189726|1|0|2|500037840|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|314097||4|3|45
500363212|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-24|2012-11-27|Followup|2012-05-24|2012-07-03|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Volunteer: Moved|66.2||2|2|1|1|F|Multi-Race (None of the above)||16||Mother|28025|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||34|28211|Associate Degree|Living w/ Significant Other|Business: Clerical|28211|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188099|7|0|2|500797130|1|0|2|500176231|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|314100||4|3|45
500186953|BBBS of Greater Charlotte|Main Office|C|Completed|2004-05-25|2012-08-09|Followup|2012-05-25|2012-07-19|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.5||1|1|2|2|M|Black||18|Yes|GrandMother|28214|Other Relative|Unknown||No||Self|General Community|Amachi|Match Support|M|White||45|28207||Single|Unknown|28209|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188126|31|0|1|500189724|1|0|1|500037838|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|314103||4|1|45
501212662|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-23|2013-04-22|Followup|2012-06-23|2012-08-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|58||1|1|1|1|M|Multi-Race (None of the above)||16|Yes|Mother|28211|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Multi-Race (None of the above)||34|28205|Bachelors Degree|Single|Business: Sales|28210|0|10|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501212937|7|0|1|501252394|7|0|1|500269647|2||-2||4|3|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|314104||4|1|45
502570396|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-08|Followup|2012-06-30|2012-06-19|Complete|Done|4|1|4|4|4|4|3.5|3|4|4|4|4|4|3.83|-8.62|3|3|4|3|3|4|3.33|4|4|3|4|2|3|3.33|0|4|4|4|4|4|4|4|4|0|3|3|5|4|3.75|3|5|3|3|3.5|7.14|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|1|3|2|50|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|51.3||1|1|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28078|Bachelors Degree|Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018987|502570850|38|0|2|502545897|31|0|2|500539251|2||-2||4|1|500005291|500005291|-2||-2|34|2|||46|2|||1|314319|296321|4|3|45
502527850|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-10-04|Followup|2012-06-30|2012-06-01|Complete|Early|4|4|4|4|4|4|4|3|3|4|3|3|3|3.17|26.18|2|4|3|4|4|4|3.5|2|3|2|2|3|3|2.5|40|3|3|3|3|4|4|4|4|-25|3|4|4|4|3.75|3|1|3|4|2.75|36.36|4|4|4|4|4|3|3|3.71|4|4|4|4|4|4|3|3.86|-3.89|4|4|3|3.67|2|4|3|3|22.33|1|2|1.5|4|4|4|-62.5|1|1|2|2|-50|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Child: Lost interest|15.2||1|1|2|2|F|Black||19|No|Mother|28027|One Parent: Female|Less than $10,000||Yes|Brochure|Media|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||42|28213|Bachelors Degree|Single|Finance: Banking|28202|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|502528298|31|0|2|502598777|31|0|2|500541242|2||-2||4|2|500005291|500005291|-2|500016374|-2|51|1|||7464|9|||1|314358|306634|4|3|45
502180719|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-04|2014-03-20|Followup|2012-06-04|2012-05-31|Complete|Done|4|4|4|4|4|4|4|4|2|4|4|4|4|3.67|8.99|2|4|4|2|2|4|3|2|4|4|4|4|4|3.67|-18.26|4|3|3|3.33|3|4|4|3.67|-9.26|5|5|4|5|4.75|5|4|4|5|4.5|5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|2|2.5|2|2|2|25|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|45.5||2|2|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|Black||42|28273|Masters Degree|Divorced|Business: Marketing||1|6|Michael Baisden|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502181148|31|0|2|502184470|31|0|2|500454904|2||500004772||4|1|500000294, 500004640, 500004901|500000294|-2|500000294|-2|7016|11|||11146|1|||1|314390|134611|4|3|45
502590651|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2013-08-22|Followup|2012-06-30|2012-07-02|Complete|Done|3|2|2|2|4|4|2.83|4|3|4|2|4|4|3.5|-19.14|2|3|4|2|2|3|2.67|2|4|3|1|2|4|2.67|0|4|4|4|4|4|4|4|4|0|5|4|4|5|4.5|5|4|5|5|4.75|-5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|3|3.67|3|4|4|3.67|0|3|4|3.5|4|3|3.5|0|2|2|1|1|100|4|4|4|4|0|Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|25.8||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||36|28205|Bachelors Degree|Single|Business: Marketing|28117|7|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011746|502591168|31|0|2|502589724|1|0|2|500542166|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|314403|294373|4|3|45
501731841|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-05|2013-08-30|Followup|2012-06-05|2012-07-29|Comprehension|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|50.8||1|1|1|1|F|Black||18|Yes|Father|28210|One Parent: Male|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||49|28277|Bachelors Degree|Single|Business: Mgt, Admin||4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|501732181|31|0|2|501182066|31|0|2|500367022|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||46|2|||1|314408||4|2|45
502646551|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-07-03|Followup|2012-06-30|2012-07-03|Comprehension|Done||||||||4|3|4|3|3|3|3.33|||||||||2|3|3|3|3|3|2.83||||||4|3|3|3.33|||||||3|4|3|4|3.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||3|2|2.5||||1|1||||4|4||Green|Project Big|Child/Family: Moved|12.1||1|1|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|White||34|28210|High School Graduate|Single|Business: Sales|28269|0|8|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502598113|31|0|2|502262622|1|0|2|500543369|2||500004641||4|1|500004640|500004640|-2|500004640|-2|0|10|||7464|9|||1|314413|312938|4|2|45
501257717|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-20|2012-10-30|Followup|2012-06-20|2012-08-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|52.3||2|2|2|2|F|Black||17|No|GrandMother|28203|Grandparents|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|White||31|28204|Bachelors Degree|Single|Finance: Banking||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|501257994|31|0|2|500839705|1|0|2|500271936|2||-2||4|1|||-2||-2|0|10|||46|2|||1|314430||4|1|45
502549829|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-30|NaT|Followup|2012-06-30|2012-07-02|Complete|Done|2|2|2|1|2|2|1.83|3|1|2|1|2|2|1.83|0|1|2|2|1|1|2|1.5|2|3|2|2|2|2|2.17|-30.88|4|4|4|4|3|2|2|2.33|71.67|3|3|4|4|3.5|3|2|2|3|2.5|40|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|3|4|4|3.67|4|4|4|4|-8.25|4|4|4|3|3|3|33.33|2|2|1|1|100|4|4||||Green|Amachi, Project Big, Project Big AND Amachi||68.5||1|1|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|Amachi, PERL 2014-2016, Project Big, Project Big AND Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Business: Engineer|30357|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|1|502594393|31|0|1|500541795|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901, 500014681|-1||-2|0|4|||7464|9|||1|314431|283404|4|3|45
502645489|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-07-03|Followup|2012-06-30|2012-07-03|Comprehension|Done||||||||4|4|4|3|4|3|3.67|||||||||3|4|3|3|3|3|3.17||||||4|3|3|3.33|||||||4|4|3|4|3.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Green|Project Big|Child/Family: Moved|12.1||1|1|1|1|F|Black||20||Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||43|28214|Masters Degree|Married|Arts, Entertainment, Sports|28202|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502508948|31|0|2|502480739|31|0|2|500543463|2||500004641||4|1|500004640|500004640, 500005291|-2||-2|0|4|||7464|9|||1|314438|313195|4|2|45
502645484|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-11-13|Baseline|2011-06-30|2011-06-30|Complete|Done|2|2|2|2|1|2|1.83|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|3|4|4|4|3.86||||||||||4|4|3|3.67||||||3|4|3.5|||||2|2||||4|4||||Green|Project Big|Child/Family: Moved|16.5||1|1|1|1|F|Black||17||Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||26|28223||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502508948|31|0|2|502291769|31|0|2|500544311|2||-2||4|1|500004640|500004640, 500005291|-2||-2|0|10|||7464|9|||1|314442|-1|4|3|44
502645484|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-11-13|Followup|2012-06-30|2012-07-03|Declined|Done||||||||2|2|2|2|1|2|1.83|||||||||4|3|4|4|4|4|3.83||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|3|4|4|4|3.86||||||4|4|3|3.67|||||3|4|3.5||||2|2||||4|4||Green|Project Big|Child/Family: Moved|16.5||1|1|1|1|F|Black||17||Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||26|28223||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502508948|31|0|2|502291769|31|0|2|500544311|2||-2||4|1|500004640|500004640, 500005291|-2||-2|0|10|||7464|9|||1|314446|314442|4|1|45
502551116|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2013-08-01|Followup|2012-06-30|2012-07-02|Complete|Done|3|2|3|2|4|4|3|2|2|2|2|1|2|1.83|63.93|2|3|4|1|3|4|2.83|4|3|4|4|4|4|3.83|-26.11|4|4|4|4|4|4|4|4|0|3|2|2|4|2.75|4|3|5|5|4.25|-35.29|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|4|3.86|0|4|4|4|4|4|4|3|3.67|8.99|4|4|4|3|4|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Moved|25.1||1|1|2|2|F|Hispanic||17|Yes|GrandFather|28216|One Parent: Male|$15,000 to $19,999||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black|Other African|36|28105||Single|Consultant|28244|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|502551569|3|0|2|500892262|31|31|2|500541956|2||500004772||4|2|500000294, 500004640, 500004901, 500005291|500004640, 500005291|-2||-2|0|4|||46|2|||1|314461|291380|4|3|45
502489575|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2012-08-29|Followup|2012-06-30|2012-08-29|Declined|Late||||||||4|2|3|1|4|4|3|||||||||3|4|3|3|4|3|3.33||||||4|4|4|4|||||||3|5|4|5|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|3|2.5||||2|2||||4|4||Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|14||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||44|28105|Masters Degree|Married|Business: Mgt, Admin|28202|3|6|Ally Financial|Workplace Partner|Big|General Site||RTBM|277|60|598|500000170|500011746|502490022|31|0|1|502432606|31|0|1|500541789|2||-2||4|3|500004640, 500005291|500005291|-2||-1|56|1|||12831|3|1209, 635|1|1|314472|307800|4|1|45
502067798|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-09|NaT|Followup|2012-07-09|2012-07-11|Complete|Done|3|2|4|4|4|4|3.5|4|1|1|1|1|4|2|75|1|4|3|2|1|3|2.33|2|3|4|1|1|4|2.5|-6.8|4|4|4|4|4|4|4|4|0|2|3|4|2|2.75|1|4|5|2|3|-8.33|4|4|4|4|4|4|4|4|3|4|4|4|2|4|3|3.43|16.62|4|4|4|4|2|2|3|2.33|71.67|3|3|3|2|4|3|0|2|2|2|2|0|4|4||||Green|||80.2||1|1|1|1|M|Black||17|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||52|28270|Bachelors Degree|Married|Business: Mgt, Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|0|1|502062408|1|0|1|500459576|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|314792|154145|4|3|45
502478700|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-09|2014-11-13|Baseline|2011-07-05|2011-08-09|Complete|Done|4|4|4|2|2|4|3.33|||||||||2|4|4|3|4|4|3.5|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|39.2||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28027|Masters Degree|Single|Business: Engineer|28262|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|277|60|598|500000170|500013781|502881024|31|0|1|502578355|1|0|1|500544505|2||-2||4|3|500005291|500005291|-2|500015184|-1|0|5|||7462|13|||1|315352|-1|4|3|44
501226882|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-21|2013-06-07|Followup|2012-04-21|2012-07-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|61.5||1|1|2|2|M|Black||18|Yes|GrandMother|28027|Grandparents|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||52|28027|Bachelors Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500002335|501227158|31|0|1|500914929|31|0|1|500259581|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||2238|7|||1|315464||4|0|45
500186952|BBBS of Greater Charlotte|Main Office|C|Active|2004-07-15|NaT|Followup|2012-07-15|2012-07-09|Complete|Done|4|4|2|2|4|4|3.33|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|Amachi||152||1|1|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||73|28203||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|500188132|31|0|2|500189723|1|0|2|500037836|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|315573||4|3|45
500186946|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-20|2012-08-23|Followup|2012-06-20|2012-07-27|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Lost contact with child/agency|62.1||2|2|1|1|F|Black||19|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||36|28262||Single|Education: Teacher||4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188139|31|0|2|500865596|31|0|2|500181565|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|315593||4|1|45
500186956|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-21|2015-03-04|Followup|2012-06-21|2012-07-21|Complete|Done|4|4|4|4|4|3|3.83|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|128.4||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28203|Bachelors Degree|Married|Law: Lawyer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|500189727|1|0|1|500037841|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|315595||4|3|45
500186107|BBBS of Greater Charlotte|Main Office|C|Completed|2006-06-22|2012-10-17|Followup|2012-06-22|2012-06-12|Complete|Done|3|3|3|3|3|3|3|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|75.9||2|2|1|1|M|Black||22||Mother|28206|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|Black||52|28210|Masters Degree|Married|Business: Mgt, Admin||0|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500012459|500187654|31|0|1|500392161|31|0|1|500102003|2||-2||4|1|||-2||-2|0|10|||2230|7|||1|315783||4|3|45
502179818|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-16|2013-02-26|Followup|2012-07-16|2012-07-03|Complete|Done|3|4|3|2|3|4|3.17|||||||||2|3|3|3|2|3|2.67|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Moved|31.4||1|1|1|1|F|Black||14|Yes|GrandMother|28216|Grandparents|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Enrollment|F|Black||28|28216||Single|Student: College||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502180247|31|0|2|502057930|31|0|2|500460281|2||500003586||4|2|500000294|500000294|-2|500000294|-2|5635|9|||7464|9|||1|315785||4|3|45
500545328|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-02|2016-09-30|Followup|2012-07-02|2012-07-30|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|99||3|3|1|1|F|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|F|Black||43|28208|Masters Degree|Single|Business: Sales|28078|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|2|501033808|31|0|2|500274449|2||-2||4|1|||-2||-2|0|10|||46|2|||1|315922||4|3|45
500186277|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2014-07-16|Followup|2012-07-08|2012-07-09|Complete|Done|3|2|2|2|3|3|2.5|||||||||1|4|3|1|1|4|2.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Child/Family: Moved|60.3||3|4|2|3|F|Black||18||Mother|28206|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||39|28210|Bachelors Degree|Married|Business: Sales||8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500187876|31|0|2|500188587|1|0|2|500373187|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|316019||4|3|45
501129794|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-14|2015-10-29|Followup|2012-06-14|2012-07-02|Complete|Done|4|1|4|2|2|2|2.5|||||||||2|3|3|4|2|3|2.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|3|2.5|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|52.5||1|2|1|2|M|Black||14||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|F|Black||45|28273|Masters Degree|Single|Tech: Research/Design||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500017777|501130068|31|0|1|500922570|31|0|2|500540937|2||-2||4|1|||-2||-2|0|4|||46|2|||1|316565||4|3|45
500187077|BBBS of Greater Charlotte|Main Office|C|Completed|2005-05-31|2013-04-02|Followup|2012-05-31|2012-05-21|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|4|1|2|4|3.17|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green||Child: Graduated|94.1||2|2|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||41|28210|Bachelors Degree|Married|Medical: Pharmacist||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500188224|31|0|1|500189824|1|0|2|500037944|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|316876||4|3|45
500740295|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2012-06-12|2012-06-06|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Yellow||Volunteer: Feels incompatible with child/family|85||1|1|1|1|M|Black||18||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|White||55|28216|Bachelors Degree|Divorced|Tech: Engineer||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500794907|1|0|1|500179696|2||-2||4|2|||-2||-2|0|5|||46|2|||1|317024||4|3|45
501631059|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-26|2012-09-10|Followup|2012-05-26|2012-07-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|39.5||1|1|1|1|F|Black||18|No|Mother|28202|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||29|28216|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|501631382|31|0|2|501589359|31|0|2|500364875|2||-2||4|2|||-2|500000294|-2|34|2|||7464|9|||1|317061||4|1|45
501609876|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-13|2016-04-29|Followup|2012-07-13|2012-07-26|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Child: Graduated|81.5||1|2|1|2|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Black||38|28269|Masters Degree|Single|Medical: Nurse|28262|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501610196|31|0|2|501425392|31|0|2|500373716|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7464|9|||1|317181||4|3|45
501604440|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-23|2014-11-19|Followup|2012-07-23|2012-09-06|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|63.9||1|1|1|1|M|Black||20|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||38|28269||Married|Govt||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501758365|3|0|1|500373108|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|317189||4|1|45
502637589|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-19|2014-06-09|Baseline|2011-07-12|2011-07-19|Complete|Done|4|2|2|1|2|4|2.5|||||||||1|4|3|3|1|1|2.17|||||||||4|4|4|4||||||2|3|2|5|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Moved|34.7||1|1|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||30|28203|Masters Degree|Single|Business: Marketing|28203|0|10|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|502638284|31|0|2|502619035|1|0|2|500545174|2||-2||4|1|500005291|500005291|-2||-2|6854|8|||131|1|||1|317220|-1|4|3|44
502606280|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-21|2012-01-05|Baseline|2011-07-14|2011-07-21|Complete|Done|2|1|3|2|3|3|2.33|||||||||1|1|2|1|1|2|1.33|||||||||4|4|4|4||||||2|2|2|2|2|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Time constraints|5.5||1|1|1|1|F|White||15|No|Mother|28081|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI|RTBM|F|White||45|28078|Bachelors Degree|Married|Business: Human Resources||2|0|BBBS National Site|Web Link|Big|General Community||RTBM|277|60|598|500000170|500002335|502606797|1|0|2|501177078|1|0|2|500546219|2||-2||4|1|500005291|500005291|-2||-2|0|4|||46|2|||1|318471|-1|4|3|44
502555551|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-21|2012-07-26|Baseline|2011-07-14|2011-07-21|Complete|Done|4|1|2|1|4|3|2.5|||||||||2|3|3|2|4|3|2.83|||||||||3|3|4|3.33||||||5|3|3|4|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||4|4|4|||||2|2|||||||||Red|Project Big|Volunteer: Moved|12.2||2|2|1|1|M|Black||16|No|Aunt|28213|One Parent: Female|$40,000 to $44,999||Yes||School|General Community|Project Big|Match Support|M|White||27|28205|Associate Degree|Single|Service: Restaurant||0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502556004|31|0|1|502629285|1|0|1|500546255|2||-2||4|3|500004640|500004640|-2||-2|0|4|||7464|9|||1|318541|-1|4|3|44
502631914|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2014-08-28|Baseline|2011-07-14|2011-07-28|Complete|Done|4|4|4|1|4|4|3.5|||||||||1|1|3|3|1|4|2.17|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|3|2|||||1|1|||||||||Red||Volunteer: Moved|37||1|1|1|1|F|Black||18|No|Mother|28215|One Parent: Female|$20,000 to $24,999||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||37|28205|Associate Degree|Single|Medical: Healthcare Worker|28205|7|10|Local Print|Media|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013781|502632569|31|0|2|502581901|1|0|2|500546271|2||-2||4|3||500005291|-2|500004640|-2|6854|8|||7439|1|||1|318565|-1|4|3|44
500478936|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-14|2013-11-11|Followup|2012-07-14|2012-07-30|Complete|Done|4|1|1|1|4|4|2.5|||||||||2|4|3|3|3|4|3.17|||||||||3|3|3|3||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green||Child: Graduated|63.9||1|1|3|3|M|Black||21|No|Mother|28078|One Parent: Female|$25,000 to $29,999||No||Neighbor/Friend|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|500479187|31|0|1|501284751|31|0|1|500275964|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|8|||132|8|||1|318857||4|3|45
500910040|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2014-05-08|Followup|2012-05-29|2012-07-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|59.3||1|1|1|1|M|White||21|No|Mother|28270|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||31|28209|||Human Services: Non-Profit|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500910310|1|0|1|501600417|1|0|1|500363806|2||||4|3|||-2||-2|0|10|||7464|9|||1|318974||4|1|45
501721760|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-22|2016-11-01|Followup|2012-06-22|2012-08-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Infraction of match rules/agency policies|88.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||59|28269|Masters Degree|Married|Clergy||0|0|Coca Cola|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|501722098|31|0|1|501755476|1|0|1|500368545|2||-2||4|1|||-2|500000294|-2|0|10|||9610|3|||1|318985||4|1|45
500771746|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2016-06-15|Followup|2012-05-29|2012-07-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Child: Graduated|84.6||3|4|1|2|F|Black||19||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||37|28012|Some College|Married|Finance: Banking|28208|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500772014|31|0|2|500996153|1|0|2|500366437|2||500004641||4|1|500004640||-2||-2|0|4|||7464|9|||1|318993||4|1|45
502544579|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-21|2013-04-25|Followup|2012-04-21|2012-04-11|Complete|Done|4|2|2|1|1|4|2.33|||||||||3|4|4|1|3|4|3.17|||||||||4|2|3|3||||||5|2|5|5|4.25|||||||4|4|4|4|4|3|2|3.57||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|24.1||1|1|1|1|F|Hispanic||14|No|Mother|28213|Two Parent|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Hispanic||35|28078|Bachelors Degree|Married|Human Services: Social Worker|28208|3|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502540313|3|0|2|501718489|3|0|2|500532120|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|319087||4|3|45
501101149|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-01|NaT|Followup|2012-07-01|2012-08-15|Complete|Done|3|2|3|3|3|4|3|||||||||3|3|3|2|3|4|3|||||||||4|4|4|4||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|||104.5||1|2|1|2|F|White||16||Mother|28270|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||55|28277|Masters Degree|Widowed|Consultant||5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|501101423|1|0|2|500834694|1|0|2|500276073|2||-2||2|2|||-2||-2|0|4|||7671|13|||1|319139||4|3|45
501014187|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-07|NaT|Followup|2011-11-07|2011-11-21|Complete|Done|3|2|3|3|3|2|2.67|||||||||2|3|2|2|2|2|2.17|||||||||4|3|3|3.33||||||4|3|3|3|3.25|||||||4|4|4|4|4|3|3|3.71||||||||||3|3|3|3||||||3|2|2.5|||||1|1||||4|4||||Green|Amachi||100.2||2|2|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||48|28205|Bachelors Degree|Living w/ Significant Other|Human Services: Non-Profit|28205|3|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501404007|1|0|2|500306699|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7671|13|||1|319260||4|3|45
500835156|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2016-11-10|Followup|2012-07-10|2012-07-23|Complete|Done||||||||||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|100||1|2|1|2|M|Black||17||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Multi-Race (None of the above)||38|29710|Bachelors Degree|Single|Architect||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500835425|31|0|1|500466903|7|0|1|500277232|2||-2||4|1|||-2||-2|0|4|||46|2|||1|319325||4|3|45
501604443|BBBS of Greater Charlotte|Main Office|C|Active|2009-07-10|NaT|Followup|2012-07-10|2012-09-04|Blank|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||92.2||1|1|1|1|M|Black||18|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||35|28209|Bachelors Degree|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501729878|1|0|1|500371104|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|319390||4|3|45
500395038|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-01|2015-02-20|Followup|2012-08-01|2012-09-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|102.7||1|1|1|1|M|White||20||Mother|28226|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|M|White||39|28211|Masters Degree|Married|Law: Lawyer|28204|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500395288|1|0|1|500392006|1|0|1|500104016|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|319393||4|1|45
501228176|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-05|2013-08-13|Followup|2012-08-05|2012-07-18|Complete|Early|4|3|3|4|4|3|3.5|||||||||2|3|4|2|2|4|2.83|||||||||4|4|4|4||||||3|4|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|60.3||1|1|1|1|M|Black||20|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|28078|Masters Degree|Married|Finance: Auditor|28202|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|501228452|31|0|1|501279790|1|0|1|500279399|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|319471||4|3|45
501347097|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-30|2014-10-16|Followup|2012-07-30|2012-10-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|74.5||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||35|28078|Bachelors Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501347376|31|0|2|501099568|1|0|2|500278256|2||-2||4|2|||-2||-2|0|10|||46|2|||1|319475||4|0|45
502171910|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2015-08-25|Followup|2012-07-30|2012-10-14|Expired|Late||||||||3|1|2|2|2|3|2.17|||||||||2|3|3|4|2|4|3||||||4|4|4|4|||||||4|3|4|3|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Red|Amachi|Volunteer: Time constraint|60.8||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28214|Some College|Married|Medical||3|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502172339|31|0|1|502141964|31|0|1|500460627|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|5|||7464|9|||1|319485|156504|4|0|45
502303088|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2016-08-29|Followup|2012-06-27|2012-05-22|Complete|Early|4|3|4|1|4|4|3.33|||||||||2|4|4|1|2|4|2.83|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Project Big|Volunteer: Time constraint|62.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community|Project Big|Enrollment|F|Black||33|28215|Bachelors Degree|Single|Human Services: Social Worker|28217|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017777|502303520|31|0|2|502445797|31|0|2|500533193|2||-2||4|1|500004640|500004640|-2|500000294, 500004640|-2|6854|8|||7464|9|||1|319588||4|3|45
502294498|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-11|2013-08-15|Baseline|2011-07-19|2011-08-11|Complete|Done|3|1|3|3|3|3|2.67|||||||||2|3|3|1|2|3|2.33|||||||||3|2|2|2.33||||||4|3|3|3|3.25|||||||3|3|3|3|4|3|3|3.14||||||||||3|4|2|3||||||3|3|3|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|24.1||1|1|1|1|M|Some Other Race||16|No|Mother|28105|One Parent: Female|Unknown||No||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||47|28227|Some College|Single|Finance: Banking|28262|22|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502294930|41|0|1|502639594|31|0|1|500546657|2||-2||4|3|500005291|500005291|-2||-2|0|5|||7464|9|||1|319638|-1|4|3|44
502183217|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-05|NaT|Followup|2012-08-05|2012-07-25|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|4|2|3|3|||||||||4|4|4|4||||||4|2|3|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|4|3|||||2|2||||4|4||||Green|Amachi||79.3||1|1|2|2|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|Black||50|28078|||Service: Restaurant|28082|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502183646|31|0|1|501733851|31|0|1|500462588|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|319641||4|3|45
500280148|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-13|NaT|Followup|2012-07-13|2012-08-24|Complete|Done|4|4|4|4|4|4|4|||||||||4|1|4|4|4|4|3.5|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi||80.1||3|3|1|1|F|Black||16|Yes|Mother|28205|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|F|Black||30|28216|Bachelors Degree|Single|Human Services: Non-Profit|28216|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188151|31|0|2|502118494|31|0|2|500460767|2||500003586||2|2|500000294|500000294|-2||-2|0|3|||7464|9|||1|319644||4|3|45
500185647|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-09|2013-10-31|Followup|2012-07-09|2012-07-21|Complete|Done|3|2|4|3|4|3|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Child: Graduated|123.8||1|2|1|2|F|Black||21|Yes|Mother|28217|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||38|28269|Bachelors Degree|Married|Unknown|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187284|31|0|2|500188649|31|0|2|500038124|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|319645||4|3|45
500896588|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2016-06-15|Followup|2012-07-20|2012-07-23|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|3|3|3|3|3|3.17|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|3|4|3|3.71||||||||||2|2|2|2||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|106.9||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28273|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||36|28269|Masters Degree|Married|Education|28205|6|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|500896858|3|15|2|500924445|1|0|2|500183434|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|319655||4|3|45
501072636|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-25|2013-06-19|Followup|2012-06-25|2012-08-10|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|47.8||2|2|1|1|M|White||18||Mother|28134|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||50|28277|Bachelors Degree|Married|Tech: Management||10|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500004169|500965396|1|0|1|501637727|1|0|1|500368653|2||-2||4|3|||-2|500000294|-2|0|10|||7462|13|||1|319659||4|1|45
502637589|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-19|2014-06-09|Followup|2012-07-19|2012-07-23|Complete|Done|4|4|2|1|3|4|3|4|2|2|1|2|4|2.5|20|1|4|3|1|2|3|2.33|1|4|3|3|1|1|2.17|7.37|4|4|4|4|4|4|4|4|0|4|3|4|5|4|2|3|2|5|3|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Moved|34.7||1|1|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||30|28203|Masters Degree|Single|Business: Marketing|28203|0|10|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|502638284|31|0|2|502619035|1|0|2|500545174|2||-2||4|1|500005291|500005291|-2||-2|6854|8|||131|1|||1|319679|317220|4|3|45
502588461|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-22|2016-04-29|Baseline|2011-07-19|2011-07-22|Complete|Done|3|3|2|2|2|3|2.5|||||||||3|4|4|3|2|4|3.33|||||||||4|3|4|3.67||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Child: Graduated|57.3||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||46|28278|Bachelors Degree|Separated|Transport: Pilot|28208|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|502588977|31|0|1|502636478|31|0|1|500546741|2||-2||4|3|500005291|500005291|-2||-2|6854|8|||46|2|||1|319772|-1|4|3|44
502335675|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-30|2016-10-31|Followup|2011-12-30|2012-01-24|Complete|Done|4|2|4|2|3|3|3|||||||||2|4|4|3|4|3|3.33|||||||||4|4|4|4||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4|||||||4||||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi|Child: Lost interest|70||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|Project Big AND Amachi|Match Support|M|White||27|28262||Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502336110|31|0|1|502305990|1|0|1|500495220|2||500004772||4|3|500000294, 500004640, 500004901|500004901|-2|500000294, 500004640|-2|0|4|||7496|10|||1|319969||4|3|45
502252828|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2015-10-13|Baseline|2011-07-20|2011-08-03|Complete|Done|4|1|4|4|1|2|2.67|||||||||1|2|1|2|2|2|1.67|||||||||1|1|1|1||||||4|3|2|1|2.5|||||||4|4|4|4|4|4|4|4||||||||||2|2|3|2.33||||||4|3|3.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|50.3||1|1|1|1|M|Black||15||GrandMother|28227|Grandparents|Unknown||No||Self|General Community|PERL 2014-2016|RTBM|M|White||27|28205|Associate Degree|Single|Law: Police Officer||0|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502253254|31|0|1|502602451|1|0|1|500547383|2||-2||4|1|500005291|500014681|-2|500005291|-2|0|10|||7496|10|||1|320066|-1|4|3|44
501185592|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-23|2016-03-03|Followup|2012-06-23|2012-07-09|Complete|Done|3|4|3|2|3|3|3|||||||||2|4|4|3|2|3|3|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Family structure changed|92.3|Y|1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||45|28211||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501255830|1|0|1|500270254|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|320476||4|3|45
502555551|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-21|2012-07-26|Followup|2012-07-21|2012-07-24|Declined|Done||||||||4|1|2|1|4|3|2.5|||||||||2|3|3|2|4|3|2.83||||||3|3|4|3.33|||||||5|3|3|4|3.75||||||||||4|4|4|4|3|4|3|3.71||||||3|4|3|3.33|||||4|4|4||||2|2|||||||Red|Project Big|Volunteer: Moved|12.2||2|2|1|1|M|Black||16|No|Aunt|28213|One Parent: Female|$40,000 to $44,999||Yes||School|General Community|Project Big|Match Support|M|White||27|28205|Associate Degree|Single|Service: Restaurant||0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502556004|31|0|1|502629285|1|0|1|500546255|2||-2||4|3|500004640|500004640|-2||-2|0|4|||7464|9|||1|320510|318541|4|1|45
501716763|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-07|2016-11-11|Followup|2012-05-07|2012-07-22|Expired|Late||||||||1|1|1|1|1|1|1|||||||||2|1|2|2|3|2|2||||||3|3|3|3|||||||2|3|2|2|2.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||1|1|||||||Red||Child/Family: Lost contact with volunteer/agency|78.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Amachi, Cabarrus County|Match Support|F|Black||39|28269||Single|Self-Employed, Entrepreneur|28027|7|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501716992|31|0|2|502112513|31|0|2|500449029|2||-2||4|3||500000294, 500016374|-2|500016374|-2|6854|8|||7458|9|||1|320757|30228|4|0|45
502588461|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-22|2016-04-29|Followup|2012-07-22|2012-07-26|Complete|Done|1|2|4|1|3|3|2.33|3|3|2|2|2|3|2.5|-6.8|3|4|3|2|3|3|3|3|4|4|3|2|4|3.33|-9.91|4|3|3|3.33|4|3|4|3.67|-9.26|5|4|5|4|4.5|4|5|4|5|4.5|0|4|3|4|4|4|4|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|3|4|3|3.33|20.12|2|4|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Child: Graduated|57.3||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||46|28278|Bachelors Degree|Separated|Transport: Pilot|28208|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|502588977|31|0|1|502636478|31|0|1|500546741|2||-2||4|3|500005291|500005291|-2||-2|6854|8|||46|2|||1|320869|319772|4|3|45
502581001|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2014-01-30|Baseline|2011-07-25|2011-07-28|Complete|Done|4|1|4|1|1|1|2|||||||||4|1|4|4|2|4|3.17|||||||||4|4|3|3.67||||||5|4|4|5|4.5|||||||4|4|4|4|3|4|3|3.71||||||||||1|4|4|3||||||1|1|1|||||1|1|||||||||Red||Volunteer: Feels incompatible with child/family|30.1||1|1|1|1|M|Black||15|No|Mother|28210|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013781|502581504|31|0|1|502650916|31|0|1|500547358|2||-2||4|3||500005291|-2|500000294|-2|34|2|||7496|10|||1|321312|-1|4|3|44
501312033|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-04|2013-02-27|Followup|2012-06-04|2012-07-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Lost interest|32.8||2|2|1|1|F|Black||17|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||35|28226|||Customer Service||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500015820|501312311|31|0|2|502053746|31|0|2|500452835|2||-2||4|3||500000294|-2||-2|0|10|||7464|9|||1|321354||4|1|45
502179379|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-25|2015-07-31|Followup|2012-07-25|2012-09-05|Complete|Done|4|3|4|2|3|4|3.33|4|4|4|4|2|4|3.67|-9.26|3|4|4|3|3|4|3.5|1|4|4|1|2|4|2.67|31.09|4|4|4|4|4|4|4|4|0|5|4|5|5|4.75|3|3|5|5|4|18.75|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|4|3|3.5|1|2|1.5|133.33|2|2|2|2|0|4|4||||Red|Project Big|Volunteer: Lost contact with child/agency|60.2||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|Black||34|28269||Single|Student: College||0|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|502179808|31|0|2|502161458|31|0|2|500461681|2||-2||4|3|500004640|500004640|-2||-2|0|10|||9221|5|||1|322403|158340|4|3|45
502631914|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2014-08-28|Followup|2012-07-28|2012-08-17|Complete|Done|3|4|4|1|4|4|3.33|4|4|4|1|4|4|3.5|-4.86|2|3|3|2|1|3|2.33|1|1|3|3|1|4|2.17|7.37|4|4|4|4|4|4|4|4|0|4|4|5|3|4|4|5|5|4|4.5|-11.11|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|3|3.86|-3.89|4|4|4|4|4|4|4|4|0|3|3|3|1|3|2|50|2|2|1|1|100|4|4||||Red||Volunteer: Moved|37||1|1|1|1|F|Black||18|No|Mother|28215|One Parent: Female|$20,000 to $24,999||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||37|28205|Associate Degree|Single|Medical: Healthcare Worker|28205|7|10|Local Print|Media|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013781|502632569|31|0|2|502581901|1|0|2|500546271|2||-2||4|3||500005291|-2|500004640|-2|6854|8|||7439|1|||1|322514|318565|4|3|45
502581001|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2014-01-30|Followup|2012-07-28|2012-07-25|Complete|Done|3|2|4|2|3|3|2.83|4|1|4|1|1|1|2|41.5|2|4|4|2|2|4|3|4|1|4|4|2|4|3.17|-5.36|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|4|5|4|4|5|4.5|-11.11|4|4|4|4|3|4|3|3.71|4|4|4|4|3|4|3|3.71|0|4|4|4|4|1|4|4|3|33.33|1|3|2|1|1|1|100|2|2|1|1|100|4|4||||Red||Volunteer: Feels incompatible with child/family|30.1||1|1|1|1|M|Black||15|No|Mother|28210|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013781|502581504|31|0|1|502650916|31|0|1|500547358|2||-2||4|3||500005291|-2|500000294|-2|34|2|||7496|10|||1|322530|321312|4|3|45
502593613|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2017-02-28|Baseline|2011-07-28|2011-08-19|Complete|Done|3|2||1|2|2||||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|3|3|3.33||||||3|3|3|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|66.4||1|1|1|1|F|Black||16|No|Mother|28208|Two Parent|$35,000 to $39,999|Y|Yes||Relative|General Community||Match Support|F|Hispanic||26|28217|Bachelors Degree|Single|Service: Restaurant||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502594130|31|0|2|502601730|3|0|2|500547881|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|322561|-1|4|3|44
502173588|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2012-08-30|Followup|2012-08-27|2012-08-13|Complete|Done|4|4|4|4|4|4|4|3|1|2|1|3|3|2.17|84.33|2|3|4|4|2|4|3.17|2|3|3|2|2|3|2.5|26.8|4|4|4|4|4|4|4|4|0|4|5|3|4|4|4|3|4|3|3.5|14.29|4|4|4|4|4|4|4|4|2|2|2|1|1|2|1|1.57|154.78|4|4|4|4|4|4|4|4|0|2|2|2|2|1|1.5|33.33|1|1|1|1|0|4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|24.1||2|2|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||No|A Child's Place|Service Organization|General Community|Amachi|Enrollment|F|White||29|28217|Bachelors Degree|Single|Customer Service||5|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502174017|31|0|2|502085998|1|0|2|500463449|2||500003586||4|2|500000294|500000294|-2||-2|7016|11|||7496|10|||1|322589|160541|4|3|45
501247286|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-14|2016-11-08|Followup|2012-05-14|2012-05-02|Complete|Done|4|3|4|4|2|4|3.5|||||||||2|3|4|4|4|4|3.5|||||||||4|2|2|2.67||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|101.8||1|1|1|1|M|White||15|No|Father|28025|One Parent: Male|Unknown||No||Self|General Community|Cabarrus County|Enrollment|M|White||49|27103|Masters Degree|Single|Education: Teacher|27282|0|0|Other|Service Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500341682|1|0|1|501247141|1|0|1|500264655|2||-2||4|1||500016374|-2|500016374|-2|0|10|||7452|6|||1|322895||4|3|45
502083456|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2013-07-22|Baseline|2011-07-29|2011-08-03|Complete|Done|2|2|1|1|3|2|1.83|||||||||1|2|3|2|2|3|2.17|||||||||4|3|3|3.33||||||3|2|3|1|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2|||||||||Green||Child/Family: Moved|23.6||1|1|1|1|F|Black||16|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||29|28262|Masters Degree|Single|Finance: Banking|28208|4|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Enrollment|277|60|598|500000170|500012459|502083880|31|0|2|502542333|31|0|2|500548042|2||-2||4|1|||-2|500014506|-1|0|10|||7671|13|||1|322957|-1|4|3|44
502492731|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-05|2012-03-29|Baseline|2011-07-29|2011-10-05|Complete|Done|3|4|3|3|4|3|3.33|||||||||2|4|3||3|4||||||||||4|4|4|4||||||2|5|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||2|3|2.5|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|5.8||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||51|28213|Bachelors Degree|Married|Medical|28208|11|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500001281|502493180|31|0|1|502677685|31|0|1|500557795|2||-2||4|2|||-2||-2|6854|8|||7438|1|||1|322981|-1|4|3|44
502453042|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2013-07-29|Baseline|2011-07-29|2011-08-03|Complete|Done|2|2|4|3|3|3|2.83|||||||||2|3|2|2|1|3|2.17|||||||||4|4|4|4||||||3|2|3|2|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|1|1.5|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|23.9||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||27|28213|Bachelors Degree|Single|Business: Marketing||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502453489|31|0|2|502632959|31|0|2|500548075|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|322995|-1|4|3|44
500186352|BBBS of Greater Charlotte|Main Office|C|Completed|2002-07-29|2014-01-02|Followup|2012-07-29|2012-08-03|Complete|Done|4|1|4|4|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|137.2||4|4|2|2|M|Black||21||Mother|28212|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|White||45|28226|Masters Degree|Married|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500187945|31|0|1|500189280|1|0|1|500037290|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|323086||4|3|45
501726201|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2015-01-30|Followup|2012-07-08|2012-08-27|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Moved|66.8||1|1|1|1|F|Black||17|Yes|Mother|28212|One Parent: Female|Unknown||Yes|YeaGod|Faith Organization|General Community|Amachi|Match Support|F|Black||51|28262|PHD|Married|Real Estate: Realtor||0|0|Weeping Willow|Faith Organization|Big|General Community||Enrollment|277|60|598|500000170|500008321|501726541|31|0|2|501734664|31|0|2|500371036|2||-2||4|3|500000294|500000294|-2||-2|5634|9|||9218|7|||1|323407||4|1|45
501213488|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-19|NaT|Followup|2012-05-19|2012-06-19|Complete|Done|3|2|3|2|3|3|2.67|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||105.9||1|1|1|1|F|White||14|No|Father|28207|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Finance: Banking|28255|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|501213764|1|0|2|501225276|1|0|2|500262655|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|326388||4|3|45
501524313|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-02|2014-04-21|Followup|2012-08-02|2012-09-06|Declined|Done||||||||2|2|3|2|3|3|2.5|||||||||3|3|3|3|3|3|3||||||3|3|3|3|||||||3|3|2|3|2.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Green|2010-2012 OJJDP JJI|Volunteer: Moved|32.6||2|2|1|1|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28208|Bachelors Degree|Single|Finance: Economist|28202|5|6|Recruitment Event|BBBS Board/Staff|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|501524605|31|0|1|502615076|1|0|1|500547406|2||-2||4|1|500005291|500005291|-2|500005291|-2|0|10|||7462|13|||1|326507|4772|4|1|45
501994951|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2014-09-18|Followup|2012-06-15|2012-07-30|Declined|Done||||||||3|3|3|1|4|4|3|||||||||4|4|3|4|4|4|3.83||||||4|4|4|4|||||||4|5|5|4|4.5||||||||||4|4|4|3|3|3|3|3.43||||||3|3|3|3|||||3|1|2||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|51.1||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|Unknown||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||36|28078||Single|Customer Service||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501843047|31|0|2|502048623|31|0|2|500455478|2||-2||4|2|||-2||-2|7294|13|||7464|9|||1|326534|139614|4|1|45
500934908|BBBS of Greater Charlotte|Main Office|C|Active|2010-06-18|NaT|Followup|2012-06-18|2012-07-24|Complete|Done|3|4|4|2|4|4|3.5|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|Amachi||80.9||2|2|1|1|M|Black||16|Yes|Aunt|28216|One Parent: Female|Less than $10,000|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||34|20175|Bachelors Degree|Single|Business: Sales|28211|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|500935173|31|0|1|502107314|1|0|1|500456443|2||500003586||2|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|326537||4|3|45
502252828|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2015-10-13|Followup|2012-08-03|2012-07-30|Complete|Done|4|2|1|2|2|4|2.5|4|1|4|4|1|2|2.67|-6.37|2|3|4|1|2|3|2.5|1|2|1|2|2|2|1.67|49.7|3|4|3|3.33|1|1|1|1|233|4|4|3|4|3.75|4|3|2|1|2.5|50|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|4|4|-7.25|4|3|3|3.33|2|2|3|2.33|42.92||||4|3|3.5||2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|50.3||1|1|1|1|M|Black||15||GrandMother|28227|Grandparents|Unknown||No||Self|General Community|PERL 2014-2016|RTBM|M|White||27|28205|Associate Degree|Single|Law: Police Officer||0|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502253254|31|0|1|502602451|1|0|1|500547383|2||-2||4|1|500005291|500014681|-2|500005291|-2|0|10|||7496|10|||1|326794|320066|4|3|45
502588295|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-27|2012-05-31|Baseline|2011-08-03|2011-09-27|Complete|Done|3|4|3|4|1|4|3.17|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|3|2|2|2.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||1|1|1|||||1|1||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Infraction of match rules/agency policies|8.1||1|1|1|1|F|Black||18|No|Mother|28208|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||38|28278|Bachelors Degree|Divorced|Business: Mgt, Admin|28269|1|0|Self|Self|Big|General Community||RTBM|277|60|598|500000170|500011746|502588811|31|0|2|502601476|1|0|2|500553687|2||-2||4|3|500004640, 500005291|500005291|-2||-2|0|10|||7464|9|||1|326814|-1|4|3|44
502083456|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2013-07-22|Followup|2012-08-03|2012-07-24|Complete|Done|2|1|1|1|2|2|1.5|2|2|1|1|3|2|1.83|-18.03|1|2|3|4|1|4|2.5|1|2|3|2|2|3|2.17|15.21|4|4|4|4|4|3|3|3.33|20.12|1|3|5|4|3.25|3|2|3|1|2.25|44.44|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3.5|14.29|2|2|2|2|0|4|4||||Green||Child/Family: Moved|23.6||1|1|1|1|F|Black||16|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||29|28262|Masters Degree|Single|Finance: Banking|28208|4|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Enrollment|277|60|598|500000170|500012459|502083880|31|0|2|502542333|31|0|2|500548042|2||-2||4|1|||-2|500014506|-1|0|10|||7671|13|||1|326972|322957|4|3|45
502453042|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2013-07-29|Followup|2012-08-03|2012-09-06|Declined|Done||||||||2|2|4|3|3|3|2.83|||||||||2|3|2|2|1|3|2.17||||||4|4|4|4|||||||3|2|3|2|2.5||||||||||4|4|4|4|4|4|3|3.86||||||3|3|3|3|||||2|1|1.5||||2|2||||4|4||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|23.9||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||27|28213|Bachelors Degree|Single|Business: Marketing||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502453489|31|0|2|502632959|31|0|2|500548075|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|326976|322995|4|1|45
502057402|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-28|2012-10-31|Followup|2012-07-28|2012-08-20|Complete|Done|3|3|4|3|3|3|3.17|4|3|4|4|3|4|3.67|-13.62|3|4|4|3|3|3|3.33|3|4|3|2|4|1|2.83|17.67|4|4|4|4|4|4|4|4|0|4|3|3|4|3.5|5|4|4|4|4.25|-17.65|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|4|3.33|4|3|4|3.67|-9.26|3|3|3|4|4|4|-25|2|2|2|2|0|4|4||||Red||Volunteer: Time constraint|27.1||1|1|1|1|M|White||17|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|White||38|28078|Some College|Married|Military||14|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502057826|1|0|1|502196301|1|0|1|500461316|2||-2||4|3|||-2|500000294|-2|0|4|||7496|10|||1|326985|157640|4|3|45
502222992|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-16|2013-12-12|Followup|2012-07-16|2012-09-04|Blank|Late||||||||3|3|3|1|2|3|2.5|||||||||2|4|3|2|2|4|2.83||||||4|4|3|3.67|||||||3|4|4|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Child: Graduated|40.9||1|1|1|1|F|Black||21|No|Aunt|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||32|28213|Bachelors Degree|Single|Education|28223|7|0|BBBS National Site|Web Link|Big|General Site||Enrollment|277|60|598|500000170|500017732|502223423|31|0|2|502085103|31|0|2|500461244|2||-2||4|1|||-2||-1|6854|8|||46|2|||1|326988|157522|4|3|45
500186174|BBBS of Greater Charlotte|Main Office|C|Completed|2005-07-28|2012-10-31|Followup|2012-07-28|2012-10-09|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|87.1||2|2|2|2|F|Black||18||Mother|28208|One Parent: Female|Unknown||No||Self|General Community||Enrollment|F|Black||48|29715|Some College|Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500187758|31|0|2|500189225|31|0|2|500038037|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|326989||4|1|45
502233621|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-14|2013-04-25|Followup|2012-08-14|2012-07-26|Complete|Early|4|3|4|3|4|4|3.67|3|4|4|4|3|4|3.67|0|4|3|4|4|4|4|3.83|4|1|4|2|4|4|3.17|20.82|4|4|4|4|4|4|4|4|0|5|4|4|3|4|5|5|4|5|4.75|-15.79|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|4|4|4|4|4|4|0|2|2|2|2|0|4|4||||Green||Child/Family: Moved|32.4||1|1|2|2|M|Multi-race (Hispanic & White)||16|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction|28208|1|1|Igniting Breakfast|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500011746|502234052|35|0|1|502255664|1|0|1|500465113|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17266|8|||1|326990|168275|4|3|45
501641337|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-07|2015-03-13|Followup|2012-08-07|2012-08-24|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|4|4|4|4|3|3.83|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|67.2||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||31|28269|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|2|500835981|31|0|2|500373972|2||-2||4|1||500000294|-2|500000294|-2|0|10|||46|2|||1|327089||4|3|45
502221904|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-06|2013-01-31|Followup|2012-08-06|2012-10-21|Expired|Late||||||||3|1|2|1|4|3|2.33|||||||||1|1|2|1|2|2|1.5||||||4|4|4|4|||||||2|2|3|3|2.5||||||||||4|4|4|4|4|4|4|4||||||2|4|1|2.33|||||3|3|3||||2|2|||||||Red|Amachi|Child/Family: Infraction of match rules/agency policies|29.9||1|1|3|3|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Arby's|Workplace Partner/Business|General Community||Match Support|F|Black||36|28078|Masters Degree|Married|Business: Marketing|28273|1|1|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|277|60|598|500000170|500015820|502222335|31|0|2|502056302|31|0|2|500464397|2||500003586||4|3|500000294||-2|500014505, 500014506|-1|3394|14|||7671|13|||1|327107|167141|4|0|45
502254067|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-10|2013-01-03|Followup|2011-09-10|2011-09-06|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|1|1|1|1|1|1.5|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|2|3.71||||||||||1|4|1|2||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|27.8||3|3|1|1|F|Black||14|No|Mother|28209|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|Black||37|28210|Bachelors Degree|Single|Insurance||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502254499|31|0|2|502214352|31|0|2|500466835|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|327327||4|3|45
502666718|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2013-07-25|Baseline|2011-08-05|2011-08-19|Complete|Done|4|2|2|1|1|4|2.33|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Child/Family: Unrealistic expectations|23.2||1|1|2|2|F|Black||16|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||38|28202|Masters Degree||Business: Clerical||7|0|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502667545|31|0|2|500932879|31|0|2|500548835|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7458|9|||1|327460|-1|4|3|44
501809541|BBBS of Greater Charlotte|Main Office|C|Active|2009-08-07|NaT|Followup|2012-08-07|2012-08-09|Complete|Done|4|4|2|3|4|4|3.5|||||||||3|3|3|4|3|4|3.33|||||||||4|3|3|3.33||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||91.3||1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||49|28031|Bachelors Degree|Married|Transport: Pilot|40223|9|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501809896|36|0|1|501620528|1|0|1|500375025|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|327736||4|3|45
502652785|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2012-04-27|Baseline|2011-08-08|2011-08-19|Complete|Done|3|3|3|3|4|4|3.33|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow|2010-2012 OJJDP JJI|Volunteer: Time constraint|8.3||1|1|1|1|M|Multi-race (Black & Hispanic)||16|No|Mother|28270|One Parent: Female|$40,000 to $44,999||No|Arby's|Workplace Partner/Business|General Community|2010-2012 OJJDP JJI|RTBM|M|Some Other Race||43|28210|Associate Degree|Married|Finance: Banking|28204|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site||RTBM|277|60|598|500000170|500001281|502653521|38|0|1|502619698|41|0|1|500548958|2||-2||4|2|500005291|500005291|-2||-1|3394|14|||7462|13|||1|327823|-1|4|3|44
501010684|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-17|2013-03-14|Baseline|2011-08-08|2011-08-12|Complete|Done|4|2|1|3|3|1|2.33|||||||||1|2|3|1|3|1|1.83|||||||||4|4|4|4||||||4|5|3|3|3.75|||||||1|4|4|3|4|4|3|3.29||||||||||3|4|2|3||||||1|2|1.5|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Child/Family: Feels incompatible with volunteer|18.9||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Less than $10,000||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|White||46|28227|Bachelors Degree|Married|Business: Mgt, Admin|28277|10|0|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500004169|503560069|31|0|1|502570658|1|0|1|500549074|2||-2||4|3|500005291|500005291|-2||-2|7016|11|||7439|1|||1|327911|-1|4|3|44
502436202|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2015-07-13|Baseline|2011-08-08|2011-09-02|Complete|Done|3|2|2|1|3|3|2.33|||||||||3|3|3|4|2|4|3.17|||||||||4|4|4|4||||||2|5|5|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|4|3|||||1|1||||4|4||||Green||Child: Graduated|46.3||1|1|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|Masters Degree|Single|Finance: Banking||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502436645|31|0|1|502642999|1|0|1|500549046|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|327937|-1|4|3|44
502478700|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-09|2014-11-13|Followup|2012-08-09|2012-08-13|Complete|Done|4|4|4|4|4|4|4|4|4|4|2|2|4|3.33|20.12|1|4|4|4|1|4|3|2|4|4|3|4|4|3.5|-14.29|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|4|5|5|4.75|5.26|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|3|3.67|8.99|3|3|3|2|2|2|50|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|39.2||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28027|Masters Degree|Single|Business: Engineer|28262|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|277|60|598|500000170|500013781|502881024|31|0|1|502578355|1|0|1|500544505|2||-2||4|3|500005291|500005291|-2|500015184|-1|0|5|||7462|13|||1|328093|315352|4|3|45
502139829|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-12|2013-08-08|Followup|2012-08-12|2012-10-25|Declined|Late||||||||3|4|4|4|4|4|3.83|||||||||2|4|4|3|2|4|3.17||||||4|3|4|3.67|||||||5|4|4|4|4.25||||||||||4|4|4|4|3|3|3|3.57||||||4|4|3|3.67|||||4|2|3||||2|2|||||||Red||Volunteer: Lost contact with child/agency|35.9||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||30|28226|Masters Degree|Single|Finance: Accountant||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502140258|31|0|1|502178005|1|0|1|500462499|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|328128|159370|4|1|45
501240369|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-10-09|Followup|2012-07-10|2012-07-31|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|75||1|1|1|1|M|Black||20|Yes|Mother|28214|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||43|28269|Masters Degree|Single|Business: Mgt, Admin|28202|3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501240645|31|0|1|501240602|1|0|1|500272039|2||500003586||4|1|500000294|500000294|-2||-2|0|3|||131|1|||1|328149||4|3|45
500186682|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2015-07-22|Followup|2012-07-20|2012-07-16|Complete|Done|4|4|4|4|4|4|4|||||||||4|1|4|2|4|4|3.17|||||||||4|4|4|4||||||3|4|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|96.1||3|4|1|1|M|Black||20|Yes|Mother|28227|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|M|Black||57|28262||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|500887363|31|0|1|500184396|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|328150||4|3|45
500186960|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-31|2013-08-15|Followup|2012-07-31|2012-09-12|Complete|Done|4|4|4|4|4|4|4|||||||||1|4|4|1|2|4|2.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|72.5||2|2|1|1|M|White||19|Yes|Mother|28227|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||40|28105|Some College|Married|Military|28112|11|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188147|1|0|1|500738970|1|0|1|500186719|2||500003586||4|3|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|328151||4|3|45
500417281|BBBS of Greater Charlotte|Main Office|C|Completed|2006-07-31|2013-01-31|Followup|2012-07-31|2012-08-17|Complete|Done|3|4|4|1|3|3|3|||||||||4|4|3|4|4|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|78.1|Y|1|1|1|1|F|White||16||Mother|28211|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||48|28211|Masters Degree|Married|Finance: Banking|28202|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500402926|1|0|2|500349297|1|0|1|500112798|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|328153||4|3|45
501725168|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-31|2013-12-18|Followup|2012-08-31|2012-10-13|Complete|Done|4|4|4|2|3|4|3.5|||||||||2|2|3|3|1|4|2.5|||||||||4|4|4|4||||||5|3|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Moved|51.6||2|2|1|1|F|Multi-Race (None of the above)||15|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28269|Bachelors Degree|Married|Human Services: Non-Profit||2|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017777|501724831|7|0|2|501824761|1|0|2|500381463|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|328456||4|3|45
502205848|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-18|NaT|Baseline|2011-08-10|2011-08-18|Complete|Done|3|4|3|2|4|4|3.33|||||||||3|2|3|4|3|3|3|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||2|4|3|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI||66.9||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Juris Doctorate (JD)|Single|Student: College|28208|0|0||Law Student Association|Big|General Community||Match Support|277|60|598|500000170|500020753|502206277|31|0|1|502624702|1|0|1|500549350|2||-2||2|1|500005291|500005291|-2||-2|0|10|||0|15|||1|328511|-1|4|3|44
500383915|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-20|2012-08-30|Followup|2012-06-20|2012-07-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|50.3||2|2|2|2|F|Black||20||GrandMother|28205|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||64|28269||Married|Finance: Economist||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|500384165|31|0|2|500540512|31|0|2|500274279|2||-2||4|1|||-2||-2|6855|8|||7464|9|||1|328783||4|1|45
502064627|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-20|NaT|Followup|2012-08-20|2012-10-25|Declined|Late||||||||2|2|4|2|3|4|2.83|||||||||3|3|4|3|2|4|3.17||||||4|3|2|3|||||||5|3|3|4|3.75||||||||||4|4|4|4|4|4|4|4||||||3|2|3|2.67|||||2|3|2.5||||1|1|||||||Green|||78.9||1|1|2|2|M|Black||16|No|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|502065051|31|0|1|500773055|3|14|1|500462574|2||-2||2|1|||-2||-2|0|10|||46|2|||1|328844|159373|4|1|45
501641325|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-24|2015-08-03|Followup|2012-06-24|2012-08-08|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|73.3||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Multi-race (Asian & White)||34|28205|Bachelors Degree|Single|Tech: Research/Design|28255|3|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|1|501715652|37|0|1|500366872|2||-2||4|1||500000294|-2|500000294|-2|6854|8|||7464|9|||1|328852||4|1|45
500910037|BBBS of Greater Charlotte|Main Office|C|Active|2009-06-22|NaT|Followup|2012-06-22|2012-08-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||92.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||46|28277||Married|Business: Mgt, Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|500910307|31|0|1|500856100|1|0|1|500368834|2||-2||2|1|||-2||-2|0|10|||46|2|||1|328853||4|1|45
500826596|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2013-12-16|Followup|2012-07-28|2012-10-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|28.6||3|3|1|1|M|Black||17|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Black||29|28226|Some College|Single|Customer Service|28210|2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500826861|31|0|1|502549323|31|0|1|500544976|2||-2||4|2|500005291||-2|500000294|-2|0|5|||7464|9|||1|328858||4|0|45
502294498|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-11|2013-08-15|Followup|2012-08-11|2012-10-25|Declined|Late||||||||3|1|3|3|3|3|2.67|||||||||2|3|3|1|2|3|2.33||||||3|2|2|2.33|||||||4|3|3|3|3.25||||||||||3|3|3|3|4|3|3|3.14||||||3|4|2|3|||||3|3|3||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|24.1||1|1|1|1|M|Some Other Race||16|No|Mother|28105|One Parent: Female|Unknown||No||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||47|28227|Some College|Single|Finance: Banking|28262|22|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502294930|41|0|1|502639594|31|0|1|500546657|2||-2||4|3|500005291|500005291|-2||-2|0|5|||7464|9|||1|328925|319638|4|1|45
502034144|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-20|2014-12-04|Followup|2012-07-20|2012-09-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|52.5||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||RTBM|M|Some Other Race||45|28210|Bachelors Degree|Married|Education: Teacher||0|0|CIS/Hidden Valley|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500018987|502034543|31|0|1|502212267|41|0|1|500460434|2||||4|1|||-2||-2|34|2|||11522|6|||1|329230||4|1|45
501300101|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-14|2015-05-11|Followup|2012-08-14|2012-08-07|Complete|Done|3|4|4|4|1|3|3.17|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|80.9||1|1|4|4|F|Black||19|Yes|GrandMother|28273|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501300379|31|0|2|500346193|31|0|2|500281421|2||500003586||4|2|500000294|500000294|-2||-2|7294|13|||46|2|||1|329881||4|3|45
502467122|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-28|2011-10-06|Baseline|2011-08-15|2011-08-28|Complete|Done|4|2|4|2|4|4|3.33|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|Amachi|Child/Family: Feels incompatible with volunteer|1.3||1|1|2|2|M|Black||14|Yes|Mother|28214|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community|Amachi|Match Support|M|White||33|28214|Associate Degree|Single|Law: Security Officer|28208|2|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012319|502467569|31|0|1|502658498|1|0|1|500550136|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|329902|-1|4|3|44
501195410|BBBS of Greater Charlotte|Main Office|C|Active|2008-08-15|NaT|Followup|2012-08-15|2012-08-07|Complete|Done|4|1|4|1|4|4|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||103||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Asian||35|28210|Bachelors Degree|Married|Business: Sales|28217|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501195684|31|0|1|501277677|4|0|1|500278978|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|330024||4|3|45
502247430|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-17|2014-01-23|Followup|2012-08-17|2012-09-12|Complete|Done|2|4|2|3|2|4|2.83|3|1|1|1|2|3|1.83|54.64|3|4|3|1|3|3|2.83|2|2|3|1|2|2|2|41.5|4|4|4|4|4|3|3|3.33|20.12|3|4|3|4|3.5|2|3|2|4|2.75|27.27|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|4|3.67|2|4|4|3.33|10.21|3|2|2.5|2|1|1.5|66.67|1|1|1|1|0|4|4||||Yellow||Child: Lost interest|41.2||1|1|1|1|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||63|28078|Bachelors Degree|Married|Medical: Nurse||10|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502247861|31|0|2|502226106|1|0|2|500465539|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|330043|166252|4|3|45
500826594|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-21|2016-06-15|Followup|2012-08-21|2012-10-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|105.8||1|1|1|1|M|Black||18|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Some Other Race||36|28209|||Business: Sales||0|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|1|500920342|41|0|1|500185735|2||-2||4|1|||-2||-2|0|5|||6450|12|||1|330045||4|1|45
502097843|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-29|2016-08-11|Baseline|2011-08-16|2011-08-29|Complete|Done|3|2|2|1|4|3|2.5|||||||||2|3|3|2|3|3|2.67|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|||||||2|2||||4|4||||Green|2010-2012 OJJDP JJI|Child: Lost interest|59.4||1|1|2|2|M|Black||17|No|Mother|28078|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500021785|502098263|31|0|1|502643791|3|0|1|500550390|2||-2||4|1|500005291||-2||-2|0|10|||7496|10|||1|330290|-1|4|3|44
502569411|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-14|2012-12-19|Baseline|2011-08-16|2011-09-14|Complete|Done|4|4|4|2|3|4|3.5|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|Amachi, 2010-2012 OJJDP JJI|Child/Family: Time constraints|15.2||1|1|1|1|F|American Indian or Alaska Native||14|Yes|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||45|28027|||Medical: Nurse|28144|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502569865|6|0|2|502642653|1|0|2|500550403|2||500003586||4|2|500000294, 500005291|500005291|-2||-2|0|10|||7496|10|||1|330300|-1|4|3|44
501010684|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-17|2013-03-14|Followup|2012-08-17|2012-08-22|Declined|Done||||||||4|2|1|3|3|1|2.33|||||||||1|2|3|1|3|1|1.83||||||4|4|4|4|||||||4|5|3|3|3.75||||||||||1|4|4|3|4|4|3|3.29||||||3|4|2|3|||||1|2|1.5||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Child/Family: Feels incompatible with volunteer|18.9||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Less than $10,000||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|White||46|28227|Bachelors Degree|Married|Business: Mgt, Admin|28277|10|0|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500004169|503560069|31|0|1|502570658|1|0|1|500549074|2||-2||4|3|500005291|500005291|-2||-2|7016|11|||7439|1|||1|330538|327911|4|1|45
502636177|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-29|2013-09-19|Baseline|2011-08-17|2011-08-29|Complete|Done|4|1|4|1|4|3|2.83|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green||Volunteer: Moved|24.7||1|1|1|1|F|Black||14|No|GrandMother|28216|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|Black||30|28212||Single|Medical||0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502636872|31|0|2|502643313|31|0|2|500551053|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|330694|-1|4|3|44
502697677|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2013-03-27|Baseline|2011-08-18|2011-09-02|Complete|Done|4|3|3|3|3|3|3.17|||||||||2|4|3|3|2|4|3|||||||||4|4|4|4||||||5|5|4|2|4|||||||4|4|4|3|4|4|2|3.57||||||||||3|3|4|3.33||||||3|3|3|||||1|1||||4|4||||Yellow||Volunteer: Moved|18.8||1|1|1|1|F|Hispanic||19|No|Mother|28027|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|F|White||32|28027|Bachelors Degree|Single|Business: Marketing|28075|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502605848|3|0|2|502590370|1|0|2|500550704|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|330902|-1|4|3|44
502627461|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-26|2012-09-27|Baseline|2011-08-18|2011-08-26|Complete|Done|3|4|2|3|4|4|3.33|||||||||4|3|4|3|2|4|3.33|||||||||4|4|4|4||||||4|3|3|2|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|2|2|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Time constraint|13.1||1|1|1|1|F|Hispanic|Mexican|20|Yes|Mother|28269|One Parent: Female|Unknown|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||52|28205|Some College|Single|Self-Employed, Entrepreneur||16|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500011746|502628116|3|10|2|502615885|1|0|2|500550750|2||-2||4|3|500005291|500005291|-2|500005291|-2|0|4|||7464|9|||1|330948|-1|4|3|44
502601023|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-31|2016-08-11|Baseline|2011-08-18|2011-08-31|Complete|Done|3|2|3|1|3|4|2.67|||||||||3|3|4|2|2|3|2.83|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|2|4|4|3|4|3|3.43||||||||||3|4|2|3||||||3|3|3|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI|Child: Graduated|59.4||1|1|1|1|F|Black||19||Mother|28216|Two Parent|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||51|28277|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502601540|31|0|2|502546883|1|0|2|500550809|2||-2||4|1|500005291|500005291|-2||-2|6854|8|||7464|9|||1|331012|-1|4|3|44
502205848|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-18|NaT|Followup|2012-08-18|2012-11-02|Expired|Late||||||||3|4|3|2|4|4|3.33|||||||||3|2|3|4|3|3|3||||||4|4|4|4|||||||4|4|5|4|4.25||||||||||4|4|4|4|3|4|4|3.86||||||4|4|3|3.67|||||2|4|3||||1|1||||4|4||Green|2010-2012 OJJDP JJI||66.9||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Juris Doctorate (JD)|Single|Student: College|28208|0|0||Law Student Association|Big|General Community||Match Support|277|60|598|500000170|500020753|502206277|31|0|1|502624702|1|0|1|500549350|2||-2||2|1|500005291|500005291|-2||-2|0|10|||0|15|||1|331123|328511|4|0|45
502593613|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2017-02-28|Followup|2012-08-19|2012-10-10|Declined|Late||||||||3|2||1|2|2||||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|3|3|3.33|||||3|3|3||||2|2||||4|4||Yellow||Volunteer: Lost contact with child/agency|66.4||1|1|1|1|F|Black||16|No|Mother|28208|Two Parent|$35,000 to $39,999|Y|Yes||Relative|General Community||Match Support|F|Hispanic||26|28217|Bachelors Degree|Single|Service: Restaurant||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502594130|31|0|2|502601730|3|0|2|500547881|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|331242|322561|4|1|45
502666718|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2013-07-25|Followup|2012-08-19|2012-08-02|Complete|Early|4|3|2|2|3|3|2.83|4|2|2|1|1|4|2.33|21.46|2|1|3|2|1|4|2.17|2|3|3|1|2|3|2.33|-6.87|4|4|||4|4|4|4||3|2|4|3|3|5|4|3|3|3.75|-20|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|3|4|3.67|3|3|3|3|22.33|1|2|1.5|4|4|4|-62.5|1|1|1|1|0|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Child/Family: Unrealistic expectations|23.2||1|1|2|2|F|Black||16|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||38|28202|Masters Degree||Business: Clerical||7|0|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502667545|31|0|2|500932879|31|0|2|500548835|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7458|9|||1|331247|327460|4|3|45
502415267|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-19|2012-12-06|Baseline|2011-08-19|2011-09-19|Complete|Done|4|1|4|1|4|4|3|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|14.6||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$25,000 to $29,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28269|Some College|Single|Unknown||0|0|Radio|Media|Big|General Community||RTBM|277|60|598|500000170|500015820|502415705|31|0|1|502657931|31|0|1|500550917|2||-2||4|3|500005291|500005291|-2||-2|0|5|||131|1|||1|331255|-1|4|3|44
502245129|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-22|NaT|Baseline|2011-08-19|2011-08-22|Complete|Done|4|3|4|2|3|3|3.17|||||||||1|4|3|2|4|3|2.83|||||||||4|3|2|3||||||5|4|3|2|3.5|||||||4|3|4|3|2|4|3|3.29||||||||||4|4|3|3.67||||||4|3|3.5|||||1|1||||4|4||||Green|Amachi||66.8||1|1|1|1|M|Multi-race (Black & Hispanic)||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||28|28262|High School Graduate|Single|Laborer||0|8|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|502245570|38|0|1|502670839|31|0|1|500551050|2||-2||2|1|500000294||-2||-2|0|10|||7671|13|||1|331272|-1|4|3|44
500826603|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2012-11-08|Followup|2012-08-19|2012-11-03|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|14.7||3|3|2|2|F|Black||16|No|Mother|28226|Two Parent|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|F|Black||39|28105|Masters Degree|Single|Business: Mgt, Admin|28204|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|500826861|31|0|2|501004437|31|0|2|500548053|2||-2||4|3|||-2||-2|0|5|||46|2|||1|331306||4|0|45
502619926|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-09|2015-05-05|Followup|2012-08-09|2012-08-17|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Volunteer: Lost contact with child/agency|44.8||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||38|28205|Bachelors Degree|Single|Law: Lawyer|28202|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502620542|31|0|2|502642260|1|0|2|500548116|2||500004641||4|1|500004640||-2||-2|0|10|||7464|9|||1|331428||4|3|45
502273093|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-01|2015-03-31|Followup|2011-10-01|2011-12-16|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|53.9||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||37|28277|PHD|Single|Medical: Healthcare Worker||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502273525|31|0|2|502252422|31|0|2|500471568|2||-2||4|1|||-2|500000294|-2|0|4|||7496|10|||1|331513||4|0|45
500465511|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-21|2013-10-31|Followup|2012-08-21|2012-09-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Graduated|86.3||1|1|1|1|M|Black||21|Yes|Mother|28262|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|M|White||54|28210|Masters Degree|Married|Finance: Accountant||0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500527675|1|0|1|500118120|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|4|||2230|7|||1|331663||4|1|45
500465506|BBBS of Greater Charlotte|Main Office|C|Active|2006-08-21|NaT|Followup|2012-08-21|2012-10-01|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi||126.8||1|1|1|1|M|Black||16|Yes|Mother|28262|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||54|28226|Bachelors Degree|Married|Arts, Entertainment, Sports||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500496966|1|0|1|500118121|2||500003586||2|2|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|331664||4|3|45
501691220|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-02|2012-08-29|Followup|2012-07-02|2012-07-31|Complete|Done|3|3|4|4|3|3|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child/Family: Moved|37.9||1|1|2|3|M|White||15|No|Mother|27949|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree||Business: Marketing|28031|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|501691558|1|0|1|501721806|1|0|1|500367645|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|331706||4|3|45
500186435|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-23|2015-08-20|Followup|2012-07-23|2012-09-06|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|144.9||1|1|1|1|M|Black||20||Mother|28216|One Parent: Female|Unknown||No|Brochure|Media|General Community||Match Support|M|White||45|28226|Bachelors Degree|Married|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187988|31|0|1|500189358|1|0|1|500037395|2||-2||4|1|||-2||-2|51|1|||7496|10|||1|331709||4|1|45
502245129|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-22|NaT|Followup|2012-08-22|2012-11-06|Expired|Late||||||||4|3|4|2|3|3|3.17|||||||||1|4|3|2|4|3|2.83||||||4|3|2|3|||||||5|4|3|2|3.5||||||||||4|3|4|3|2|4|3|3.29||||||4|4|3|3.67|||||4|3|3.5||||1|1||||4|4||Green|Amachi||66.8||1|1|1|1|M|Multi-race (Black & Hispanic)||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||28|28262|High School Graduate|Single|Laborer||0|8|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|502245570|38|0|1|502670839|31|0|1|500551050|2||-2||2|1|500000294||-2||-2|0|10|||7671|13|||1|331819|331272|4|0|45
502000252|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-22|NaT|Followup|2012-08-22|2012-10-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||78.8||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020910|502000651|31|0|1|502127058|1|0|1|500465318|2||-2||2|1|||-2||-2|0|10|||130|1|||1|331855||4|1|45
500474486|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-23|2015-08-18|Followup|2012-08-23|2012-10-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|107.8||1|1|1|1|M|Black||20||Mother|28214|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||38|28209|Bachelors Degree|Single|Construction|28247|0|2|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500474735|31|0|1|500491064|31|0|1|500118168|2||-2||4|3|||-2||-2|34|2|||7447|3|||1|331858||4|1|45
502234504|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-28|NaT|Followup|2012-07-28|2012-09-05|Complete|Done|3|2|3|2|3|3|2.67|4|4|4|4|2|4|3.67|-27.25|2|3|4|2|3|4|3|1|4|4|1|2|4|2.67|12.36|4|4|4|4|4|4|4|4|0|3|4|4|4|3.75|3|3|5|5|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|3|3|3|1|3|2|50|2|2|2|2|0|4|4||||Yellow|Project Big||79.6||1|1|2|2|F|Black||16|No|GrandMother|28208|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|Project Big|Match Support|F|Black||37|28216|Bachelors Degree|Single|Customer Service||8|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500008321|502234935|31|0|2|502129464|31|0|2|500463451|2||500004641||2|2|500004640|500004640|-2||-1|0|4|||11247|3|1204|3|1|332243|155881|4|3|45
501318837|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-04|2013-02-27|Followup|2012-08-04|2012-08-20|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|30.8||2|2|1|1|M|Black||17|No|Mother|28205|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Retail: Sales||0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|501319115|31|0|1|502170420|1|0|1|500459741|2||-2||4|3|||-2||-2|6854|8|||7496|10|||1|332263||4|1|45
502183420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-28|2015-01-15|Followup|2011-09-28|2011-10-10|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|4|4|4|4|||||||||3|3|3|3||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Time constraint|51.6||2|2|1|1|M|Multi-race (Black & White)||14|Yes|GrandMother|28215|Grandparents|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||58|28226|Masters Degree|Married|Tech: Sales, Mktg|28202|6|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502183840|36|0|1|502264770|1|0|1|500473793|2||500003586||4|2|500000294|500000294|-2||-2|7016|11|||7464|9|||1|332762||4|3|45
502615628|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-09|2011-12-28|Baseline|2011-08-25|2011-09-09|Complete|Done|3|2|2|1|3|2|2.17|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|||||||2|2||||4|4||||Green||Volunteer: Time constraint|3.6||1|1|2|2|M|Black||16|No|Mother|28215|One Parent: Female|$10,000 to $14,999||Yes||Therapist/Counselor|General Community||RTBM|M|Black||27|28262|Associate Degree|Divorced|Medical: Nurse|28203|1|0|Self|Self|Big|General Site||Match Support|277|60|598|500000170|500001281|502616240|31|0|1|502635965|31|0|1|500551985|2||-2||4|1|||-2||-1|0|5|||7464|9|||1|333011|-1|4|3|44
501457406|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-20|2013-07-16|Followup|2012-08-20|2012-10-10|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|46.9||1|1|1|1|M|Black||21|No|Mother|28269|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28205|||Finance: Banking|28217|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|501457691|31|0|1|501720969|1|0|1|500375964|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|333287||4|1|45
501529924|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2017-02-28|Followup|2012-08-27|2012-10-10|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|78.1||2|2|1|1|F|Black||15|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||30|28209|Bachelors Degree|Single|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501530213|31|0|2|502199360|1|0|2|500465517|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|333289||4|1|45
502636177|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-29|2013-09-19|Followup|2012-08-29|2012-08-28|Complete|Done|4|3|4|1|4|4|3.33|4|1|4|1|4|3|2.83|17.67|4|4|4|4|4|4|4|4|4|4|4|3|4|3.83|4.44|4|4|4|4|4|4|4|4|0|5|5|5|5|5|4|4|4|4|4|25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Moved|24.7||1|1|1|1|F|Black||14|No|GrandMother|28216|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|Black||30|28212||Single|Medical||0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502636872|31|0|2|502643313|31|0|2|500551053|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|333720|330694|4|3|45
502097843|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-29|2016-08-11|Followup|2012-08-29|2012-08-23|Complete|Done|2|3|3|3|3|3|2.83|3|2|2|1|4|3|2.5|13.2|3|4|4|3|3|4|3.5|2|3|3|2|3|3|2.67|31.09|4|4|4|4|4|4|4|4|0|4|4|4|5|4.25|3|3|3|4|3.25|30.77|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3|3|3|33.33|3|3|3|3||||2|2|2|2|0|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child: Lost interest|59.4||1|1|2|2|M|Black||17|No|Mother|28078|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500021785|502098263|31|0|1|502643791|3|0|1|500550390|2||-2||4|1|500005291||-2||-2|0|10|||7496|10|||1|333817|330290|4|3|45
502630686|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2014-08-06|Baseline|2011-08-29|2011-09-02|Complete|Done|3|4|3|1|1|3|2.5|||||||||2|3|4|4|3|3|3.17|||||||||1|4|3|2.67||||||3|2|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Yellow|Amachi, Project Big AND Amachi|Volunteer: Lost contact with child/agency|35.1||1|1|1|1|M|Black||16|Yes|Mother|28216|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Multi-race (Black & Hispanic)||39|28208|Bachelors Degree|Single|Business: Marketing||1|6|Recruitment Event|BBBS Board/Staff|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500015820|502631341|31|0|1|502630052|38|0|1|500552346|2||500003586||4|2|500000294, 500004901|500000294|-2|500005291|-2|0|5|||7462|13|||1|333868|-1|4|3|44
502602958|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-11|2017-02-23|Baseline|2011-08-29|2011-09-11|Complete|Done|4|1|1|2|3|4|2.5|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|65.4||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||52|28207|Masters Degree|Married|Business|28202|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501480402|31|0|1|502578040|1|0|1|500552390|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|333955|-1|4|3|44
500761491|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2013-03-22|Followup|2012-08-27|2012-09-05|Complete|Done|4|3|4|2|3|3|3.17|||||||||4|3|3|2|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|30.8||3|3|1|1|F|Black||16||Aunt|28213|One Parent: Female|$40,000 to $44,999|Y|No||Self|General Community||Enrollment|F|Black||61|28269|Bachelors Degree|Divorced|Education: Teacher|28215|1|1|LPL Financial|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500761759|31|0|2|502189613|31|0|2|500465204|2||-2||4|1|||-2||-2|0|10|||11247|3|||1|334025||4|3|45
502670076|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-12|2013-06-06|Baseline|2011-08-30|2011-10-12|Complete|Done|4|4|3|4|3|4|3.67|||||||||3|4|4|2|2|4|3.17|||||||||3|3|2|2.67||||||5|3|4|3|3.75|||||||4|3|4|4|4|4|3|3.71||||||||||3|3|3|3||||||4|3|3.5|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|19.8||2|2|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|Black||31|29223|||Human Services: Youth Worker||0|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502670904|31|0|2|502655392|31|0|2|500552412|2||-2||4|2||500000294, 500016374|-2||-2|0|10|||7459|10|||1|334127|-1|4|3|44
502619301|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-21|2012-07-31|Baseline|2011-08-31|2011-09-21|Complete|Done|3|2|4|3|2|4|3|||||||||2|3|3|3|4|4|3.17|||||||||2|2|2|2||||||5|2|4|4|3.75|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|4|3.67||||||4|2|3|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|10.3||1|1|1|1|F|Hispanic||15|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||RTBM|F|Hispanic||34|28078|Some College|Single|Education: Teacher|28269|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502619917|3|0|2|502590110|3|0|2|500552773|2||500003586||4|3|500005291||-2|500004640|-2|0|10|||7462|13|||1|334718|-1|4|3|44
502307352|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-31|2013-02-28|Followup|2012-08-31|2012-10-15|Declined|Done||||||||3|3|3|3|3|3|3|||||||||3|3|3|3|3|3|3||||||3|4|3|3.33|||||||3|4|3|3|3.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|3|3||||1|1|||||||Red|Amachi, Project Big AND Amachi|Volunteer: Lost contact with child/agency|18||2|2|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big AND Amachi|Match Support|F|Black||33|28217|PHD|Single|Medical: Doctor, Provider||0|0|Recruitment Event|Other Big|Big|General Community||Match Support|277|60|598|500000170|500015820|502307784|31|0|2|502636073|31|0|2|500552236|2||500004772||4|3|500000294, 500004901|500004901|-2||-2|0|4|||7460|12|||1|334754|196663|4|1|45
501776333|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-08|2013-07-25|Followup|2012-09-08|2012-10-23|Complete|Done|4|3|4|2|4|3|3.33|3|2|3|2|4|4|3|11|2|3|4|2|2|4|2.83|3|3|3|2|3|3|2.83|0|4|4|3|3.67|3|3|3|3|22.33|3|4|3|3|3.25|4|4|4|4|4|-18.75|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Green||Volunteer: Moved|46.5||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28210|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011746|501776688|31|0|1|501832599|31|0|1|500381636|2||-2||4|1|||-2|500000294|-2|34|2|||7464|9|||1|334791|9814|4|3|45
502601023|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-31|2016-08-11|Followup|2012-08-31|2012-11-15|Expired|Late||||||||3|2|3|1|3|4|2.67|||||||||3|3|4|2|2|3|2.83||||||4|4|4|4|||||||3|3|4|5|3.75||||||||||4|2|4|4|3|4|3|3.43||||||3|4|2|3|||||3|3|3||||2|2||||4|4||Green|2010-2012 OJJDP JJI|Child: Graduated|59.4||1|1|1|1|F|Black||19||Mother|28216|Two Parent|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||51|28277|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502601540|31|0|2|502546883|1|0|2|500550809|2||-2||4|1|500005291|500005291|-2||-2|6854|8|||7464|9|||1|335061|331012|4|0|45
502627470|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-12|2014-05-19|Baseline|2011-09-01|2011-09-12|Complete|Done|4|4|4|3|2|4|3.5|||||||||2|2|4|1|4|4|2.83|||||||||3|4|4|3.67||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|32.2||1|1|1|1|M|Hispanic|Mexican|16|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|Asian||26|28105|Some College|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502628116|3|10|1|502672424|4|0|1|500552887|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|335186|-1|4|3|44
501872144|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-30|NaT|Followup|2012-07-30|2012-10-14|Expired|Late||||||||4|4|3|1|3|3|3|||||||||2|3|2|1|2|2|2||||||2|3|2|2.33|||||||2|2|1|2|1.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||1|1|1||||2|2|||||||Green|||79.5||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown|Y|Yes||Relative|General Community||Match Support|M|White||35|28205|Masters Degree|Married|Tech: Engineer|28115|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501872517|31|31|1|502063676|1|0|1|500460156|2||-2||2|1|||-2||-2|0|3|||46|2|||1|335198|155585|4|0|45
502668768|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-17|2012-11-13|Baseline|2011-09-01|2011-09-17|Complete|Done|3|4|1|2|1|1|2|||||||||2|1|3|1|1|3|1.83|||||||||3|3|3|3||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||1|4|2.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|13.9||1|1|1|1|F|Hispanic||15|No|Mother|28212|One Parent: Female|$10,000 to $14,999||Yes||School|General Community||Match Support|F|Hispanic||30|28226|Bachelors Degree|Married|Law: Paralegal|28226|4|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502669595|3|0|2|502571563|3|0|2|500552927|2||-2||4|2|||-2||-2|0|4|||7462|13|||1|335238|-1|4|3|44
502436202|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2015-07-13|Followup|2012-09-02|2012-10-24|Declined|Late||||||||3|2|2|1|3|3|2.33|||||||||3|3|3|4|2|4|3.17||||||4|4|4|4|||||||2|5|5|5|4.25||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||2|4|3||||1|1||||4|4||Green||Child: Graduated|46.3||1|1|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|Masters Degree|Single|Finance: Banking||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502436645|31|0|1|502642999|1|0|1|500549046|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|335452|327937|4|1|45
502630686|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2014-08-06|Followup|2013-09-02|2013-10-09|Complete|Done|4|4|4|4|4|4|4|3|4|3|1|1|3|2.5|60|4|4|4|4|3|4|3.83|2|3|4|4|3|3|3.17|20.82|4|4|4|4|1|4|3|2.67|49.81|3|4|3|3|3.25|3|2|2|3|2.5|30|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|2|2|2|100|1|1|1|1|0|4|4|4|4|0|Yellow|Amachi, Project Big AND Amachi|Volunteer: Lost contact with child/agency|35.1||1|1|1|1|M|Black||16|Yes|Mother|28216|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Multi-race (Black & Hispanic)||39|28208|Bachelors Degree|Single|Business: Marketing||1|6|Recruitment Event|BBBS Board/Staff|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500015820|502631341|31|0|1|502630052|38|0|1|500552346|2||500003586||4|2|500000294, 500004901|500000294|-2|500005291|-2|0|5|||7462|13|||1|335457|333868|4|3|45
502697677|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2013-03-27|Followup|2012-09-02|2012-08-24|Complete|Done|3|3|3|2|3|4|3|4|3|3|3|3|3|3.17|-5.36|2|3|3|2|3|4|2.83|2|4|3|3|2|4|3|-5.67|4|4|4|4|4|4|4|4|0|2|4|4|3|3.25|5|5|4|2|4|-18.75|4|4|4|4|3|4|2|3.57|4|4|4|3|4|4|2|3.57|0|4|3|2|3|3|3|4|3.33|-9.91|3|2|2.5|3|3|3|-16.67|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Moved|18.8||1|1|1|1|F|Hispanic||19|No|Mother|28027|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|F|White||32|28027|Bachelors Degree|Single|Business: Marketing|28075|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502605848|3|0|2|502590370|1|0|2|500550704|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|335531|330902|4|3|45
502549830|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-30|NaT|Followup|2012-06-30|2012-07-02|Complete|Done|4|1|2|1|2|4|2.33|||||||||1|4|4|1|1|4|2.5|||||||||2|4|4|3.33||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||68.5||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|Amachi, Project Big, Project Big AND Amachi|Match Support|M|Black||25|28211||Single|Transport: Driver||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|1|502462453|31|0|1|500538768|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-1||-2|0|4|||7464|9|||1|335613||4|3|45
502254067|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-10|2013-01-03|Followup|2012-09-10|2012-08-29|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|1|1|1|1|1|1.5|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|27.8||3|3|1|1|F|Black||14|No|Mother|28209|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|Black||37|28210|Bachelors Degree|Single|Insurance||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502254499|31|0|2|502214352|31|0|2|500466835|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|335863||4|3|45
501261979|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-22|2014-10-13|Followup|2012-07-22|2012-08-13|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|74.7||1|1|3|3|F|Black||15|No|Mother|28134|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||55|28173||Married|Human Services: Non-Profit|28205|0|0|Coworker|Workplace Partner|Big|General Community|VOL - Maximizing Match Impact|Match Support|277|60|598|500000170|500011349|501262256|31|0|2|500418936|31|0|2|500278634|2||-2||4|1|||-2|500011314|-2|0|10|||7447|3|||1|335875||4|3|45
502108064|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2014-02-06|Followup|2012-07-22|2012-09-07|Declined|Late||||||||3|4|4|4|4|4|3.83|||||||||1|4|3|1|1|3|2.17||||||4|4|4|4|||||||5|5|5|5|5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||1|1|1||||1|1|||||||Yellow||Child: Graduated|42.5||1|1|1|1|F|White||21|No|Father|28277|One Parent: Male|Unknown||No||Relative|General Community||Match Support|F|White||48|28277|High School Graduate|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502108491|1|0|2|502146885|1|0|2|500460150|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|335877|155579|4|1|45
500881634|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-14|NaT|Followup|2012-07-14|2012-08-23|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|4|3|3|4|4|3.5|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||104||1|2|1|2|M|Black||18||Mother|28213|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||38|28213||Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500881903|31|0|1|500816190|31|0|2|500277615|2||-2||2|1|||-2||-2|0|4|||46|2|||1|335926||4|3|45
502455004|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-20|NaT|Baseline|2011-09-06|2011-09-20|Complete|Done|4|2|4|1|1|4|2.67|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||4|2|3|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI||65.8||1|1|1|1|M|Black|Other African|15|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|29720|Bachelors Degree|Married|Business: Sales|28134|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|31|1|502680045|1|0|1|500553363|2||-2||2|1|500005291|500005291|-2||-2|0|4|||7464|9|||1|336027|-1|4|3|44
500970495|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-10|2017-03-09|Followup|2012-09-10|2012-10-24|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|101.9||3|3|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$35,000 to $39,999||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black|Other African|44|28212||Single|Consultant||1|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500970766|31|0|2|500965698|31|31|2|500285645|2||-2||4|2|||-2||-2|7294|13|||46|2|||1|336064||4|1|45
501597228|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-04|NaT|Followup|2012-09-04|2012-10-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||90.3||1|1|1|1|F|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||40|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28204|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501597548|31|0|2|501397328|31|0|2|500379964|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|336211||4|1|45
500186675|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-23|2013-08-29|Followup|2012-08-23|2012-08-07|Complete|Early|4|1|2|1|4|4|2.67|||||||||2|3|4|2|2|3|2.67|||||||||4|4|4|4||||||4|5|3|4|4|||||||3|4|4|4|4|4|4|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|72.2||4|4|1|1|F|Black||20|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||38|28221||Single|Human Services: Youth Worker||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188055|31|0|2|500865601|31|0|2|500185332|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|336300||4|3|45
501825910|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-24|2016-09-23|Followup|2012-08-24|2012-08-14|Complete|Done|3|4|3|3|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|3|3.67||||||5|4|5|3|4.25|||||||4|4|3|4|3|4|3|3.57||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|85||1|1|1|1|M|Black||16|Yes|Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|White||51|28214|Masters Degree|Married|Business: Sales|94108|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|501196986|1|0|1|500380446|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||7496|10|||1|336304||4|3|45
500961274|BBBS of Greater Charlotte|Main Office|C|Active|2007-08-27|NaT|Followup|2012-08-27|2012-10-02|Complete|Done|4|1|4|1|4|4|3|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi||114.6||1|1|2|2|F|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28216|Bachelors Degree|Divorced|Business: Clerical|28204|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500934638|31|0|2|500403000|31|0|2|500186952|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|336306||4|3|45
500185972|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-01|2012-12-21|Followup|2012-09-01|2012-08-27|Complete|Done|3|2|2|2|1|4|2.33|||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|3|3|||||1|1||||4|4||||Green|Amachi|Child: Graduated|75.7||2|3|1|1|F|Black||22|Yes|Mother|28206|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|F|Black||38|28213|Bachelors Degree|Single|Education: Teacher|28202|2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187610|31|0|2|500492482|31|0|2|500120588|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|336311||4|3|45
501831581|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-29|NaT|Followup|2012-09-29|2012-09-04|Complete|Early|4|2|4|4|4|2|3.33|||||||||2|2|3|4|1|3|2.5|||||||||4|4|4|4||||||3|2|2|2|2.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Green|Amachi||89.5||1|1|2|3|F|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||38|28273||Single|Tech: Engineer||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501831944|31|0|2|500715453|31|0|2|500387624|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|336598||4|3|45
501305368|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-09|2013-06-19|Followup|2012-09-09|2012-08-02|Complete|Early|4|4|4|4|4|4|4|||||||||3|4|4|4|2|4|3.5|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2||||4|4||||Green||Volunteer: Moved|21.3||2|2|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|M|White||29|28202|Bachelors Degree|Single|Finance: Banking|28202|0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|501305646|31|0|1|502665365|1|0|1|500552025|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|336870||4|3|45
502696388|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-27|2012-03-23|Baseline|2011-09-09|2011-09-27|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|3|3|4|4|4|3.67|||||||||4|4|4|4||||||5|4|5|3|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Moved|5.8||1|1|1|1|F|Black||17|No|Mother|28212|One Parent: Female|Unknown|Y|Yes||Self|General Community||RTBM|F|White||28|28105|Masters Degree|Single|Medical: Healthcare Worker|28078|0|1|Recruitment Event|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008629|502697233|31|0|2|502609046|1|0|2|500553973|2||-2||4|1|500005291||-2||-2|0|10|||7460|12|||1|336951|-1|4|3|44
502602958|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-11|2017-02-23|Followup|2012-09-11|2012-10-23|Complete|Done|4|3|3|2|3|4|3.17|4|1|1|2|3|4|2.5|26.8|2|4|4|2|3|3|3|4|3|4|4|4|4|3.83|-21.67|4|4|||4|4|4|4||3|4|3|3|3.25|5|3|5|5|4.5|-27.78|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|4|4|4|2|3|2.5|60|2|2|2|2|0|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|65.4||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||52|28207|Masters Degree|Married|Business|28202|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501480402|31|0|1|502578040|1|0|1|500552390|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|337265|333955|4|3|45
500185624|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-28|2013-02-26|Followup|2012-06-28|2012-07-10|Complete|Done|4|4|4|1|3|4|3.33|||||||||4|3|4|2|4|3|3.33|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Yellow|Amachi|Child/Family: Moved|68||1|1|1|1|M|Black||16|Yes|Mother|28213|Other/Unknown|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||61|28205||Married|Tech: Management||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|500187258|31|0|1|500923420|31|0|1|500182113|2||500003586||4|2|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|337329||4|3|45
502538068|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-27|2012-01-31|Baseline|2011-09-12|2011-09-27|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|4.1||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||28|28215||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|502538521|31|0|1|502672354|1|0|1|500554099|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|337368|-1|4|3|44
502627470|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-12|2014-05-19|Followup|2012-09-12|2012-09-17|Complete|Done|4|2|3|3|3|3|3|4|4|4|3|2|4|3.5|-14.29|2|4|3|2|3|3|2.83|2|2|4|1|4|4|2.83|0|4|4|4|4|3|4|4|3.67|8.99|4|3|3|2|3|4|5|3|4|4|-25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|4|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Lost contact with child/agency|32.2||1|1|1|1|M|Hispanic|Mexican|16|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|Asian||26|28105|Some College|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502628116|3|10|1|502672424|4|0|1|500552887|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|337434|335186|4|3|45
501309634|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-12|NaT|Followup|2012-09-12|2012-10-24|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||102.1||1|1|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||46|27704|Associate Degree|Divorced|Medical: Admin||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501309912|31|0|2|501046221|31|0|2|500281317|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7462|13|||1|337835||4|1|45
500186665|BBBS of Greater Charlotte|Main Office|C|Completed|2004-07-20|2013-02-28|Followup|2012-07-20|2012-08-30|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|103.3||1|1|1|1|M|Black||21||Mother|28202|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|Black||40|28207||Single|Medical: Nurse||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500188050|31|0|1|500189566|31|0|1|500037664|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|337859||4|1|45
502172536|BBBS of Greater Charlotte|Main Office|C|Active|2010-10-13|NaT|Followup|2012-10-13|2012-10-05|Complete|Done|3|4|4|4|4|4|3.83|3|2|4|3|1|1|2.33|64.38|2|4|4|2|4|4|3.33|2|4|4|2|2|4|3|11|4|4|4|4|4|4|4|4|0|5|5|4|5|4.75|5|4|4|4|4.25|11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|2|3|0|2|2|2|2|0|4|4||||Green|||77.1||1|1|1|1|F|Black||17|No|Mother|28269|Two Parent|Unknown||Yes||Relative|General Community||Match Support|F|Multi-race (Asian & White)||33|28205|Masters Degree|Married|Finance: Economist|28223|7|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502172965|31|0|2|501279665|37|0|2|500475431|2||-2||2|1|||-2||-2|0|3|||129|1|||1|338103|184611|4|3|45
502359051|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-28|2017-02-28|Followup|2011-10-28|2012-01-05|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|76.1||1|1|1|1|F|Black||14|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||35|28213|Masters Degree|Married|Business: Clerical||3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502359489|31|0|2|502242295|31|0|2|500483954|2||500004772||4|3|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|10|||131|1|||1|338144||4|1|45
501614157|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-29|2013-04-04|Followup|2012-07-29|2012-10-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|44.2||1|1|1|1|F|Black||21|No|Mother|28202|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28273|||Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|501614477|31|0|2|501596246|31|0|2|500374258|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|338406||4|0|45
500934906|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-31|2013-02-12|Followup|2012-07-31|2012-10-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Lost contact with child/agency|66.5||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||52|28216|Bachelors Degree|Married|Tech: Engineer||13|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500935173|31|0|2|500859806|31|0|2|500186448|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|338415||4|0|45
502569411|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-14|2012-12-19|Followup|2012-09-14|2012-09-04|Complete|Done|2|2|4|2|3|2|2.5|4|4|4|2|3|4|3.5|-28.57|2|4|2|1|2|4|2.5|2|3|3|1|2|3|2.33|7.3|4|3|3|3.33|4|4|4|4|-16.75|5|3|4|2|3.5|5|3|3|4|3.75|-6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|4|4|4|4|-25|2|4|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Yellow|Amachi, 2010-2012 OJJDP JJI|Child/Family: Time constraints|15.2||1|1|1|1|F|American Indian or Alaska Native||14|Yes|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||45|28027|||Medical: Nurse|28144|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502569865|6|0|2|502642653|1|0|2|500550403|2||500003586||4|2|500000294, 500005291|500005291|-2||-2|0|10|||7496|10|||1|338526|330300|4|3|45
502229042|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-30|2013-02-22|Followup|2012-09-30|2012-10-11|Complete|Done|4|2|4|1|4|4|3.17|||||||||2|4|4|4|1|4|3.17|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|28.8||3|3|1|1|F|Black||14|No|Mother|28269|Two Parent|Unknown||Yes||Relative|General Community||Match Support|F|White||35|28211||Single|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502172965|31|0|2|502272069|1|0|2|500470500|2||-2||4|2|||-2|500000294|-2|0|3|||7496|10|||1|338624||4|3|45
500186106|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-18|2015-08-13|Followup|2012-10-18|2012-11-27|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|3|3|3|1|3|2.5|||||||||4|4|4|4||||||3|4|2|3|3|||||||4|3|4|4|3|3|2|3.29||||||||||3|4|3|3.33||||||2|4|3|||||2|2||||4|4||||Green||Child: Graduated|93.8||2|2|1|1|F|Black||20||Mother|28217|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||35|28211|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187698|31|0|2|500778380|1|0|2|500202993|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|338626||4|3|45
502062624|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-30|2012-12-19|Followup|2012-08-30|2012-08-29|Complete|Done|4|4|4|4|4|4|4|3|3|3|2|1|4|2.67|49.81|4|4|4|4|4|4|4|2|4|3|3|3|4|3.17|26.18|3|3|3|3|4|4|4|4|-25|4|5|5|5|4.75|3|5|3|5|4|18.75|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|4|4|4|4|-16.75|3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Yellow||Volunteer: Feels incompatible with child/family|27.7||1|1|1|1|F|Black||16|No|Mother|28081|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||32|28083|Bachelors Degree|Single|Tech: Computer/Programmer|28216|1|7|LPL Financial|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|502063048|31|0|2|502067861|31|0|2|500460279|2||-2||4|2|||-2||-2|0|10|||11247|3|||1|338690|155833|4|3|45
500480596|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-13|2014-01-16|Followup|2012-09-13|2012-08-31|Complete|Done|3|4|4|3|4|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|88.1||1|1|1|1|M|Black||21|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Married|Business: Sales|28203|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500480847|31|0|1|500491267|1|0|1|500120915|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|338742||4|3|45
501788776|BBBS of Greater Charlotte|Main Office|C|Active|2010-01-25|NaT|Followup|2012-01-25|2012-03-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||85.7||1|1|1|1|M|Black||14|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||64|28117||Married|Business: Sales|28031|0|0|Alpha Kappa Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500020752|501789128|31|0|1|501698382|1|0|1|500418170|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||8697|14|||1|339343||4|1|45
500896018|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-03|2014-08-14|Followup|2012-07-03|2012-06-18|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|4|1|4|4|3|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Child: Graduated|73.4||1|1|1|1|F|Black||20|Yes|Mother|28027|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||40|28027|Bachelors Degree|Separated|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500896288|31|0|2|501225232|31|0|2|500269506|2||-2||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|339360||4|3|45
502668768|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-17|2012-11-13|Followup|2012-09-17|2012-09-26|Declined|Done||||||||3|4|1|2|1|1|2|||||||||2|1|3|1|1|3|1.83||||||3|3|3|3|||||||4|4|4|3|3.75||||||||||4|4|4|4|4|4|4|4||||||3|4|4|3.67|||||1|4|2.5||||2|2||||4|4||Yellow||Volunteer: Time constraint|13.9||1|1|1|1|F|Hispanic||15|No|Mother|28212|One Parent: Female|$10,000 to $14,999||Yes||School|General Community||Match Support|F|Hispanic||30|28226|Bachelors Degree|Married|Law: Paralegal|28226|4|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502669595|3|0|2|502571563|3|0|2|500552927|2||-2||4|2|||-2||-2|0|4|||7462|13|||1|339370|335238|4|1|45
500399844|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-20|2017-02-24|Followup|2012-08-20|2012-10-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|114.2||1|2|1|2|F|Black||16||Mother|28208|One Parent: Female|Unknown||No||School|General Site||Match Support|F|White||35|28210|Bachelors Degree|Single|Business: Mgt, Admin|29715|0|0|Radio|Media|Big|General Site||Match Support|277|60|598|500000170|500008321|500400094|31|0|2|500188569|1|0|2|500190707|2||-2||4|3|||-1||-1|0|4|||131|1|||1|339374||4|1|45
501604446|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-19|NaT|Followup|2012-09-19|2012-10-24|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|2010-2012 OJJDP JJI||65.9||2|2|1|1|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28213|Bachelors Degree|Married|Tech: Support, Writing|28273|11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|502664359|31|0|1|500555050|2||-2||2|1|500005291|500005291|-2||-2|0|10|||7462|13|||1|339616||4|1|45
502415267|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-19|2012-12-06|Followup|2012-09-19|2012-10-09|Complete|Done|4|1|2|1|4|4|2.67|4|1|4|1|4|4|3|-11|2|4|3|2|1|3|2.5|2|4|4|2|4|4|3.33|-24.92|4|4|4|4|4|4|4|4|0|4|5|3|3|3.75|3|5|5|5|4.5|-16.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|14.6||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$25,000 to $29,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28269|Some College|Single|Unknown||0|0|Radio|Media|Big|General Community||RTBM|277|60|598|500000170|500015820|502415705|31|0|1|502657931|31|0|1|500550917|2||-2||4|3|500005291|500005291|-2||-2|0|5|||131|1|||1|339632|331255|4|3|45
500187090|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-04|2013-08-29|Followup|2012-10-04|2012-09-07|Complete|Early|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|82.8||2|2|3|3|F|Black||20||Mother|28216|Two Parent|Unknown||No||School|General Community||Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|500188103|31|0|2|500189320|31|0|2|500125754|2||-2||4|1|||-2|500016374|-2|0|4|||7464|9|||1|339639||4|3|45
500187075|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-21|2014-01-16|Followup|2012-09-21|2012-10-22|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|111.8||1|1|6|6|F|Black||21||Mother|28205|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||38|28209|Bachelors Degree|Single|Human Services: Non-Profit||0|0|Recruitment Event|Self|Big|General Site||Match Support|277|60|598|500000170|500012459|500188223|31|0|2|500189550|1|0|2|500037643|2||-2||4|1|||-2||-1|0|10|||7458|9|||1|339683||4|3|45
500267459|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-19|2013-02-27|Followup|2012-09-19|2012-12-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|77.3||1|1|1|1|M|Black||16||Mother|28203|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28202|Bachelors Degree|Single|Finance: Accountant||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|500187395|31|0|1|500464544|1|0|1|500121193|2||-2||4|3|||-2||-2|0|10|||46|2|||1|340059||4|0|45
502455004|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-20|NaT|Followup|2012-09-20|2012-09-18|Complete|Done|4|2|4|4|4|4|3.67|4|2|4|1|1|4|2.67|37.45|2|3|4|2|4|4|3.17|4|4|4|2|4|4|3.67|-13.62|4|4|4|4|4|4|4|4|0|5|5|3|4|4.25|5|5|4|5|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|3|4|3.5|4|2|3|16.67|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||65.8||1|1|1|1|M|Black|Other African|15|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|29720|Bachelors Degree|Married|Business: Sales|28134|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|31|1|502680045|1|0|1|500553363|2||-2||2|1|500005291|500005291|-2||-2|0|4|||7464|9|||1|340176|336027|4|3|45
502186245|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-18|2013-08-22|Followup|2012-08-18|2012-07-26|Complete|Early|3|2|2|2|3|3|2.5|||||||||2|4|4|3|4|4|3.5|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Volunteer: Moved|24.1||3|3|1|1|F|Black||14|No|Mother|28216|Two Parent|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|White||33|28203||Single|Business|28211|3|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500004169|501610196|31|0|2|502605983|1|0|2|500548277|2||500004641||4|1|500004640||-2|500000294, 500004640|-2|0|10|||7464|9|||1|340396||4|3|45
502436198|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-17|2012-10-31|Followup|2012-03-17|2012-05-01|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|19.5||2|2|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||51|28205|Masters Degree|Married|Education: Teacher|28212|14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502436641|31|0|2|502446619|1|0|2|500520591|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|340904||4|1|45
502240205|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-22|2014-06-11|Followup|2012-09-22|2012-11-30|Declined|Late||||||||4|2|4|3|3|3|3.17|||||||||2|3|3|2|2|3|2.5||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||4|2|3||||2|2|||||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|32.6||3|3|2|2|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||48|28203|Bachelors Degree|Married|Business: Mgt, Admin|28202|1|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002334|502240634|31|0|2|502657850|31|0|2|500553471|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|341039|156483|4|1|45
502670071|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-26|2014-03-20|Baseline|2011-09-22|2011-10-26|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Yellow|Amachi, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|28.8||1|1|1|1|F|Black||16|Yes|Mother|28083|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|Black||36|28269|Masters Degree|Single|Human Services: Youth Worker|28027|2|2|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|502670906|31|0|2|502685522|31|0|2|500557057|2||500003586||4|2|500000294, 500005291|500005291|-2||-2|0|10|||9229|13|||1|341113|-1|4|3|44
502206673|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-13|2015-06-23|Baseline|2011-09-22|2011-10-13|Complete|Done|3|2|3|2|3|4|2.83|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||4|5|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Red|Amachi|Child: Lost interest|44.3||1|1|1|1|M|Black||17|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||47|28216|Bachelors Degree|Married|Business: Engineer|28255|18|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500013781|502207102|31|0|1|502668179|1|0|1|500557233|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|341305|-1|4|3|44
502567552|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-07|2012-07-31|Followup|2012-06-07|2012-06-20|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|13.8||1|1|2|2|F|Hispanic||14|Yes|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community|Project Big AND Amachi|Match Support|277|60|598|500000170|500011746|502568002|3|0|2|502208867|31|0|2|500538510|2||500004772||4|3|500000294, 500004640, 500004901|500004640, 500004901|-2|500004901|-2|0|4|||7464|9|||1|341422||4|1|45
502698363|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-18|2013-12-06|Baseline|2011-09-23|2011-10-18|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|4|4|4|4|1|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Lost contact with child/agency|25.6||1|1|1|1|M|Black||18|Yes|GrandMother|28203|Grandparents|Unknown||Yes||Self|General Community|Amachi|Enrollment|M|Black||43|28208|Bachelors Degree|Single|Education|28217|0|0|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500015820|502699208|31|0|1|502641410|31|0|1|500557390|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7452|6|||1|341569|-1|4|3|44
500863413|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-23|2013-02-28|Followup|2012-09-23|2012-11-05|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Moved|17.2||2|2|2|2|M|White||18|No|Mother|28227|One Parent: Female|$25,000 to $29,999||No||School|General Community||Match Support|M|White||36|28226|Some College|Single|Business: Marketing||2|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500004169|500863682|1|0|1|502632871|1|0|1|500551916|2||-2||4|3|||-2||-2|0|4|||46|2|||1|341759||4|1|45
502404516|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-23|2013-06-19|Followup|2012-08-23|2012-07-31|Complete|Early|2|3|2|3|2|2|2.33|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Moved|21.9||1|1|1|1|M|White||14|No|Mother|28273|One Parent: Female|Unknown||No|Yahoo!|Web Link|General Community||Enrollment|M|White||49|19711|Bachelors Degree|Living w/ Significant Other|Business: Marketing|28278|15|2|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500004169|502404954|1|0|1|502624164|1|0|1|500548056|2||-2||4|3|||-2|500004640|-2|30|2|||7464|9|||1|341884||4|3|45
500382177|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-18|2015-08-25|Followup|2012-09-18|2012-10-24|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|107.2||1|1|2|2|M|Black||16||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||43|28215|Bachelors Degree|Single|Finance: Banking|28262|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|500382427|31|0|1|500188566|31|0|1|500122093|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|342184||4|1|45
502221847|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-27|NaT|Followup|2012-09-27|2012-09-05|Complete|Early|1|1|1|1|3|1|1.33|3|1|2|1|4|2|2.17|-38.71|3|4|4|4|4|4|3.83|4|4|4|2|4|4|3.67|4.36|4|4|4|4|4|4|4|4|0|4|3|5|5|4.25|5|4|5|5|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|2|2|1|1.67|3|4|4|3.67|-54.5|4|4|4|2|4|3|33.33|2|2|2|2|0|4|4||||Green|Amachi||65.6||2|2|1|1|F|Black||16|Yes|GrandMother|28213|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||24|28027|Some College|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502222278|31|0|2|502654877|31|0|2|500556560|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|343129|154081|4|3|45
500483980|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-01|2014-03-24|Followup|2012-09-01|2012-10-24|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|90.7||1|1|2|2|M|Black||21||Mother|28227|One Parent: Female|$10,000 to $14,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||71|28270||Single|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500484231|31|0|1|500423426|31|0|1|500120592|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|345084||4|1|45
501831576|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-30|2012-10-17|Followup|2012-09-30|2012-08-29|Complete|Early|3|4|4|2|4|4|3.5|4|4|4|3|3|4|3.67|-4.63|2|4|4|4|2|4|3.33|2|4|4|2|2|4|3|11|4|4|4|4|4|4|4|4|0|4|5|5|4|4.5|4|2|4|4|3.5|28.57|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|2|3|2.5|2|2|2|25|1|1|2|2|-50|4|4||||Yellow|Amachi|Volunteer: Unrealistic expectations|12.6||3|3|1|1|F|Black||18|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|White||26|28262|Some College|Single|Retail: Sales||0|6|UNCC|College Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501831944|31|0|2|502697749|1|0|2|500556209|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||9221|5|1208|5|1|345121|11655|4|3|45
501750507|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-30|2013-06-13|Followup|2012-09-30|2012-12-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Infraction of match rules/agency policies|20.4||2|2|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|Black||35|28212|Masters Degree|Single|Human Services: Social Worker|28204|2|5|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500015820|501750847|31|0|2|502275127|31|0|2|500557811|2||-2||4|3||500005291|-2|500004640|-2|0|10|||7464|9|||1|345165||4|1|45
502264006|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-22|2017-02-26|Followup|2012-09-22|2012-09-28|Complete|Done|3|2|2|3|3|3|2.67|2|1|3|1|2|3|2|33.5|3|4|4|4|3|4|3.67|1|3|2|2|1|3|2|83.5|4|4|4|4|4|4|4|4|0|4|3|5|4|4|4|2|3|4|3.25|23.08|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|3|3.33|20.12|4|4|4|4|3|3.5|14.29|2|2|1|1|100|4|4||||Red||Child: Lost interest|77.2||1|1|1|1|F|Hispanic||16|No|Mother|28211|One Parent: Female|Unknown||Yes|Spanish Print|Media|General Community||Match Support|F|Hispanic||38|28202|Bachelors Degree|Single|Tech: Engineer|28202|12|0|Big Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020753|502264438|3|0|2|502274748|3|0|2|500470897|2||-2||4|3|||-2||-2|7063|1|||7456|8|||1|345620|178842|4|3|45
501771263|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-02-28|Followup|2012-09-29|2012-11-05|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|89||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||31|28262|Bachelors Degree|Single|Medical: Admin|28216|0|8|Recruitment Event|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501741899|31|0|2|501622704|31|0|2|500379993|2||-2||4|1|||-2||-2|0|10|||7443|2|||1|345706||4|1|45
501645192|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-21|2016-08-19|Followup|2012-07-21|2012-07-21|Complete|Done|3|4|4|4|3|4|3.67|||||||||2|3|4|3|3|3|3|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red||Child: Graduated|85||1|1|2|2|M|Hispanic||19|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501645515|3|0|1|501519306|1|0|1|500374818|2||-2||4|3||500016374|-2|500016374|-2|0|10|||7464|9|||1|346686||4|3|45
502241349|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2013-09-04|Followup|2012-07-22|2012-10-06|Expired|Late||||||||2|2|2|1|2|2|1.83|||||||||2|3|3|3|3|3|2.83||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Child/Family: Moved|37.5||1|1|2|2|M|Black||19|No|Aunt|28081|Two Parent|Unknown||No|Other|Faith Organization|General Community||Match Support|M|Black||54|28025||Married|Clergy|28025|23|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500002335|502241780|31|0|1|502240986|31|0|1|500461089|2||-2||4|1|||-2|500016374|-2|5635|9|||7671|13|||1|347619|157252|4|0|45
500930976|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-13|2013-04-26|Followup|2012-08-13|2012-09-25|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green||Child: Lost interest|56.4||1|1|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|Y|No||Service Organization|General Community||Match Support|F|Black||66|28205|Masters Degree|Single|Self-Employed, Entrepreneur||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500931243|31|0|2|501176751|31|0|2|500280106|2||-2||4|1|||-2||-2|0|11|||46|2|||1|347643||4|3|45
502499851|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2015-07-07|Baseline|2011-10-07|2011-11-11|Complete|Done|3|1|1|1|2|2|1.67|||||||||4|4|4|2|2|4|3.33|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|4|3|||||2|2||||4|4||||Red||Agency: Concern with Volunteer re: child safety|43.8||1|1|1|1|M|White||18|No|Mother|28210|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||39|28210|Masters Degree|Single|Finance|28106|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|502500300|1|0|1|502690262|1|0|1|500562789|2||-2||4|3|||-2||-2|0|10|||46|2|||1|348364|-1|4|3|44
501332658|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-01-19|Followup|2012-09-29|2012-09-25|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Severity of challenges|87.7||1|1|1|1|M|Black||15|Yes|GrandMother|28213|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||46|28227|High School Graduate|Single|Medical: Healthcare Worker|28269|4|0|Coworker|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500020752|501332937|31|0|1|501814288|1|0|1|500384166|2||-2||4|1|500000294|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||7447|3|||1|348991||4|3|45
502183420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-28|2015-01-15|Followup|2012-09-28|2012-12-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Time constraint|51.6||2|2|1|1|M|Multi-race (Black & White)||14|Yes|GrandMother|28215|Grandparents|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||58|28226|Masters Degree|Married|Tech: Sales, Mktg|28202|6|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502183840|36|0|1|502264770|1|0|1|500473793|2||500003586||4|2|500000294|500000294|-2||-2|7016|11|||7464|9|||1|348997||4|0|45
501811375|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-27|2013-08-28|Followup|2012-07-27|2012-07-16|Complete|Done|4|4|4|2|3|4|3.5|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||4|2|3|||||2|2||||4|4||||Yellow||Child: Graduated|49.1||1|1|3|3|F|Black||21|No|Mother|28027|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||41|28027|PHD|Single|Medical: Doctor, Provider|28075|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|501811730|31|0|2|501391123|31|0|2|500374230|2||-2||4|2|||-2|500016374|-2|0|8|||7464|9|||1|349458||4|3|45
502698998|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2014-03-13|Baseline|2011-10-12|2011-11-11|Complete|Done|3|2|2|1|3|3|2.33|||||||||3|2|3|3|3|3|2.83|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|28||1|1|1|1|F|Black||18|No|GrandMother|28211|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28203|Masters Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500012459|502699843|31|0|2|502692148|1|0|2|500564380|2||-2||4|2||500005291|-2||-2|0|4|||7464|9|||1|350301|-1|4|3|44
502670076|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-12|2013-06-06|Followup|2012-10-12|2012-09-25|Complete|Early|4|3|3|3|4|4|3.5|4|4|3|4|3|4|3.67|-4.63|3|4|4|2|3|4|3.33|3|4|4|2|2|4|3.17|5.05|3|4|4|3.67|3|3|2|2.67|37.45|5|4|3|4|4|5|3|4|3|3.75|6.67|4|4|4|4|4|4|4|4|4|3|4|4|4|4|3|3.71|7.82|2|4|1|2.33|3|3|3|3|-22.33|4|4|4|4|3|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Lost contact with child/agency|19.8||2|2|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|Black||31|29223|||Human Services: Youth Worker||0|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502670904|31|0|2|502655392|31|0|2|500552412|2||-2||4|2||500000294, 500016374|-2||-2|0|10|||7459|10|||1|350716|334127|4|3|45
502206673|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-13|2015-06-23|Followup|2012-10-13|2012-10-09|Complete|Done|3|4|4|1|1|4|2.83|3|2|3|2|3|4|2.83|0|2|4|3|4|2|3|3|2|3|3|3|3|3|2.83|6.01|4|4|4|4|4|4|4|4|0|4|5|4|3|4|4|5|3|3|3.75|6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Red|Amachi|Child: Lost interest|44.3||1|1|1|1|M|Black||17|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||47|28216|Bachelors Degree|Married|Business: Engineer|28255|18|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500013781|502207102|31|0|1|502668179|1|0|1|500557233|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|350896|341305|4|3|45
502638767|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-27|2012-06-29|Baseline|2011-10-13|2011-10-27|Complete|Done|4|4|4|3|3|4|3.67|||||||||4|4|3|4|1|3|3.17|||||||||4|4|4|4||||||5|3|5|3|4|||||||4|4|4|4|3|4|1|3.43||||||||||4|4|4|4||||||2|4|3|||||1|1||||4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|8.1||1|1|1|1|M|Black||18|No||28206|One Parent: Female|$60,000 to $74,999||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||47|28205||Divorced|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502639463|31|0|1|502570705|1|0|1|500565299|2||-2||4|3|500004640, 500005291|500005291|-2||-2|0|10|||7464|9|||1|351297|-1|4|3|44
502760967|BBBS of Greater Charlotte|Main Office|C|Active|2011-12-08|NaT|Baseline|2011-10-14|2011-12-08|Complete|Done|1|2|4|1|3|3|2.33|||||||||4|4|4|4|3|4|3.83|||||||||4|2|2|2.67||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|||63.2||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|$25,000 to $29,999|Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||29|28120|Bachelors Degree|Single|Govt: Clerical||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502761879|31|0|2|502666332|31|0|2|500579826|2||-2||2|1||500005291|-2||-2|2203|12|||7464|9|||1|351583|-1|4|3|44
502212598|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-18|2013-08-15|Followup|2012-10-18|2012-12-07|Declined|Late||||||||4|1|3|3|2|4|2.83|||||||||2|4|4|1|2|3|2.67||||||3|4|4|3.67|||||||2|3|3|4|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Red|Amachi|Volunteer: Moved|21.9||2|2|1|1|F|Black||17|Yes|Mother|28215|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||28|28202|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|502213028|31|0|2|502715153|1|0|2|500558562|2||500003586||4|3|500000294|500000294|-2||-2|7016|11|||7464|9|||1|353512|151061|4|1|45
502698363|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-18|2013-12-06|Followup|2012-10-18|2013-01-02|Expired|Late||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4|4|1|3.5||||||4|4|4|4|||||||4|4|4|4|4||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||2|4|3||||2|2||||4|4||Red|Amachi|Volunteer: Lost contact with child/agency|25.6||1|1|1|1|M|Black||18|Yes|GrandMother|28203|Grandparents|Unknown||Yes||Self|General Community|Amachi|Enrollment|M|Black||43|28208|Bachelors Degree|Single|Education|28217|0|0|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500015820|502699208|31|0|1|502641410|31|0|1|500557390|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7452|6|||1|353665|341569|4|0|45
501023408|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-05|NaT|Followup|2012-11-05|2013-01-09|Complete|Late|4|1|4|2|3|3|2.83||||||||||||||||||||||||4|3|3|3.33||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||100.3||1|1|1|1|M|Hispanic|Other South American|17|No|Mother|28273|One Parent: Female|Less than $10,000||Yes||Self|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501023677|3|15|1|501356600|1|0|1|500296545|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|353690||4|3|45
500185734|BBBS of Greater Charlotte|Main Office|C|Completed|2003-10-15|2013-08-15|Followup|2012-10-15|2012-11-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|118||1|1|1|1|F|Black||21||Mother|28203|One Parent: Female|Unknown||No||Neighbor/Friend|General Community||Match Support|F|White||45|28202|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187476|31|0|2|500188688|1|0|2|500036688|2||-2||4|3|||-2||-2|0|8|||7464|9|||1|354320||4|1|45
500185723|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-05|2015-06-25|Followup|2012-09-05|2012-09-05|Complete|Done|3|2|3|3|3|3|2.83|||||||||2|3|3|3|3|3|2.83|||||||||4|3|3|3.33||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|81.6||2|2|1|1|M|Black||19||Mother|28214|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|M|Black||36|28214|Bachelors Degree|Single|Tech: Computer/Programmer|28147|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187335|31|0|1|501310677|31|0|1|500284133|2||-2||4|3|||-2||-2|6855|8|||7464|9|||1|354446||4|3|45
502699353|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-31|2014-01-30|Baseline|2011-10-20|2011-10-31|Complete|Done|3|3|4|2|4|4|3.33|||||||||3|3|3|4|4|3|3.33|||||||||3|3|3|3||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||1|1||||4|4||||Yellow|Project Big|Volunteer: Moved|27||2|2|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown||No||School|General Community|PERL 2014-2016, Project Big|Match Support|F|White||29|28204|Bachelors Degree|Single|Business|28255|0|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502700198|31|0|2|502530062|1|0|2|500568290|2||-2||4|2|500004640|500004640, 500014681|-2|500000294|-2|0|4|||7464|9|||1|355021|-1|4|3|44
502371558|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-31|NaT|Baseline|2011-10-20|2011-10-31|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|2|3|||||1|1||||4|4||||Green|||64.5||1|1|2|2|M|Black||17|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020752|502371997|31|0|1|502528355|1|0|1|500568298|2||-2||2|1||500000294, 500005291|-2||-2|0|10|||132|8|||1|355033|-1|4|3|44
502580335|BBBS of Greater Charlotte|Main Office|C|Active|2011-11-30|NaT|Baseline|2011-10-20|2011-11-30|Complete|Done|3|2|1|1|1|3|1.83|||||||||2|4|3|1|4|3|2.83|||||||||4|4|3|3.67||||||5|2|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|||63.5||1|1|1|1|F|Black||16||GrandMother|28269|Grandparents|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28269|Masters Degree|Single|Finance: Banking|28255|15|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502580838|31|0|2|502677590|31|0|2|500571804|2||-2||2|1||500005291|-2||-2|0|10|||7464|9|||1|355336|-1|4|3|44
502681369|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-26|2013-08-29|Baseline|2011-10-21|2011-10-26|Complete|Done|3|3|4|4|2|4|3.33|||||||||3|1|4|4|1|4|2.83|||||||||4|3|4|3.67||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|2|3.71||||||||||2|3|1|2||||||3|4|3.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Child: Lost interest|22.1||1|1|1|1|F|White||16|No|Mother|28262|One Parent: Female|$25,000 to $29,999||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||36|28205|Bachelors Degree|Single|Business: Human Resources|28202|4|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502682197|1|0|2|502726053|1|0|2|500568638|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|355566|-1|4|3|44
502613782|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-17|2013-09-12|Baseline|2011-10-21|2011-11-17|Complete|Done|1|4|1|2|1|1|1.67|||||||||4|4|4|3|4|4|3.83|||||||||4|2|2|2.67||||||5|5|5|5|5|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||2|1|1.5|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|21.8||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28202|Bachelors Degree|Single|Consultant||12|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500004169|502614394|31|0|1|502719849|1|0|1|500568690|2||-2||4|3||500005291|-2||-2|0|10|||46|2|||1|355624|-1|4|3|44
502604900|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-15|2015-05-14|Baseline|2011-10-24|2011-11-15|Complete|Done|3|1|1|1|1|1|1.33|||||||||1|1|2|1|1|3|1.5|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|41.9||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||30|28211|Bachelors Degree|Single|Finance: Accountant|28204|0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502605417|1|0|1|502582742|1|0|1|500577855|2||-2||4|1|||-2|500000294|-2|6854|8|||7464|9|||1|356462|-1|4|3|44
501101153|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-30|2013-08-30|Followup|2012-09-30|2012-10-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Severity of challenges|59||1|2|2|3|M|Black||19||Mother|28205|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||62|28214|Bachelors Degree|Married|Human Services: Non-Profit|28214|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501101427|31|0|1|500789916|1|0|1|500293277|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|357379||4|1|45
500970267|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-29|NaT|Followup|2012-09-29|2012-10-30|Complete|Done|3|3|3|3|3|4|3.17|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Green|Amachi||77.5||1|1|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||61|28204||Divorced|Self-Employed, Entrepreneur||0|0|Billboard|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|2|502084649|1|0|2|500468192|2||500003586||2|1|500000294|500000294|-2|500000294|-2|5635|9|||125|1|||1|357694|174196|4|3|45
500931662|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-07|NaT|Followup|2012-09-07|2012-10-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||114.3||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$60,000 to $74,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||58|28270|Bachelors Degree|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500931932|31|0|1|500894084|1|0|1|500193824|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|357720||4|1|45
502529397|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-11|NaT|Followup|2012-08-11|2012-08-09|Complete|Done|4|1|4|2|4|4|3.17|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||4|5|2|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Green|Project Big||67.2||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||48|28216|Bachelors Degree|Married|Finance: Banking|28255|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502529850|31|0|1|500188946|31|0|1|500548763|2||500004641||2|1|500004640||-2||-2|6854|8|||7464|9|||1|357817||4|3|45
502681369|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-26|2013-08-29|Followup|2012-10-26|2012-11-02|Complete|Done|4|2|2|2|3|3|2.67|3|3|4|4|2|4|3.33|-19.82|2|3|3|2|2|2|2.33|3|1|4|4|1|4|2.83|-17.67|3|3|3|3|4|3|4|3.67|-18.26|2|1|2|1|1.5|3|5|5|4|4.25|-64.71|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|4|4|2|3|1|2|100|4|4|4|3|4|3.5|14.29|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child: Lost interest|22.1||1|1|1|1|F|White||16|No|Mother|28262|One Parent: Female|$25,000 to $29,999||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||36|28205|Bachelors Degree|Single|Business: Human Resources|28202|4|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502682197|1|0|2|502726053|1|0|2|500568638|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|357888|355566|4|3|45
502555105|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2012-08-30|Baseline|2011-10-26|2011-11-11|Complete|Done|3|4|3|4|1|2|2.83|||||||||2|3|2|3|3|2|2.5|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|2|3|2.67||||||4|1|2.5|||||2|2||||4|4||||Yellow||Child/Family: Moved|9.6||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|$25,000 to $29,999||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28205|Bachelors Degree|Married|Self-Employed, Entrepreneur|28205|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|502555558|31|0|1|502598372|1|0|1|500570292|2||-2||4|2|||-2||-2|6854|8|||46|2|||1|357924|-1|4|3|44
502670071|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-26|2014-03-20|Followup|2012-10-26|2012-09-25|Complete|Early|4|1|4|1|4|4|3|4|4|4|1|4|4|3.5|-14.29|2|3|4|2|4|4|3.17|4|3|4|4|4|4|3.83|-17.23|4|4|4|4|4|4|4|4|0|1|1|4|2|2|5|5|5|5|5|-60|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|3|3|3|3|4|3|3.33|-9.91|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Yellow|Amachi, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|28.8||1|1|1|1|F|Black||16|Yes|Mother|28083|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|Black||36|28269|Masters Degree|Single|Human Services: Youth Worker|28027|2|2|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|502670906|31|0|2|502685522|31|0|2|500557057|2||500003586||4|2|500000294, 500005291|500005291|-2||-2|0|10|||9229|13|||1|358058|341113|4|3|45
501250109|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-11|2013-02-27|Followup|2012-09-11|2012-11-26|Expired|Late||||||||3|1|3|1|3|3|2.33|||||||||3|3|3|3|4|3|3.17||||||3|3|3|3|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Red||Volunteer: Lost contact with child/agency|41.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28227|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|501250385|31|0|1|501790515|31|0|1|500381167|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|358684|13945|4|0|45
500186428|BBBS of Greater Charlotte|Main Office|C|Completed|2005-10-03|2013-09-30|Followup|2012-10-03|2012-11-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|95.9||1|2|2|3|M|Black||21||Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||40|28211|Bachelors Degree|Single|Unknown||0|0|Brochure|Media|Big|General Community||Match Support|277|60|598|500000170|500004169|500187986|31|0|1|500189441|1|0|1|500044683|2||-2||4|1|||-2||-2|0|10|||127|1|||1|360045||4|1|45
500948385|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-28|2013-01-09|Followup|2012-08-28|2012-10-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|64.4||1|1|1|1|F|Black||17|No|Mother|28214|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Asian|Chinese|32|28216|||Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|500948655|31|0|2|500885771|4|16|2|500187434|2||-2||4|2|||-2||-2|34|2|||46|2|||1|360634||4|1|45
502510347|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-31|2016-08-30|Followup|2012-10-31|2012-10-23|Complete|Done|3|2|3|4|3|2|2.83|4|1|2|1|4|4|2.67|5.99|2|3|2|2|4|3|2.67|1|4|2|2|2|2|2.17|23.04|4|3|3|3.33|4|4|4|4|-16.75|4|3|2|3|3|3|4|2|4|3.25|-7.69|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|4|4|3|2|1|2|100|3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child: Graduated|58||1|1|1|1|F|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28262|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502510796|31|0|2|502677833|31|0|2|500557844|2||-2||4|1|500005291|500005291|-2||-2|0|5|||7464|9|||1|361626|310349|4|3|45
502699353|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-31|2014-01-30|Followup|2012-10-31|2013-01-12|Declined|Late||||||||3|3|4|2|4|4|3.33|||||||||3|3|3|4|4|3|3.33||||||3|3|3|3|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||3|3|3||||1|1||||4|4||Yellow|Project Big|Volunteer: Moved|27||2|2|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown||No||School|General Community|PERL 2014-2016, Project Big|Match Support|F|White||29|28204|Bachelors Degree|Single|Business|28255|0|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502700198|31|0|2|502530062|1|0|2|500568290|2||-2||4|2|500004640|500004640, 500014681|-2|500000294|-2|0|4|||7464|9|||1|361683|355021|4|1|45
502371558|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-31|NaT|Followup|2012-10-31|2012-12-26|Declined|Late||||||||3|2|3|3|3|3|2.83|||||||||3|4|4|3|2|4|3.33||||||4|4|4|4|||||||4|4|4|5|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|2|3||||1|1||||4|4||Green|||64.5||1|1|2|2|M|Black||17|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020752|502371997|31|0|1|502528355|1|0|1|500568298|2||-2||2|1||500000294, 500005291|-2||-2|0|10|||132|8|||1|361691|355033|4|1|45
501234606|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-16|NaT|Followup|2012-09-16|2012-12-01|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||101.9||1|1|1|1|F|Black||16|No|Mother|28216|Grandparents|Unknown||No|TV|Media|General Community||Match Support|F|Black||42|28212|Bachelors Degree|Single|Unknown|28202|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501234882|31|0|2|501233675|31|0|2|500287478|2||-2||2|1|||-2||-2|56|1|||7464|9|||1|361940||4|0|45
502370669|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-07|2012-11-29|Baseline|2011-11-01|2011-12-07|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||2|4|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Moved|11.8||2|2|1|1|M|Black||18|No|Mother|28269|One Parent: Female|$40,000 to $44,999|Y|Yes||Self|General Community||Match Support|M|Some Other Race||31|28205|Masters Degree|Single|Finance|28777|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500001281|502371107|31|0|1|502731507|41|0|1|500573204|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|362162|-1|4|3|44
500186765|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-05|2013-08-15|Followup|2012-09-05|2012-10-24|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|107.3||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||46|28078|Masters Degree|Widowed|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500004169|500188083|31|0|2|500189359|31|0|2|500037396|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|362503||4|1|45
500868942|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-20|NaT|Followup|2012-09-20|2012-11-05|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||113.8|Y|1|1|1|1|M|Black||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|M|White||54|28207||Married|Business: Sales||0|0|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500869211|31|0|1|500947018|1|0|1|500195082|2||-2||2|1|||-2||-2|0|10|||7458|9|||1|362504||4|1|45
502217445|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-14|2012-10-31|Baseline|2011-11-02|2011-11-11|Complete|Done|3|4|4|2|4|4|3.5|||||||||4|3|4|1|2|4|3|||||||||4|4|3|3.67||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|2|3.33||||||4|2|3|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|11.6||1|1|1|1|M|Black||19|No|Mother|28226|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||42|28277|Some College|Single|Self-Employed, Entrepreneur||5|0|Local Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500011746|502217876|31|0|1|502685222|31|0|1|500573483|2||-2||4|3|||-2||-2|0|10|||7437|1|||1|362521|-1|4|3|44
501938282|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-17|NaT|Followup|2012-11-17|2012-11-07|Complete|Done|4|2|2|1|2|2|2.17|||||||||1|1|1|1|2|1|1.17|||||||||2|2|2|2||||||1|1|2|2|1.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|1|2.5|||||2|2||||4|4||||Green|Amachi, Cabarrus County||75.9||1|1|1|1|F|White||14|Yes|Mother|28025|Two Parent|Unknown|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||63|28027|High School Graduate|Married|Self-Employed, Entrepreneur|28027|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501938680|1|0|2|502356100|1|0|2|500493871|2||500016307||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|362571||4|3|45
502753870|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2014-10-30|Baseline|2011-11-03|2011-11-30|Complete|Done|3|3|3|2|3|3|2.83|||||||||4|1|2|3|3|3|2.67|||||||||4|4|4|4||||||3||2|2||||||||4|4|4|4|4|4|4|4||||||||||3|2|3|2.67||||||3|4|3.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|35||2|2|1|1|F|Hispanic||16|No|Mother|28262|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|F|White||31|28210|Masters Degree|Single|Medical: Doctor, Provider||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502751081|3|0|2|502785389|1|0|2|500574313|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|363493|-1|4|3|44
501863951|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-18|2015-05-29|Followup|2011-12-18|2011-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Lost interest|65.3||1|1|2|2|F|Black||14|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28078|Bachelors Degree|Single|Business: Human Resources|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501864324|31|0|2|501601161|31|0|2|500421259|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|363835||4|1|45
502138562|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-14|2013-06-06|Followup|2012-12-14|2013-01-09|Complete|Done|4|1|1|2|3|3|2.33|2|3|4|3|1|1|2.33|0|2|3|3|3|2|3|2.67|1|2|1|4|4|4|2.67|0|4|4|4|4|3|3|3|3|33.33|5|5|5|5|5|5|4|4|5|4.5|11.11|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|2|3|33.33|2|2|2|2|0|4|4||||Green||Child: Lost interest|29.7||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||38|28216|Masters Degree|Single|Finance: Auditor|28217|3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500011746|502138991|31|0|1|502380370|31|0|1|500502780|2||-2||4|1|||-2||-2|0|10|||12183|14|||1|364555|220057|4|3|45
502255225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-08|2016-08-26|Followup|2012-11-08|2012-11-13|Complete|Done|4|3|4|2|3|3|3.17|2|2|2|4|1|4|2.5|26.8|2|3|3|2|2|3|2.5|2|3|3|2|2|3|2.5|0|4|4|4|4|4|3|3|3.33|20.12|4|4|3|4|3.75|5|3|5|3|4|-6.25|4|4|4|4|4|4|4|4|4|3|4|4|4|4|4|3.86|3.63|4|4|4|4|4|4|4|4|0|4|3|3.5|1|1|1|250|2|2|1|1|100|4|4||||Red||Volunteer: Moved|69.6||1|1|1|1|M|Hispanic||15||Mother|28212|One Parent: Female|Unknown||No|Spanish Radio|Media|General Community||Match Support|M|White||33|28226|Bachelors Degree|Single|Education: Teacher||3|0|Spanish Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502255655|3|0|1|502312682|1|0|1|500487118|2||-2||4|3|||-2||-2|7068|1|||11662|1|||1|364564|199091|4|3|45
500867579|BBBS of Greater Charlotte|Main Office|C|Completed|2007-09-22|2013-04-02|Followup|2012-09-22|2012-10-13|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|66.3||1|1|1|1|M|Black||23|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|No||Faith Organization|General Community|Amachi|Match Support|M|Black||42|28269||Single|Finance: Banking||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008629|500867843|31|0|1|500577903|31|0|1|500195387|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|9|||2238|7|||1|365852||4|1|45
501123191|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-20|2015-12-21|Followup|2012-10-20|2012-11-27|Complete|Done|3|1|4|1|4|4|2.83|||||||||2|4|4|3|1|4|3|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|4|3.67||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Moved|62||2|2|1|1|F|Black||15|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||48|28210|Some College|Single|Human Services||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500915629|31|0|2|502153920|1|0|2|500478644|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|366277||4|3|45
500829028|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-30|NaT|Followup|2012-11-30|2012-12-12|Complete|Done|1|4|2|2|3|3|2.5|||||||||2|4|4|2|4|3|3.17|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|4|3.33||||||2|4|3|||||2|2||||4|4||||Green|||75.5||3|3|2|2|F|Black||17|No|Mother|28209|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||39|28210|Masters Degree|Single|Education|28212|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502254499|31|0|2|501978180|1|0|2|500498594|2||-2||2|1|||-2|500000294, 500004640|-2|0|10|||7464|9|||1|366856||4|3|45
501288021|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-27|2016-02-01|Followup|2012-08-27|2012-08-08|Complete|Early|4|4|4|4|4|4|4|||||||||2|1|4|1|1|4|2.17|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||1|1|1|||||2|2||||4|4||||Green||Volunteer: Moved|89.2||1|1|1|1|F|Black||16|No|Mother|28211|Two Parent|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28027|PHD|Single|Education: College Professor|27411|1|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501288299|31|0|2|501249338|31|0|2|500281778|2||-2||4|1|||-2||-2|0|10|||46|2|||1|367514||4|3|45
502499851|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2015-07-07|Followup|2012-11-11|2012-11-27|Complete|Done|2|2|2|2|2|2|2|3|1|1|1|2|2|1.67|19.76|3|3|4|2|3|4|3.17|4|4|4|2|2|4|3.33|-4.8|4|4|4|4|4|4|4|4|0|2|4|4|4|3.5|5|5|5|4|4.75|-26.32|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|4|3|3.33|0|2|4|3|2|4|3|0|2|2|2|2|0|4|4|4|4|0|Red||Agency: Concern with Volunteer re: child safety|43.8||1|1|1|1|M|White||18|No|Mother|28210|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||39|28210|Masters Degree|Single|Finance|28106|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|502500300|1|0|1|502690262|1|0|1|500562789|2||-2||4|3|||-2||-2|0|10|||46|2|||1|367558|348364|4|3|45
501342393|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-22|2014-06-06|Followup|2012-10-22|2012-12-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|67.4||1|1|1|1|F|White||19|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Business: Sales||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501342672|1|0|2|501210017|1|0|2|500293459|2||-2||4|1|||-2||-2|0|10|||46|2|||1|367635||4|1|45
500713817|BBBS of Greater Charlotte|Main Office|C|Active|2009-10-30|NaT|Followup|2012-10-30|2012-12-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||88.5||2|2|1|1|M|Black||16||Mother|28216|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28078|||Medical: Pharmacist|28210|10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|500714084|31|0|1|501834795|1|0|1|500396466|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|367661||4|1|45
501614040|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-11|2013-02-28|Followup|2012-11-11|2013-01-26|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|39.6||1|1|1|1|M|Hispanic||16|No|Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||29|28273|||Facilities/Maintenance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|501614360|3|0|1|501864748|1|0|1|500404360|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|367700||4|0|45
502698998|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2014-03-13|Followup|2012-11-11|2012-10-31|Complete|Done|4|4|4|4|4|4|4|3|2|2|1|3|3|2.33|71.67|4|4|4|4|4|4|4|3|2|3|3|3|3|2.83|41.34|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3|4|4|4|3.75|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|3|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Yellow||Child/Family: Lost contact with volunteer/agency|28||1|1|1|1|F|Black||18|No|GrandMother|28211|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28203|Masters Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500012459|502699843|31|0|2|502692148|1|0|2|500564380|2||-2||4|2||500005291|-2||-2|0|4|||7464|9|||1|367756|350301|4|3|45
500867581|BBBS of Greater Charlotte|Main Office|C|Completed|2007-09-28|2014-02-06|Followup|2012-09-28|2012-10-09|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|76.3||1|1|2|2|M|Black||21|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999||No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||40|28269|Masters Degree|Single|Finance: Accountant|28255|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|500867843|31|0|1|500708515|1|0|1|500195388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|367807||4|3|45
502714405|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-08|2015-08-06|Baseline|2011-11-11|2011-12-08|Complete|Done|3|3|2|2|3|4|2.83|||||||||2|3|3|3|4|4|3.17|||||||||4|4|4|4||||||3|5|3|3|3.5|||||||4|3|4|4|4|4|4|3.86||||||||||3|4|4|3.67||||||1|1|1|||||1|1||||4|4||||Green||Child: Graduated|43.9||1|1|1|1|M|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||33|28213|Associate Degree|Single|Transport: Driver|28205|5|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500017732|502715293|31|0|1|502764673|31|0|1|500577475|2||-2||4|1||500005291|-2||-2|56|1|||7446|3|||1|367813|-1|4|3|44
502714414|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-08|2012-08-29|Baseline|2011-11-11|2011-12-08|Complete|Done|2|2|2|2|3|3|2.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|3|4|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|1|1.5|||||1|1||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|8.7||1|1|1|1|M|Black||18|No|Mother|28206|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||26|28213|Some College|Single|Business||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500001281|502715293|31|0|1|502769005|31|0|1|500577485|2||-2||4|1||500005291|-2||-2|56|1|||7462|13|1208|5|1|367824|-1|4|3|44
502604900|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-15|2015-05-14|Followup|2012-11-15|2012-11-29|Complete|Done|3|2|2|2|3|3|2.5|3|1|1|1|1|1|1.33|87.97|3|2|3|2|3|3|2.67|1|1|2|1|1|3|1.5|78|4|3|3|3.33|4|4|4|4|-16.75|4|3|3|4|3.5|4|4|3|3|3.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|2|3|33.33|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Lost contact with child/agency|41.9||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||30|28211|Bachelors Degree|Single|Finance: Accountant|28204|0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502605417|1|0|1|502582742|1|0|1|500577855|2||-2||4|1|||-2|500000294|-2|6854|8|||7464|9|||1|369047|356462|4|3|45
501129781|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-15|2015-01-15|Followup|2012-11-15|2012-12-19|Complete|Done|4|1|4|4|4|4|3.5|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Family structure changed|50||1|2|4|6|F|Black||17||Mother|28217|Two Parent|Unknown||No||School|General Community||Match Support|F|Black||48|28273|Bachelors Degree|Married|Business: Mgt, Admin|28273|4|0|Recruitment Event|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500018987|501130055|31|0|2|500189245|31|0|2|500494855|2||-2||4|1|||-2||-2|0|4|||7459|10|||1|369572||4|3|45
502613782|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-17|2013-09-12|Followup|2012-11-17|2013-02-01|Expired|Late||||||||1|4|1|2|1|1|1.67|||||||||4|4|4|3|4|4|3.83||||||4|2|2|2.67|||||||5|5|5|5|5||||||||||4|4|4|4|3|4|4|3.86||||||4|4|3|3.67|||||2|1|1.5||||2|2||||4|4||Red||Volunteer: Lost contact with child/agency|21.8||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28202|Bachelors Degree|Single|Consultant||12|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500004169|502614394|31|0|1|502719849|1|0|1|500568690|2||-2||4|3||500005291|-2||-2|0|10|||46|2|||1|370288|355624|4|0|45
502738004|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2012-03-23|Baseline|2011-11-17|2011-11-30|Complete|Done|3|3|3|2|2|3|2.67|||||||||3|3|3|3|4|3|3.17|||||||||3|2|2|2.33||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Infraction of match rules/agency policies|3.7||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28262|Two Parent: Not Married|Unknown|Y|No||Self|General Community||Match Support|F|Hispanic||36|28202||Single|Finance: Banking||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502738904|3|15|2|502620216|3|0|2|500579434|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|370646|-1|4|3|44
500185846|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-28|2014-10-23|Followup|2012-09-28|2012-09-18|Complete|Done|1|4|4|4|4|4|3.5|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|1|2.67||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|120.8||1|2|1|2|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||65|28256|Bachelors Degree||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187437|31|0|2|500188764|31|0|2|500038142|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|372105||4|3|45
500191820|BBBS of Greater Charlotte|Main Office|C|Completed|2005-09-30|2013-08-29|Followup|2012-09-30|2012-11-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|94.9|Y|2|2|2|2|M|Black||19||Mother|28227||Unknown||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||72|28214||Married|Retired||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500191823|31|0|1|500191501|31|0|1|500044434|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|8|||2238|7|||1|372106||4|1|45
500871683|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-01|2016-02-22|Followup|2012-10-01|2012-11-09|Complete|Done|1|1|2|1|4|4|2.17|||||||||4|4|4|2|2|4|3.33|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|100.7||1|1|1|1|M|Black||19|Yes|Aunt|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|M|White||46|28209|Masters Degree|Single|Self-Employed, Entrepreneur|28209|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500871952|31|0|1|500933829|1|0|1|500199601|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|372111||4|3|45
501340102|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-03|2013-04-25|Followup|2012-10-03|2012-10-04|Complete|Done|3|4|4|4|3|3|3.5|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||2|2||||4|4||||Red|Amachi|Child/Family: Time constraints|54.7||1|1|1|1|M|Multi-race (Black & Hispanic)||18|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||50|28269|Masters Degree|Married|Customer Service|28269|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340381|38|0|1|501316292|1|0|1|500287888|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|372112||4|3|45
501114443|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-08|2013-07-25|Followup|2012-10-08|2012-11-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|57.5||1|1|2|2|M|Black||22|No|Uncle|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||34|28205|Juris Doctorate (JD)|Married|Law: Lawyer||0|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501114708|31|0|1|501180846|1|0|1|500290376|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||46|2|||1|372114||4|1|45
501253195|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-24|NaT|Followup|2012-10-24|2012-10-19|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|3|4|2|1|4|3|||||||||4|4|4|4||||||5|3|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi||100.7||1|1|2|2|M|Black||15|Yes|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28203|Masters Degree|Single|Medical: Doctor, Provider|28211|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501253471|31|0|1|500395148|1|0|1|500282924|2||500003586||2|1|500000294||-2||-2|0|10|||7464|9|||1|372116||4|3|45
500185907|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2015-02-18|Followup|2012-10-29|2012-11-09|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|99.7||2|3|1|1|F|Black||19|Yes|Mother|28262|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||48|28212||Single|Medical: Healthcare Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187470|31|0|2|500697782|31|0|2|500134557|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|372117||4|3|45
501224287|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-30|2014-01-23|Followup|2012-10-30|2012-10-30|Complete|Done|4|3|4|2|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Child: Lost interest|62.8||1|1|1|1|M|Black||19|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||43|28262|Bachelors Degree|Married|Customer Service|28211|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501224558|31|0|1|501343190|31|0|1|500298289|2||-2||4|3|500000294|500000294|-2|500000294|-2|5635|9|||2230|7|||1|372118||4|3|45
501014187|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-07|NaT|Followup|2012-11-07|2012-11-12|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||100.2||2|2|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||48|28205|Bachelors Degree|Living w/ Significant Other|Human Services: Non-Profit|28205|3|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501404007|1|0|2|500306699|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7671|13|||1|372119||4|3|45
502380578|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-22|2014-05-15|Followup|2013-11-22|2013-11-20|Complete|Done|4|4|4|4|4|4|4|4|4|4|3|4|4|3.83|4.44|3|2|3|3|4|4|3.17|2|1|3|3|1|3|2.17|46.08|4|4|4|4|4|4|4|4|0|4|5|5|5|4.75|2|3|2|3|2.5|90|4|4|4|4|3|4|4|3.86|4|4|4|4|1|3|1|3|28.67|3|3|3|3|4|4|4|4|-25|3|3|3|3|4|3.5|-14.29|1|1|2|2|-50|4|4||||Yellow||Child/Family: Moved|29.7||2|2|3|3|F|Black||16||Mother|28213|Other/Unknown|Unknown||Yes||School|General Community||Match Support|F|Black||29|28262|Bachelors Degree|Single|Student: College||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|502381016|31|0|2|502138981|31|0|2|500579112|2||-2||4|2|||-2||-2|0|4|||7496|10|||1|372907|204339|4|3|45
502672482|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-18|2013-08-29|Followup|2012-10-18|2012-10-23|Complete|Done|3|2|2|1|3|4|2.5|||||||||4|3|2|3|3|4|3.17|||||||||4||3|||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Project Big|Volunteer: Lost contact with child/agency|22.4||1|1|1|1|M|Hispanic||14|No|Mother|28208|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Project Big|Match Support|M|White||27|28209|Bachelors Degree|Single|Tech: Support, Writing|29707|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502673310|3|0|1|502621665|1|0|1|500566301|2||500004641||4|3|500004640|500004640|-2||-2|0|10|||7464|9|||1|373723||4|3|45
502674024|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-07|2016-05-17|Baseline|2011-11-28|2011-12-07|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|4|4|4|4|3|3.5|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green||Child: Lost interest|53.3||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Sales||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018851|502674852|31|0|2|502660051|1|0|2|500581910|2||-2||4|1||500005291|-2||-2|0|10|||7496|10|||1|374331|-1|4|3|44
500826592|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-08|2016-10-18|Followup|2012-10-08|2012-11-12|Complete|Done|3|4|4|1|4|4|3.33|||||||||3|4|4|1|2|4|3|||||||||4|4|4|4||||||4|4|2|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|84.3||3|3|1|1|F|Black||20|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|F|White||33|28277|Bachelors Degree|Living w/ Significant Other|Unknown|28209|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|2|501314246|1|0|2|500382768|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|375016||4|3|45
500186190|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-13|2014-08-20|Followup|2012-10-13|2012-12-21|Complete|Late|4|4|4|4|4|4|4|||||||||4|4|4|1|2|4|3.17|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|118.2||1|1|2|2|F|Black||20||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187761|31|0|2|500189140|31|0|2|500037140|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|375018||4|3|45
502702145|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-21|2016-05-24|Baseline|2011-11-30|2011-12-21|Complete|Done|3|3|4|3|4|4|3.5|||||||||3|4|4|4|4|4|3.83|||||||||3|3|3|3||||||5|4|2|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|2|3|2.67||||||3|2|2.5|||||2|2||||4|4||||Red||Child: Graduated|53.1||1|1|2|2|F|Black||17|No|Mother|28083|One Parent: Female|$60,000 to $74,999||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020753|502702991|31|0|2|502204211|31|0|2|500582836|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|375724|-1|4|3|44
502753870|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2014-10-30|Followup|2012-11-30|2012-12-12|Complete|Done|4|4|4|4|3|4|3.83|3|3|3|2|3|3|2.83|35.34|4|4|4|4|4|4|4|4|1|2|3|3|3|2.67|49.81|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3||2|2|||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|2|3|2.67|49.81|4|4|4|3|4|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Time constraint|35||2|2|1|1|F|Hispanic||16|No|Mother|28262|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|F|White||31|28210|Masters Degree|Single|Medical: Doctor, Provider||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502751081|3|0|2|502785389|1|0|2|500574313|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|375730|363493|4|3|45
502838696|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2012-03-28|Baseline|2011-11-30|2011-11-30|Comprehension|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Feels incompatible with child/family|3.9||1|1|1|1|F|Hispanic||15|No|Mother|28031|Two Parent|Unknown||Yes||School|General Community||Match Support|F|White||51|28031|Some College|Married|Real Estate: Realtor|28031|5|0||Relative|Big|General Community||RTBM|277|60|598|500000170|500011746|502839988|3|0|2|502445477|1|0|2|500582889|2||-2||4|3|||-2||-2|0|4|||0|11|||1|375787|-1|4|2|44
502580335|BBBS of Greater Charlotte|Main Office|C|Active|2011-11-30|NaT|Followup|2012-11-30|2013-02-10|Declined|Late||||||||3|2|1|1|1|3|1.83|||||||||2|4|3|1|4|3|2.83||||||4|4|3|3.67|||||||5|2|4|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||3|2|2.5||||2|2||||4|4||Green|||63.5||1|1|1|1|F|Black||16||GrandMother|28269|Grandparents|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28269|Masters Degree|Single|Finance: Banking|28255|15|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502580838|31|0|2|502677590|31|0|2|500571804|2||-2||2|1||500005291|-2||-2|0|10|||7464|9|||1|375938|355336|4|1|45
502307545|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2013-08-29|Followup|2012-11-30|2012-11-21|Complete|Done|3|2|2|2|3|4|2.67|3|3|3|2|3|3|2.83|-5.65|2|4|3|3|3|3|3|2|3|3|3|3|3|2.83|6.01|4|3|3|3.33|3|3|3|3|11|3|2|3|3|2.75|3|3|3|4|3.25|-15.38|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|4|4|4|2|1|1.5|166.67|2|2|1|1|100|4|4||||Green|Project Big|Child/Family: Lost contact with volunteer/agency|21||2|2|1|1|F|Hispanic||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Hispanic||38|28209|Bachelors Degree||Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502307977|3|0|2|502782829|3|0|2|500582593|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7464|9|||1|375968|194334|4|3|45
502589869|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2015-10-29|Followup|2012-11-30|2012-12-19|Complete|Done|4|1|3|1|2|4|2.5|4|2|2|3|1|1|2.17|15.21|3|4|4|4|4|4|3.83|2|4|4|4|4|4|3.67|4.36|4|4|4|4|4|4|4|4|0|5|5|5|5|5|4|5|4|5|4.5|11.11|4|4|4|4|4|4|4|4|4|3|4|4|4|4|3|3.71|7.82|4|4|4|4|4|3|4|3.67|8.99|4|4|4|2|3|2.5|60|2|2|2|2|0|4|4|4|4|0|Green|Project Big|Child/Family: Lost contact with volunteer/agency|46.9||2|2|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28205|Bachelors Degree|Married|Business|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502590381|31|0|2|502701252|1|0|2|500582617|2||500004641||4|1|500004640|500004640, 500005291|-2|500000294|-2|0|4|459|3|7496|10|||1|375969|290937|4|3|45
501353940|BBBS of Greater Charlotte|Main Office|C|Active|2011-11-30|NaT|Followup|2012-11-30|2013-01-10|Complete|Done|4|3|3|2|3|4|3.17|||||||||2|2|3|2|3|3|2.5|||||||||4|3|3|3.33||||||3|3|2|2|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Green|Amachi||63.5||3|3|1|1|M|Black||16|No|Relative: Other|28205|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||33|28226|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|10|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500020752|501354219|31|0|1|502710990|1|0|1|500574615|2||500003586||2|1|500000294|500000294, 500005291|-2||-2|34|2|||17161|11|||1|376460||4|3|45
502745717|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-12|2013-02-28|Baseline|2011-12-01|2012-01-12|Complete|Done|3|1|4|1|4|4|2.83|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||3|4|3|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|2|3|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|13.6||1|1|1|1|F|Multi-race (Black & White)||17|No|Mother|28278|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|F|Asian||34|28278|Bachelors Degree|Single|Govt|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|502746625|36|0|2|502712044|4|0|2|500583497|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|376817|-1|4|3|44
502328599|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-10-31|Baseline|2011-12-01|2012-02-22|Complete|Done|4|1|4|1|4|3|2.83|||||||||2|4|4|2|2|4|3|||||||||2|2|2|2||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Red||Volunteer: Time constraint|32.3||1|1|1|1|M|Black||15|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||73|28226|Bachelors Degree|Widowed|Construction||7|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502329034|31|0|1|502732347|1|0|1|500594124|2||-2||4|3|||-2||-2|0|10|||131|1|||1|376848|-1|4|3|44
502260656|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-18|2013-03-19|Followup|2012-10-18|2012-10-22|Complete|Done|3|2|2|1|4|4|2.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Moved|29||2|2|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28078|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||33|28078|Associate Degree|Married|Education: Teacher Asst/Aid||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502261088|38|0|2|502249984|1|0|2|500475564|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|377216|170947|4|3|45
502247579|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-02|2016-05-10|Followup|2012-12-02|2012-12-14|Complete|Done|4|3|3|1|4|4|3.17|4|3|3|2|3|4|3.17|0|3|4|4|2|2|4|3.17|2|3|2|2|2|3|2.33|36.05|4|4|4|4|4|4|4|4|0|5|3|4|3|3.75|3|3|3|3|3|25|4|3|4|4|2|3|3|3.29|4|4|4|4|4|4|4|4|-17.75|4|4|3|3.67|4|4|4|4|-8.25|2|2|2|3|3|3|-33.33|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|53.3||2|2|1|1|F|Black||15|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||47|28226|Bachelors Degree|Single|Education: Teacher||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500017732|502248010|31|0|2|502681447|31|0|2|500575685|2||500003586||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|10|||2238|7|||1|377223|194970|4|3|45
500958307|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-19|NaT|Followup|2012-09-19|2012-08-29|Complete|Early|3|4|4|4|4|4|3.83|||||||||2|3|2|1|2|2|2|||||||||4|4|4|4||||||3|2|2|2|2.25|||||||4|4|4|4|4|3|2|3.57||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi, Cabarrus County||113.9|Y|1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$40,000 to $44,999|Y|No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|Black||62|28213||Married|Finance: Economist||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500958577|31|0|1|500876132|31|0|1|500193868|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|377685||4|3|45
502708670|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-23|2014-02-06|Baseline|2011-12-05|2011-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|25.5||1|1|1|1|F|Black||18|No|Mother|28209|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||28|28215|Bachelors Degree|Single|Customer Service|28078|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500015820|502709557|31|0|2|502756331|1|0|2|500584031|2||-2||4|3|||-2||-2|0|4|||7462|13|||1|377810|-1|4|1|44
502256918|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-07|2013-04-25|Followup|2012-12-07|2013-01-09|Declined|Done||||||||4|4|4|1|3|4|3.33|||||||||3|3|4|2|4|3|3.17||||||4|4|4|4|||||||3|3|2|5|3.25||||||||||4|4|4|4|4|4|4|4||||||4|3|4|3.67|||||3|3|3||||2|2|||||||Red||Child/Family: Moved|28.6||1|1|1|1|M|Hispanic||16|No|Mother|28212|One Parent: Female|Unknown||No|Spanish Print|Media|General Community||Match Support|M|White||38|28209|Juris Doctorate (JD)|Single|Law||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502257350|3|0|1|502143354|1|0|1|500501039|2||-2||4|3|||-2||-2|7063|1|||7464|9|||1|378147|217658|4|1|45
500186646|BBBS of Greater Charlotte|Main Office|C|Completed|2005-10-20|2013-09-23|Followup|2012-10-20|2013-01-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|95.1||3|3|3|3|F|Some Other Race||21||Mother|28217|Other/Unknown|Unknown||No||Neighbor/Friend|General Community||Match Support|F|Black||39|28216|Some College||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500188044|41|0|2|500189263|31|0|2|500047741|2||-2||4|2|||-2||-2|0|8|||7464|9|||1|378403||4|0|45
501725162|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2016-10-14|Followup|2012-10-29|2012-10-29|Complete|Done|3|1|3|2|4|3|2.67|4|1|2|1|4|4|2.67|0|2|4|3|3|3|3|3|3|4|2|3|3|3|3|0|4|4|4|4|1|4|4|3|33.33|4|5|4|4|4.25|5|1|5|5|4|6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|2|3.33|20.12|4|4|4|4|3|3.5|14.29|2|2|2|2|0|4|4||||Green||Agency: Challenges with program/partnership|83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501724831|39|0|1|501833178|1|0|1|500394157|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|378556|16143|4|3|45
501729405|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-14|2013-06-16|Followup|2012-12-14|2013-01-25|Complete|Done|4|4|4|4|3|4|3.83|||||||||3|4|3|4|3|3|3.33|||||||||4|3|3|3.33||||||2|4|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|30.1||2|2|1|1|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|RTBM|F|White||33|28204|Bachelors Degree|Single|Business: Sales|28210|0|7|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501729745|31|0|2|502361956|1|0|2|500501689|2||500004772||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|4|||7464|9|||1|378909||4|3|45
502419933|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-07|2014-09-04|Followup|2012-12-07|2012-11-28|Complete|Done|2|2|3|3|2|2|2.33|3|2|3|3|3|3|2.83|-17.67|3|2|3|1|3|3|2.5|3|3|3|2|3|4|3|-16.67|3|4|3|3.33|4|4|4|4|-16.75|3|3|2|3|2.75|4|4|4|4|4|-31.25|4|4|4|4|4|4|3|3.86||4|4|4|4|4|4|||4|4|4|4|4|4|4|4|0|4|1|2.5|4|4|4|-37.5|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Time constraint|32.9||2|2|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$40,000 to $44,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||58|28031|Bachelors Degree|Living w/ Significant Other|Business: Mgt, Admin||22|0|Big Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500011349|502371107|31|0|1|502669194|1|0|1|500571419|2||-2||4|2||500005291|-2||-2|0|10|||7456|8|||1|379031|254462|4|3|45
500186192|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2014-10-13|Followup|2012-11-18|2012-11-30|Complete|Done|3|3|3|4|3|3|3.17|||||||||2|3|2|2|2|3|2.33|||||||||4|4|4|4||||||4|3|2|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|46.8||2|2|1|1|F|Black||20||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|Black||33|28208||Single|Service: Restaurant||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187762|31|0|2|502323059|31|0|2|500490136|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|379103||4|3|45
502674024|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-07|2016-05-17|Followup|2012-12-07|2012-11-28|Complete|Done|1|4|4|1|4|4|3|4|4|4|3|4|4|3.83|-21.67|4|4|4|4|4|4|4|2|4|4|4|4|3|3.5|14.29|4|4|4|4|4|4|4|4|0|4|5|2|5|4|4|4|4|3|3.75|6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|3|4|3|3.33|20.12|3|2|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Green||Child: Lost interest|53.3||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Sales||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018851|502674852|31|0|2|502660051|1|0|2|500581910|2||-2||4|1||500005291|-2||-2|0|10|||7496|10|||1|379188|374331|4|3|45
502760967|BBBS of Greater Charlotte|Main Office|C|Active|2011-12-08|NaT|Followup|2012-12-08|2012-12-14|Complete|Done|1|1|4|2|1|3|2|1|2|4|1|3|3|2.33|-14.16|4|4|4|4|4|4|4|4|4|4|4|3|4|3.83|4.44|4|4|4|4|4|2|2|2.67|49.81|4|5|5|5|4.75|5|5|5|5|5|-5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Green|||63.2||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|$25,000 to $29,999|Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||29|28120|Bachelors Degree|Single|Govt: Clerical||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502761879|31|0|2|502666332|31|0|2|500579826|2||-2||2|1||500005291|-2||-2|2203|12|||7464|9|||1|379553|351583|4|3|45
502714405|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-08|2015-08-06|Followup|2012-12-08|2013-02-22|Expired|Late||||||||3|3|2|2|3|4|2.83|||||||||2|3|3|3|4|4|3.17||||||4|4|4|4|||||||3|5|3|3|3.5||||||||||4|3|4|4|4|4|4|3.86||||||3|4|4|3.67|||||1|1|1||||1|1||||4|4||Green||Child: Graduated|43.9||1|1|1|1|M|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||33|28213|Associate Degree|Single|Transport: Driver|28205|5|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500017732|502715293|31|0|1|502764673|31|0|1|500577475|2||-2||4|1||500005291|-2||-2|56|1|||7446|3|||1|379583|367813|4|0|45
502805818|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-14|2013-12-19|Baseline|2011-12-09|2011-12-14|Complete|Done|3|1|4|1|3|3|2.5|||||||||2|3|3|2|2|4|2.67|||||||||4|3|3|3.33||||||3|2|4|4|3.25|||||||4|4|4|3|4|3|3|3.57||||||||||4|4|3|3.67||||||1|3|2|||||2|2||||4|4||||Green|Amachi|Child/Family: Moved|24.2||1|1|1|1|F|Black||18|Yes|GrandMother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||45|28213|Some College|Single|Business: Mgt, Admin|28202|1|3|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500015820|502807093|31|0|2|502704456|31|0|2|500585665|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|380178|-1|4|3|44
501142903|BBBS of Greater Charlotte|Main Office|C|Active|2008-06-05|NaT|Followup|2012-06-05|2012-06-08|Complete|Done|3|2|4|4|3|4|3.33|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||105.3||1|1|1|1|M|Black||14|Yes|GrandMother|28208|One Parent: Female|Less than $10,000||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|M|White||53|28204|Juris Doctorate (JD)|Married|Law: Lawyer|28244|16|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501143177|31|0|1|501236825|1|0|1|500268808|2||500003586||2|1|500000294|500000294|-2|500000294|-2|7294|13|||2238|7|||1|380590||4|3|45
501721579|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-24|2016-06-17|Followup|2012-07-24|2012-08-15|Complete|Done|1|1|4|1|1|4|2|||||||||2|1|4|1|2|3|2.17|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Moved|82.8||2|2|1|1|F|Multi-Race (None of the above)||14|No|Mother|28211|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||50|28227|Some College|Single|Human Services: Social Worker||2|5|St. Paul Baptist|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501721919|7|0|2|501687513|31|0|2|500375006|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||9609|7|||1|380674||4|3|45
502758832|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-17|2014-10-23|Baseline|2011-12-12|2011-12-17|Complete|Done|4|4|4|4|3|3|3.67|||||||||1|3|3|2|1|3|2.17|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Family structure changed|34.2||1|1|1|1|F|White||14|No|Mother|28027|One Parent: Female|$50,000 to $59,999||No||Relative|General Community||Match Support|F|White||33|28027|Masters Degree|Single|Education: Teacher|28027|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502759744|1|0|2|502666962|1|0|2|500586238|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|381135|-1|4|3|44
502310004|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-26|2014-05-01|Followup|2012-10-26|2012-12-26|Declined|Late||||||||4|4|4|4|3|3|3.67|||||||||2|3|4|4|3|4|3.33||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Yellow|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|42.2||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||No||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Enrollment|F|White||37|28078||Single|Business||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502310436|31|0|2|502331000|1|0|2|500483762|2||500003586||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7496|10|||1|381605|194875|4|1|45
501686310|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-30|2013-03-13|Followup|2012-10-30|2013-01-14|Expired|Late||||||||3|4|4|4|3|4|3.67|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||4|5|5|5|4.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|4|4||||1|1|||||||Red||Child/Family: Lost contact with volunteer/agency|40.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28211|One Parent: Female|Unknown||No|Radio|Media|General Community||Match Support|M|Black||34|28202|Juris Doctorate (JD)|Single|Law: Lawyer||1|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501686648|36|0|1|501818631|31|0|1|500392214|2||-2||4|3|||-2||-2|55|1|||7446|3|||1|381633|14832|4|0|45
502571727|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-13|2017-03-09|Baseline|2011-12-14|2012-01-13|Complete|Done|3|4|4|3|1|4|3.17|||||||||2|4|2|3|4|3|3|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|2|3.33||||||3|4|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|61.8||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|M|Black||45|28207|Masters Degree|Married|Tech: Management|28081|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|502572181|31|0|1|502769619|31|0|1|500586830|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|382185|-1|4|3|44
502805818|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-14|2013-12-19|Followup|2012-12-14|2013-02-10|Declined|Late||||||||3|1|4|1|3|3|2.5|||||||||2|3|3|2|2|4|2.67||||||4|3|3|3.33|||||||3|2|4|4|3.25||||||||||4|4|4|3|4|3|3|3.57||||||4|4|3|3.67|||||1|3|2||||2|2||||4|4||Green|Amachi|Child/Family: Moved|24.2||1|1|1|1|F|Black||18|Yes|GrandMother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||45|28213|Some College|Single|Business: Mgt, Admin|28202|1|3|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500015820|502807093|31|0|2|502704456|31|0|2|500585665|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|382225|380178|4|1|45
502280284|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-13|2013-07-31|Followup|2012-12-13|2013-01-25|Complete|Done|3|3|4|4|4|4|3.67|4|3|3|2|4|4|3.33|10.21|2|4|4|2|4|4|3.33|3|4|4|2|3|4|3.33|0|3|3|3|3|4|4|4|4|-25|4|3|3|3|3.25|3|3|3|3|3|8.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|2|2.5|3|3|3|-16.67|2|2|1|1|100|4|4||||Red|Project Big|Volunteer: Lost contact with child/agency|31.6||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|White||31|28205|Associate Degree|Married|Business: Human Resources||3|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502280719|31|0|2|502241391|1|0|2|500500329|2||500004641||4|3|500004640|500004640|-2|500004640|-2|0|10|||46|2|||1|382313|216597|4|3|45
502763567|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-30|2012-10-17|Baseline|2011-12-15|2011-12-30|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|3|3|2|2|3|2.67|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||2|4|3|||||2|2||||4|4||||Red|Project Big|Child/Family: Lost contact with volunteer/agency|9.6||1|1|2|2|F|Black||15|No|Mother|28211|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||34|28215|Some College|Single|Finance: Banking|28270|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|502764479|31|0|2|502672644|31|0|2|500587190|2||-2||4|3|500004640||-2||-2|0|4|||7464|9|||1|382782|-1|4|3|44
500936718|BBBS of Greater Charlotte|Main Office|C|Completed|2007-12-20|2016-06-16|Followup|2012-12-20|2012-11-27|Complete|Early|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||2|3|3|2.67||||||1|4|2.5|||||2|2||||4|4||||Green||Agency: Challenges with program/partnership|101.9||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28210|Bachelors Degree|Married|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500017732|500915629|31|0|1|501027885|1|0|1|500224574|2||-2||4|1|||-2|500014505, 500015184|-1|34|2|||46|2|||1|382858||4|3|45
500185637|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-29|2014-12-11|Followup|2012-12-29|2013-02-28|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|107.4||1|1|2|2|M|Black||20||Mother|28206|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Black||55|28297|Masters Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500187271|31|0|1|500189284|31|0|1|500073080|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|382867||4|1|45
500801567|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-26|2013-12-12|Followup|2012-10-26|2012-11-12|Complete|Done|2|4|4|4|3|3|3.33|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|4|5|3|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|49.5||2|2|1|1|M|Black||20||Mother|28213|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||62|28078|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500801835|31|0|1|501834907|1|0|1|500391790|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|382948||4|3|45
502787524|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-25|2014-08-29|Baseline|2011-12-15|2012-01-25|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|4|4|4|3.5|||||||||4|3|3|3.33||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4||||||||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|31.1||1|1|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28205|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Asian||29|28202||Single|Tech: Computer/Programmer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502788707|38|0|2|502272989|4|0|2|500587325|2||-2||4|3|||-2|500004640|-2|0|10|||7496|10|||1|382987|-1|4|3|44
502273093|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-01|2015-03-31|Followup|2012-10-01|2012-11-19|Complete|Late|3|3|3|2|3|3|2.83|||||||||3|3|3|2|3|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|4|3.33||||||3|3|3|||||2|2||||4|4||||Green||Child/Family: Moved|53.9||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||37|28277|PHD|Single|Medical: Healthcare Worker||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502273525|31|0|2|502252422|31|0|2|500471568|2||-2||4|1|||-2|500000294|-2|0|4|||7496|10|||1|383284||4|3|45
502317500|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-08|2015-07-31|Baseline|2011-12-16|2012-02-08|Complete|Done|4|2|1|2|4|4|2.83|||||||||2|3|4|2|2|4|2.83|||||||||4|4|4|4||||||4|3|2|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|2|2.5|||||2|2||||4|4||||Red|Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|41.7||1|1|2|2|M|Black||15|No|Mother|28214|One Parent: Female|Unknown||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|M|White||33|28214|Associate Degree|Single|Law: Security Officer|28208|2|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502317931|31|0|1|502658498|1|0|1|500587614|2||-2||4|3|500004640, 500004901|500004640, 500004901|-2||-2|0|4|||7464|9|||1|383492|-1|4|3|44
502758832|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-17|2014-10-23|Followup|2012-12-17|2012-12-12|Complete|Done|4|2|4|1|4|4|3.17|4|4|4|4|3|3|3.67|-13.62|2|4|4|2|2|3|2.83|1|3|3|2|1|3|2.17|30.41|4|4|4|4|4|4|4|4|0|5|5|5|5|5|4|5|4|5|4.5|11.11|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|4|3|3.33|0|4|4|4|3|4|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Green||Child: Family structure changed|34.2||1|1|1|1|F|White||14|No|Mother|28027|One Parent: Female|$50,000 to $59,999||No||Relative|General Community||Match Support|F|White||33|28027|Masters Degree|Single|Education: Teacher|28027|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502759744|1|0|2|502666962|1|0|2|500586238|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|383687|381135|4|3|45
502861536|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-08|2012-11-16|Baseline|2011-12-19|2012-02-08|Complete|Done|3|3|4|3|3|4|3.33|||||||||2|4|4|3|4|4|3.5|||||||||4|3|3|3.33||||||5|5|3|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child/Family: Infraction of match rules/agency policies|9.3||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||31|28213|Bachelors Degree|Single|Insurance|28262|3|0|BBBS National Site|Web Link|Big|General Community||RTBM|277|60|598|500000170|500011349|502862935|31|0|2|502876160|31|0|2|500595490|2||-2||4|3|||-2||-2|0|4|||46|2|||1|383944|-1|4|3|44
502570185|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2014-05-15|Followup|2012-06-30|2012-07-05|Complete|Done|3|1|4|3|3|4|3|||||||||3|4|3|3|3|4|3.33|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|34.5||1|1|1|1|F|Black||14|No|Mother|28206|Other/Unknown|Unknown||Yes||Relative|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||58|28226|Masters Degree|Single|Tech: Management|28078|0|2|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500017777|502570639|31|0|2|502191626|31|0|2|500542078|2||500004641||4|2|500000294, 500004640, 500004901, 500005291|500004640, 500005291|-2|500004640|-2|0|3|459|3|46|2|||1|384438||4|3|45
501853848|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-30|2014-08-29|Followup|2012-11-30|2012-12-23|Complete|Done|4|3|3|2|4|4|3.33|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|56.9||1|1|1|1|M|Black||15|Yes|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|M|Black||33|28273|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501854219|31|0|1|501839466|31|0|1|500405366|2||-2||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|384779||4|3|45
502732602|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-25|2013-06-18|Baseline|2011-12-21|2012-01-25|Complete|Done|4|2|4|1|1|4|2.67|||||||||2|2|3|4|3|4|3|||||||||4|4|4|4||||||3|3|5|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Yellow||Volunteer: Moved|16.8||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|White||29|28203|Masters Degree|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502733499|31|0|2|502766077|1|0|2|500588408|2||-2||4|2||500005291|-2||-2|0|5|||7464|9|||1|385114|-1|4|3|44
502702145|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-21|2016-05-24|Followup|2012-12-21|2012-12-12|Complete|Done|4|4|4|3|4|4|3.83|3|3|4|3|4|4|3.5|9.43|1|4|4|4|4|4|3.5|3|4|4|4|4|4|3.83|-8.62|4|4|4|4|3|3|3|3|33.33|5|5|5|5|5|5|4|2|4|3.75|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|3|3|3|2|3|2.67|12.36|4|4|4|3|2|2.5|60|2|2|2|2|0|4|4|4|4|0|Red||Child: Graduated|53.1||1|1|2|2|F|Black||17|No|Mother|28083|One Parent: Female|$60,000 to $74,999||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020753|502702991|31|0|2|502204211|31|0|2|500582836|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|385210|375724|4|3|45
500186133|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-14|2016-06-28|Followup|2012-10-14|2012-11-13|Complete|Done|3|2|3|2|3|3|2.67|||||||||3|3|3|3|4|3|3.17|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|140.5||1|1|1|1|M|White||18||Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||51|28262|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500187724|1|0|1|500188930|1|0|1|500036930|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|385337||4|3|45
500545326|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2016-09-02|Followup|2012-10-29|2012-10-19|Complete|Done|4|1|1|1|1|4|2|||||||||1|1|4|1|1|4|2|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|118.1|Y|1|1|1|1|M|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|Black||55|28214||Married|Clergy||12|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|1|500697845|31|0|1|500134545|2||-2||4|3|||-2||-2|0|10|||2238|7|||1|385625||4|3|45
502861544|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-03|2012-11-16|Baseline|2011-12-22|2012-01-03|Complete|Done|3|4|4|3|3|4|3.5|||||||||2|2|4|3|1|3|2.5|||||||||4|2|2|2.67||||||4|1|3|3|2.75|||||||2|2|2|4|4|3|3|2.86||||||||||3|4|2|3||||||1|1|1|||||2|2||||4|4||||Red||Child/Family: Infraction of match rules/agency policies|10.4||1|1|1|1|M|Black||20|No|Mother|28205|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Black||45|28210|Some College|Married|Tech: Production Line||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011349|502862935|31|0|1|502817316|31|0|1|500588737|2||-2||4|3|||-2||-2|0|4|||7496|10|||1|385730|-1|4|3|44
501744683|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-06|2012-11-28|Followup|2012-11-06|2012-10-20|Declined|Early||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|36.7||1|1|1|1|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||56|28270|Some College|Separated|Unknown|28277|7|7|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500013781|501745023|31|0|1|501863268|31|0|1|500405317|2||-2||4|1|||-2||-2|0|10|||46|2|||1|385737||4|1|45
501863951|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-18|2015-05-29|Followup|2012-12-18|2013-01-16|Complete|Done|3|2|4|2|4|4|3.17|||||||||4|3|3|3|4|4|3.5|||||||||3|3|3|3||||||4|3|3|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Child: Lost interest|65.3||1|1|2|2|F|Black||14|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28078|Bachelors Degree|Single|Business: Human Resources|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501864324|31|0|2|501601161|31|0|2|500421259|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|386093||4|3|45
501313839|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-11|2013-06-18|Followup|2012-11-11|2013-01-26|Expired|Late||||||||3|2|3|3|4|4|3.17|||||||||2|3|4|4|2|4|3.17||||||3|4|4|3.67|||||||4|5|5|5|4.75||||||||||4|4|4|3|2|2|1|2.86||||||3|4|3|3.33|||||3|3|3||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|43.2||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||36|28204|Bachelors Degree|Single|Consultant||4|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501314117|31|0|1|501788563|1|0|1|500396680|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|386101|590|4|0|45
502708670|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-23|2014-02-06|Followup|2012-12-23|2012-12-31|Complete|Done|4|2|4|1|4|4|3.17|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|2|3.33||||||2|3|2.5|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|25.5||1|1|1|1|F|Black||18|No|Mother|28209|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||28|28215|Bachelors Degree|Single|Customer Service|28078|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500015820|502709557|31|0|2|502756331|1|0|2|500584031|2||-2||4|3|||-2||-2|0|4|||7462|13|||1|386128|377810|4|3|45
500252077|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-24|2016-01-20|Followup|2012-11-24|2012-11-21|Complete|Done|4|1|2|2|3|4|2.67|||||||||2|3|3|1|1|3|2.17|||||||||4|3|3|3.33||||||3|3|4|5|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|85.8||3|3|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Tech: Computer/Programmer||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501750989|31|0|1|501365749|1|0|1|500317108|2||500003586||4|3|500000294|500000294|-2||-2|7295|11|||46|2|||1|386167||4|3|45
500186742|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-08|2016-06-30|Followup|2012-12-08|2012-12-12|Complete|Done|1|4|4|4|4|4|3.5|||||||||4|3|1|4|3|3|3|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|2|2|||||1|1||||4|4||||Green|Amachi|Child: Graduated|66.7||4|4|1|1|M|Black||19|Yes|Mother|28227|One Parent: Female|Unknown|Y|No||School|General Community|Amachi|Match Support|M|Black||52|28227|Masters Degree|Married|Education: Teacher|28227|2|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|502397541|31|0|1|500501282|2||500003586||4|1|500000294|500000294|-2|500000294, 500004640|-2|0|4|||12183|14|635|1|1|386169||4|3|45
501292079|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-11|2013-07-18|Followup|2012-12-11|2013-01-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Lost interest|55.2||1|1|1|1|F|Black||17|Yes|GrandMother|28214|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||31|28203|Bachelors Degree|Single|Consultant|28204|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501292357|31|0|2|501519897|1|0|2|500323243|2||500003586||4|1|500000294|500000294|-2||-2|7294|13|||7464|9|||1|386170||4|1|45
502180724|BBBS of Greater Charlotte|Main Office|C|Active|2010-12-30|NaT|Followup|2012-12-30|2012-12-14|Complete|Early|4|4|4|4|4|4|4|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||74.5|Y|2|2|2|2|M|Black||15|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502181148|31|0|1|502391505|31|0|2|500505039|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7438|1|||1|386562||4|3|45
501967613|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2013-02-26|Followup|2012-12-31|2013-01-24|Declined|Done||||||||4|3|3|3|3|4|3.33|||||||||3|4|3|3|3|2|3||||||4|3|3|3.33|||||||3|4|4|3|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Yellow||Volunteer: Time constraint|25.9||1|1|1|1|F|Black||20|No|Mother|28273|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Finance: Accountant|28277|3|5|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500012459|501968011|31|0|2|502311344|1|0|2|500498762|2||-2||4|2|||-2|500000294, 500004640|-2|34|2|||7496|10|||1|386748|148519|4|1|45
500733695|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-26|2015-03-03|Followup|2012-12-26|2012-12-22|Complete|Done|3|4|4|2|4|4|3.5|||||||||4|4|3|4|2|4|3.5|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.2||1|1|1|1|F|Black||19|Yes|GrandMother|28217|Grandparents|Less than $10,000|Y|No|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||34|28210|Bachelors Degree|Married|Finance: Accountant|28202|0|2|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500733962|31|0|2|500307108|1|0|2|500150172|2||500003586||4|3|500000294|500000294|-2||-2|7294|13|||2238|7|||1|386975||4|3|45
501340105|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2013-06-27|Followup|2012-12-12|2012-12-31|Complete|Done|1|2|1|2|3|3|2|||||||||3|3|4|2|3|4|3.17|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|4|3.33||||||3|2|2.5|||||1|1||||4|4||||Red|Amachi|Child: Graduated|54.5||1|1|1|1|F|Multi-race (Black & Hispanic)||21|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||53|28269||Married|Medical: Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340376|38|0|2|501514453|1|0|2|500322778|2||-2||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|387197||4|3|45
501114434|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-23|2014-06-12|Followup|2012-12-23|2013-01-21|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|65.6||1|1|1|1|M|Black||20|No|Uncle|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||33|28207|Masters Degree|Single|Finance: Accountant|28244|0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501114708|31|0|1|501315131|1|0|1|500324423|2||-2||4|3|500000294|500000294|-2||-2|0|10|||130|1|11|3|1|387234||4|3|45
501296349|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-01|2014-02-27|Followup|2012-12-01|2013-02-01|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|62.9||1|1|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||42|28214|Bachelors Degree|Single|Business: Mgt, Admin|28205|3|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501296627|31|0|2|501471640|31|0|2|500318555|2||||4|2|||-2|500000294|-2|0|4|||7464|9|||1|387263||4|1|45
502236953|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-17|2015-01-30|Followup|2012-08-17|2012-08-14|Complete|Done|3|1|2|4|4|3|2.83|||||||||2|3|3|1|2|4|2.5|||||||||4|4|4|4||||||3|4|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Red||Volunteer: Time constraint|53.5||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||50|28212|Some College|Married|Law: Police Officer||2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502237384|31|0|1|502232559|31|0|1|500464143|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|387706||4|3|45
500998933|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-19|2013-12-06|Followup|2012-11-19|2013-01-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|36.6||1|1|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|F|White||37|28210|Masters Degree|Single|Medical|28210|1|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500015820|500999202|31|0|2|502274159|1|0|2|500497430|2||500003586||4|3|500000294|500000294|-2|500000294, 500004640|-2|0|10|||7496|10|||1|388067||4|1|45
502290880|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-20|2014-03-31|Followup|2013-10-20|2013-11-18|Complete|Done|4|3|4|2|4|4|3.5|4|3|3|1|4|4|3.17|10.41|2|3|3|2|3|3|2.67|3|4|4|3|3|4|3.5|-23.71|4|3|3|3.33|4|4|4|4|-16.75|3|3|3|2|2.75|5|4|5|4|4.5|-38.89|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|4|4|4|4|4|4|0|2|4|3|2|4|3|0|2|2|2|2|0|4|4||||Green|Project Big|Child/Family: Time constraints|41.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|M|White||35|28202|Bachelors Degree|Single|Real Estate: Realtor|28208|2|10|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502291312|31|0|1|502261364|1|0|1|500471473|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7496|10|||1|388188|179708|4|3|45
502725760|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2014-09-24|Baseline|2012-01-04|2012-01-23|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|32||1|1|1|1|M|Black||16|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|Amachi|Match Support|M|Black||28|28226|Bachelors Degree|Single|Business: Sales|28217|0|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502726656|31|0|1|502687867|31|0|1|500589763|2||-2||4|2|500000294|500000294|-2||-2|0|10|||4748|14|633|1|1|388386|-1|4|3|44
502825916|BBBS of Greater Charlotte|Main Office|C|Active|2012-01-23|NaT|Baseline|2012-01-04|2012-01-23|Complete|Done|4|2|1|2|2|4|2.5|||||||||2|3|4|3|4|3|3.17|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Yellow|Amachi||61.7||1|1|2|2|F|Black||14|Yes|Mother|28273|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28208|Some College|Single|Education: Teacher|28226|1|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502827199|31|0|2|502367677|31|0|2|500589764|2||-2||2|2|500000294|500000294|-2|500000294, 500004640|-2|0|10|||7464|9|||1|388387|-1|4|3|44
502861539|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-10|2012-11-16|Baseline|2012-01-04|2012-01-10|Complete|Done|4|3|2|1|2|3|2.5|||||||||3|4|3|2|3|3|3|||||||||4|4|4|4||||||4|3|5|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Red||Child/Family: Infraction of match rules/agency policies|10.2||1|1|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Asian||25|28105|Some College|Single|Business: Sales|28134|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502862935|31|0|2|502683556|4|0|2|500589768|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|388391|-1|4|3|44
502063945|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-21|2016-08-05|Followup|2013-10-21|2014-01-05|Expired|Late||||||||3|3|3|2|2|3|2.67|||||||||2|3|3|1|3|2|2.33||||||3|2|2|2.33|||||||3|2|4|2|2.75||||||||||4|4|4|4|4|3|2|3.57||||||3|4|3|3.33|||||1|4|2.5||||2|2|||||||Yellow||Volunteer: Time constraint|69.5||1|1|1|1|M|White||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community||Match Support|M|White||37|28205||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502064367|1|0|1|502295138|1|0|1|500478943|2||500004641||4|2|||-2||-2|0|5|||7496|10|||1|388529|189168|4|0|45
502635070|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-05|2012-08-31|Baseline|2012-01-05|2012-01-05|Complete|Done|3|1|2|2|4|4|2.67|||||||||1|4|4|2|2|3|2.67|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||1|1|1|1|1|1|1|1||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|7.9||1|1|1|1|M|Multi-race (Black & Hispanic)||14|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community|Amachi|RTBM|M|White||31|28202|Masters Degree|Single|Finance: Auditor|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500001281|502635764|38|0|1|502823119|1|0|1|500581061|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|388592|-1|4|3|44
500970264|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2013-06-17|Followup|2012-10-27|2012-11-30|Complete|Done|3|2|3|2|3|3|2.67|4|3|3|2|3|3|3|-11|3|4|3|4|3|3|3.33|2|4|3|3|2|3|2.83|17.67|4|4|4|4|4|4|4|4|0|3|3|3|3|3|2|3|3|3|2.75|9.09|4|4|4|4|4|4|4|4|4|4|4|4|4|4||||4|4|3|3.67|4|4|4|4|-8.25|3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Red|Amachi|Volunteer: Lost contact with child/agency|31.7||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Enrollment|M|Black||44|28269|Some High School|Single|Insurance||0|2|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|1|502250629|31|0|1|500478922|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||12183|14|1209|1|1|388658|189150|4|3|45
502173821|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2014-08-29|Followup|2012-11-18|2012-12-23|Complete|Done|4|3|3|3|4|4|3.5|4|1|1|1|4|4|2.5|40|3|4|4|3|3|4|3.5|3|4|4|3|3|4|3.5|0|4|4|4|4|4|4|4|4|0|5|5|3|3|4|5|5|4|4|4.5|-11.11|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|2|2|2|50|2|2|1|1|100|4|4||||Red|Amachi|Volunteer: Time constraint|45.3||2|2|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||32|28262|Masters Degree|Single|Finance: Banking|28262|3|11|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502174240|31|0|2|502264706|1|0|2|500491573|2||500003586||4|3|500000294|500000294|-2|500000294, 500004640|-2|7016|11|||7464|9|||1|388663|148526|4|3|45
502308593|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-23|2015-05-28|Followup|2012-11-23|2013-02-07|Expired|Late||||||||4|2|3|1|3|4|2.83|||||||||3|3|4|4|3|3|3.33||||||3|2|3|2.67|||||||3|4|5|2|3.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|3|2.5||||1|1|||||||Red||Child/Family: Moved|54.1||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||40|28278|Bachelors Degree|Married|Tech: Computer/Programmer||3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502309025|31|0|1|502262702|31|0|1|500492994|2||-2||4|3|||-2||-2|0|10|||12183|14|1209|1|1|388665|206463|4|0|45
502359051|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-28|2017-02-28|Followup|2012-10-28|2012-11-30|Complete|Done|4|3|4|3|4|4|3.67|||||||||3|4|3|3|3|4|3.33|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|76.1||1|1|1|1|F|Black||14|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||35|28213|Masters Degree|Married|Business: Clerical||3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502359489|31|0|2|502242295|31|0|2|500483954|2||500004772||4|3|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|10|||131|1|||1|388672||4|3|45
502610186|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-26|NaT|Baseline|2012-01-05|2012-03-26|Complete|Done|4|1|4|1|4|4|3|||||||||3|3|3|2|2|3|2.67|||||||||4|4|4|4||||||2|4|2|4|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|||59.7||1|1|1|1|F|Black||16|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Asian||35|28210|Masters Degree|Married|Arts, Entertainment, Sports|28202|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|502610737|31|0|2|502913393|4|0|2|500601697|2||-2||2|1|||-2||-2|6854|8|||7671|13|||1|388768|-1|4|3|44
502308197|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-03|2016-05-09|Followup|2012-12-03|2012-12-12|Complete|Done|3|4|4|1|4|3|3.17|||||||||1|4|4|2|1|4|2.67|||||||||4|4|4|4||||||5|2|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|2|3||||||3|4|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|65.2||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Enrollment|F|White||35|28210|Bachelors Degree|Living w/ Significant Other|Business: Sales|18034|2|7|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big AND Amachi|Match Support|277|60|598|500000170|500021785|502308629|31|0|2|502325667|1|0|2|500493122|2||500003586||4|1||500000294|-2|500000294, 500004901|-2|0|10|||7496|10|||1|388871||4|3|45
500496598|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-23|NaT|Followup|2013-10-23|2014-01-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi, Cabarrus County||100.7||2|2|1|1|M|White||15|Yes|Mother|28083|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi, Cabarrus County|Match Support|M|White||35|28083|Masters Degree|Single|Business: Mgt, Admin|28027|2|3|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500496849|1|0|1|501383928|1|0|1|500299090|2||500003586||2|2|500000294, 500016374|500000294, 500016374|-2|500016374|-2|34|2|||7464|9|||1|389197||4|0|45
502431042|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-10|2013-12-20|Followup|2013-02-10|2013-02-25|Complete|Done|4|2|2|3|3|4|3|3|4|2|3|4|4|3.33|-9.91|3|4|4|4|4|4|3.83|2|3|3|3|4|3|3|27.67|4|4|4|4|4|4|4|4|0|4|4|5|5|4.5|3|4|5|3|3.75|20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|34.3||1|1|1|1|F|Black||17|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||34|28226|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502431483|31|0|2|502447496|1|0|2|500515174|2||-2||4|2|500005291|500005291|-2||-2|0|10|||7464|9|||1|389412|240749|4|3|45
502673798|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-30|2014-04-24|Baseline|2012-01-10|2012-01-30|Complete|Done|4|1|1|3|4|4|2.83|||||||||1|1|3|2|1|4|2|||||||||4|4|3|3.67||||||5|5|3|3|4|||||||4|4|4|4|1|4|4|3.57||||||||||4|3|4|3.67||||||2|1|1.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|26.8||1|1|1|1|M|Black||17|No|Mother|28105|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|White||36|28173|Bachelors Degree|Separated|Business: Mgt, Admin|28110|15|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502674626|31|0|1|502860952|1|0|1|500590803|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|389961|-1|4|3|44
502338225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2016-05-26|Followup|2013-10-27|2013-11-18|Complete|Done|4|4|4|3|4|4|3.83|3|2|3|1|4|4|2.83|35.34|3|4||4|4|4||2|3|2|2|3|3|2.5||4|4|4|4|3|3|3|3|33.33|5|5|4|4|4.5|2|3|2|3|2.5|80|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|2|3|2.5|20|2|2|1|1|100|4|4||||Yellow|Project Big|Volunteer: Lost contact with child/agency|67||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|White||33|28227|Bachelors Degree|Single|Unknown||9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502338658|31|0|2|502312449|1|0|2|500483095|2||500004641||4|2|500004640|500004640|-2|500004640|-2|0|4|||7496|10|||1|390183|194054|4|3|45
502725777|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2015-08-30|Baseline|2012-01-11|2012-01-23|Complete|Done|3|3|2|3|1|4|2.67|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||3|5|3|3|3.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Red|Amachi|Volunteer: Moved|43.2||1|1|1|1|F|Black||17|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||31|28217||Single|Customer Service||0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502726673|31|0|2|502710032|31|0|2|500590950|2||-2||4|3|500000294|500000294|-2||-2|34|2|||7464|9|||1|390244|-1|4|3|44
502860019|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-02-24|Baseline|2012-01-11|2012-02-22|Complete|Done|3|3|4|3|3|4|3.33|||||||||2|4|4|4|3|4|3.5|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||2|1|1.5|||||1|1||||4|4||||Green||Volunteer: Time constraint|24.1||1|1|1|1|F|Hispanic||19|No|Mother|28213|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|White||36|28205|Bachelors Degree||Tech: Engineer|28204|1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502861418|3|0|2|502873149|1|0|2|500596129|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|390412|-1|4|3|44
502627466|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-18|2014-05-15|Baseline|2012-01-11|2012-01-18|Complete|Done|3|3|4|2|2|4|3|||||||||4|4|4|2|4|4|3.67|||||||||4|3|4|3.67||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|4|3.5|||||1|1||||4|4||||Green||Volunteer: Moved|27.9||1|1|1|1|M|Hispanic|Mexican|18|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Multi-race (Hispanic & White)||28|28202|Bachelors Degree|Single|Finance||0|3|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502628116|3|10|1|502800101|35|0|1|500591158|2||-2||4|1|||-2||-2|0|4|||7438|1|||1|390452|-1|4|3|44
502745717|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-12|2013-02-28|Followup|2013-01-12|2013-01-31|Declined|Done||||||||3|1|4|1|4|4|2.83|||||||||2|4|4|2|2|4|3||||||4|4|4|4|||||||3|4|3|5|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||4|2|3||||2|2||||4|4||Red||Child/Family: Lost contact with volunteer/agency|13.6||1|1|1|1|F|Multi-race (Black & White)||17|No|Mother|28278|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|F|Asian||34|28278|Bachelors Degree|Single|Govt|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|502746625|36|0|2|502712044|4|0|2|500583497|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|390718|376817|4|1|45
500186260|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-29|2015-12-17|Followup|2013-10-29|2014-01-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|133.6||3|3|1|1|M|Black||19|No|Mother|28025|One Parent: Female|Unknown||No||Self|General Site||Match Support|M|Black||42|28025|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|500187857|31|0|1|500189139|31|0|1|500037139|2||-2||4|2|||-1||-2|0|10|||7464|9|||1|390952||4|0|45
501361902|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-23|NaT|Followup|2013-01-23|2013-03-13|Complete|Late|4|3|3|3|3|3|3.17|||||||||3|2|3|3|3|3|2.83|||||||||4|4|4|4||||||3|4|5|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||4|3|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi||97.7||1|1|1|1|M|White||17|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28227|Bachelors Degree|Divorced|Business: Sales|28273|9|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501249611|1|0|1|501307192|1|0|1|500328424|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|391037||4|3|45
502571727|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-13|2017-03-09|Followup|2013-01-13|2013-03-30|Expired|Late||||||||3|4|4|3|1|4|3.17|||||||||2|4|2|3|4|3|3||||||4|4|4|4|||||||4|3|4|5|4||||||||||4|4|4|4|3|4|4|3.86||||||4|4|2|3.33|||||3|4|3.5||||2|2||||4|4||Green||Volunteer: Lost contact with child/agency|61.8||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|M|Black||45|28207|Masters Degree|Married|Tech: Management|28081|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|502572181|31|0|1|502769619|31|0|1|500586830|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|391144|382185|4|0|45
502830103|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-31|2012-05-31|Baseline|2012-01-13|2012-01-31|Complete|Done|4|4|4|4|4|4|4|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|3|4|4|4|4|4|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Red||Volunteer: Moved|4||1|1|1|1|F|Hispanic||16|No|Mother|28213|One Parent: Female|Less than $10,000||Yes||Self|General Community|Amachi|RTBM|F|White||28|28205|Bachelors Degree|Single|Retail: Mgt|28056|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502831393|3|0|2|502819928|1|0|2|500592797|2||-2||4|3||500000294|-2||-2|0|10|||7464|9|||1|391205|-1|4|3|44
502507408|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-13|2016-08-22|Followup|2012-10-13|2012-11-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|58.3||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Less than $10,000||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||71|28277|Bachelors Degree|Married|Retired||0|0||Relative|Big|General Community||Match Support|277|60|598|500000170|500017732|502507857|31|0|1|502673562|31|0|1|500559678|2||-2||4|2|500005291||-2||-2|34|2|||0|11|||1|391372||4|1|45
501092957|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-09|2014-05-15|Followup|2012-11-09|2013-01-09|Complete|Late|3|2|2|3|2|2|2.33|||||||||4|4|4|1|2|4|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|42.2||2|2|1|1|M|Black||17|No|Mother|28027|One Parent: Female|$30,000 to $34,999||No|Radio|Media|General Community||Match Support|M|White||44|28269||Married|Finance: Banking||5|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|501093231|31|0|1|502294662|1|0|1|500484597|2||-2||4|1|||-2||-2|55|1|||7459|10|||1|391783||4|3|45
501060196|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-26|2015-08-03|Followup|2012-11-26|2012-12-12|Complete|Done|4|4|4|3|3|4|3.67|||||||||2|3|2|3|2|2|2.33|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|3|3|4|3|3|3.43||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green||Child/Family: Moved|92.2||1|1|1|1|M|Black||19|No|Mother|28205|One Parent: Female|$15,000 to $19,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28226|Masters Degree|Single|Finance: Accountant||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501060469|31|0|1|501036081|1|0|1|500223215|2||-2||4|1|||-2||-2|34|2|||46|2|||1|391959||4|3|45
502627466|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-18|2014-05-15|Followup|2014-01-18|2014-02-03|Complete|Done|4|3|3|3|4|4|3.5|3|3|4|2|2|4|3|16.67|3|4|4|2|3|4|3.33|4|4|4|2|4|4|3.67|-9.26|4|4|4|4|4|3|4|3.67|8.99|5|3|3|4|3.75|5|4|3|5|4.25|-11.76|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|2|3.33|3|4|4|3.67|-9.26|3|3|3|3|4|3.5|-14.29|1|1|1|1|0|4|4|4|4|0|Green||Volunteer: Moved|27.9||1|1|1|1|M|Hispanic|Mexican|18|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Multi-race (Hispanic & White)||28|28202|Bachelors Degree|Single|Finance||0|3|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502628116|3|10|1|502800101|35|0|1|500591158|2||-2||4|1|||-2||-2|0|4|||7438|1|||1|392249|390452|4|3|45
501428903|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-21|2015-02-25|Followup|2013-01-21|2013-04-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|73.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|White||53|15001|Masters Degree|Single|Consultant|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501429188|31|0|1|501441245|1|0|1|500331206|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|393057||4|0|45
502627468|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-17|2014-05-19|Baseline|2012-01-20|2013-05-17|Complete|Done|2|4|4|4|3|3|3.33|||||||||4|2|2|3|4|4|3.17|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Lost interest|12.1||1|1|1|1|M|Hispanic|Mexican|18|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||30|28036|Some College|Single|Business|28078|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500017777|502628116|3|10|1|503419352|1|0|1|500696276|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|393156|-1|4|3|44
502197477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-10|2016-10-03|Followup|2013-02-10|2013-04-27|Expired|Late||||||||4|3|4|4|4|4|3.83|||||||||2|3|3|4|3|3|3||||||3|3|3|3|||||||5|3|3|5|4||||||||||4|4|4|3|3|4|4|3.71||||||4|4|3|3.67|||||4|4|4||||1|1||||4|4||Green|2010-2012 OJJDP JJI|Volunteer: Moved|67.7||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28202|Bachelors Degree|Single|Business: Sales|27560|1|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017732|502197915|31|0|1|502422929|1|0|1|500515536|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|4|||7464|9|||1|393171|241218|4|0|45
500340183|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-18|2013-08-30|Followup|2012-12-18|2013-02-04|Complete|Late|3|2|2|1|3|3|2.33|||||||||1|4|4|1|2|4|2.67|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|44.4||3|3|1|1|M|Black||17|No|Relative: Other|28208|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction||0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|500340317|31|0|1|501933993|1|0|1|500419988|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|393311||4|3|45
501069450|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-07|2017-02-28|Followup|2013-11-07|2014-01-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|111.7||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||66|28075||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501048131|31|0|1|500887364|31|0|1|500212043|2||-2||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|393503||4|0|45
501786018|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2013-06-28|Followup|2013-01-23|2013-01-09|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|3|3|4|4|3|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Moved|17.1||4|4|1|1|M|Black||17|Yes|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Asian||28|28203||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|501786373|31|0|1|502800403|4|0|1|500589712|2||500003586||4|3|500000294||-2||-2|0|10|||7496|10|||1|393631||4|3|45
502725760|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2014-09-24|Followup|2013-01-23|2013-03-25|Declined|Late||||||||4|4|4|4|4|4|4|||||||||2|4|4|2|4|4|3.33||||||4|4|4|4|||||||5|4|4|5|4.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|2|3||||2|2||||4|4||Yellow|Amachi|Volunteer: Lost contact with child/agency|32||1|1|1|1|M|Black||16|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|Amachi|Match Support|M|Black||28|28226|Bachelors Degree|Single|Business: Sales|28217|0|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502726656|31|0|1|502687867|31|0|1|500589763|2||-2||4|2|500000294|500000294|-2||-2|0|10|||4748|14|633|1|1|393654|388386|4|1|45
502725777|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2015-08-30|Followup|2013-01-23|2013-03-25|Declined|Late||||||||3|3|2|3|1|4|2.67|||||||||3|4|4|4|4|4|3.83||||||4|4|4|4|||||||3|5|3|3|3.5||||||||||4|4|4|4|4|4|2|3.71||||||4|4|3|3.67|||||4|4|4||||1|1||||4|4||Red|Amachi|Volunteer: Moved|43.2||1|1|1|1|F|Black||17|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||31|28217||Single|Customer Service||0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502726673|31|0|2|502710032|31|0|2|500590950|2||-2||4|3|500000294|500000294|-2||-2|34|2|||7464|9|||1|393670|390244|4|1|45
502825916|BBBS of Greater Charlotte|Main Office|C|Active|2012-01-23|NaT|Followup|2013-01-23|2013-03-25|Declined|Late||||||||4|2|1|2|2|4|2.5|||||||||2|3|4|3|4|3|3.17||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||4|4|4||||2|2||||4|4||Yellow|Amachi||61.7||1|1|2|2|F|Black||14|Yes|Mother|28273|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28208|Some College|Single|Education: Teacher|28226|1|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502827199|31|0|2|502367677|31|0|2|500589764|2||-2||2|2|500000294|500000294|-2|500000294, 500004640|-2|0|10|||7464|9|||1|393702|388387|4|1|45
500337327|BBBS of Greater Charlotte|Main Office|C|Active|2006-12-14|NaT|Followup|2013-12-14|2013-12-23|Complete|Done|4|4|4|1|1|1|2.5|||||||||2|4|3|4|2|3|3|||||||||4|4|4|4||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||123||2|3|4|5|M|Black||16||GrandMother|28208|Grandparents|Unknown||No||School|General Site||Match Support|M|Black||49|28217|Associate Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site||Match Support|277|60|598|500000170|500017732|500251937|31|0|1|500189300|31|0|1|500148262|2||-2||2|1|||-1||-1|0|4|||7464|9|||1|393719||4|3|45
501904094|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-15|2013-06-19|Followup|2013-01-15|2013-04-01|Expired|Late||||||||4|1|4|2|4|4|3.17|||||||||2|4|4|3|4|4|3.5||||||4|4|4|4|||||||3|4|2|5|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Red||Volunteer: Lost contact with child/agency|41.1||1|1|1|1|F|Black||16|No|Mother|28214|One Parent: Female|Unknown|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||56|28208|Some College|Single|Finance: Accountant|28203|19|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500004169|501904482|31|0|2|501342148|31|0|2|500420809|2||-2||4|3|||-2|500000294|-2|34|2|||7446|3|||1|393772|23717|4|0|45
501454635|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-19|2013-09-30|Followup|2013-01-19|2013-02-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|44.4||1|1|2|2|M|Black||15|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Some Other Race||40|28216|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|501454920|31|0|1|500188923|41|0|1|500424889|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|393800||4|1|45
502244776|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-19|NaT|Followup|2013-01-19|2013-02-06|Complete|Done|4|2|1|2|4|3|2.67|4|2|2|1|3|4|2.67|0|2|4|4|2|3|3|3|2|3|3|2|3|2|2.5|20|4|3|4|3.67|4|3|2|3|22.33|5|5|5|5|5|2|3|3|4|3|66.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|2|4|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|2010-2012 OJJDP JJI||73.9||1|1|2|2|F|Black||16|No|Mother|28216|Two Parent|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28209|Bachelors Degree|Single|Law|28273|5|0|Relative|Relative|Big|General Community|Amachi|Match Support|277|60|598|500000170|500021785|502245202|31|0|2|502143351|1|0|2|500511171|2||-2||2|1|500005291|500005291|-2|500000294|-2|0|4|||17161|11|||1|393963|233727|4|3|45
501529921|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2015-04-06|Followup|2013-01-23|2013-01-28|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|4|2|4|3.17|||||||||4|4|4|4||||||3|1|5|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|38.4||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||48|28031|Some College|Divorced|Medical|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501530213|31|0|2|502554719|1|0|2|500581908|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|393998||4|3|45
500791567|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-31|2013-04-11|Followup|2013-01-31|2013-02-06|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|4|2|4|4|3.5|||||||||4|3|3|3.33||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow||Volunteer: Time constraint|74.3||1|1|2|2|M|Multi-Race (None of the above)||18|No|Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|M|Black||32|28215||Married|Finance: Banking||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|500187654|7|0|1|500578720|31|0|1|500155823|2||-2||4|2|||-2||-2|0|10|||7447|3|||1|394344||4|3|45
502335675|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-30|2016-10-31|Followup|2012-12-30|2013-02-09|Complete|Done|3|3|3|2|4|4|3.17|||||||||3|4|4|3|4|3|3.5|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi|Child: Lost interest|70||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|Project Big AND Amachi|Match Support|M|White||27|28262||Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502336110|31|0|1|502305990|1|0|1|500495220|2||500004772||4|3|500000294, 500004640, 500004901|500004901|-2|500000294, 500004640|-2|0|4|||7496|10|||1|394443||4|3|45
502188863|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-31|2013-10-31|Followup|2012-12-31|2013-02-09|Complete|Done|3|3|4|2|3|4|3.17|4|2|3|2|3|3|2.83|12.01|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|4|4|4|4|4|25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|4|2|3|16.67|2|2|1|1|100|4|4||||Red|Project Big|Volunteer: Moved|34||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|M|Some Other Race||30|28202|Some College|Single|Tech: Support, Writing|28210|0|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502189292|31|0|1|502288935|41|0|1|500498784|2||-2||4|3|500004640|500004640|-2|500004640|-2|0|10|||46|2|||1|394458|191872|4|3|45
500847570|BBBS of Greater Charlotte|Main Office|C|Active|2012-01-25|NaT|Followup|2013-01-25|2013-01-30|Complete|Done|4|1|2|1|3|3|2.33|||||||||4|4|4|1|2|4|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Yellow|Amachi||61.7||2|2|1|1|F|Black||16|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||52|28227|Bachelors Degree|Married|Insurance|28277|14|0|AA Task Force|Special Event|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188056|31|0|2|502542379|31|0|2|500592215|2||500003586||2|2|500000294|500000294|-2|500000294|-2|0|10|||11098|8|||1|394660||4|3|45
502888277|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-31|2012-08-29|Baseline|2012-01-25|2012-01-31|Complete|Done|3|3|3|2|3|2|2.67|||||||||2|3|2|2|2|3|2.33|||||||||4|4|4|4||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Child: Lost interest|6.9||1|1|1|1|M|Black||18|Yes|Mother|28205|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||63|28269|Bachelors Degree|Married|Business: Sales||9|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502889684|31|0|1|502853546|1|0|1|500593701|2||500003586||4|3|500000294|500000294|-2||-2|6854|8|||7464|9|||1|394807|-1|4|3|44
502787524|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-25|2014-08-29|Followup|2013-01-25|2013-03-06|Complete|Done|4|3|4|3|4|4|3.67|3|4|4|4|4|4|3.83|-4.18|3|4|4|4|4|4|3.83|2|4|3|4|4|4|3.5|9.43|4|4|4|4|4|3|3|3.33|20.12|4|5|5|4|4.5|4|5|5|5|4.75|-5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|3|3.5|4|4|4|-12.5|2|2||||4|4|4|4|0|Red||Child/Family: Lost contact with volunteer/agency|31.1||1|1|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28205|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Asian||29|28202||Single|Tech: Computer/Programmer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502788707|38|0|2|502272989|4|0|2|500587325|2||-2||4|3|||-2|500004640|-2|0|10|||7496|10|||1|394867|382987|4|3|45
502732602|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-25|2013-06-18|Followup|2013-01-25|2013-02-09|Declined|Done||||||||4|2|4|1|1|4|2.67|||||||||2|2|3|4|3|4|3||||||4|4|4|4|||||||3|3|5|3|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||1|1|1||||2|2||||4|4||Yellow||Volunteer: Moved|16.8||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|White||29|28203|Masters Degree|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502733499|31|0|2|502766077|1|0|2|500588408|2||-2||4|2||500005291|-2||-2|0|5|||7464|9|||1|394874|385114|4|1|45
500185865|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-15|2014-08-20|Followup|2012-12-15|2013-03-01|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|68.1||2|2|2|2|F|Black||19||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187761|31|0|2|500189140|31|0|2|500326656|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|395240||4|0|45
500914579|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-16|2014-12-04|Followup|2012-12-16|2013-01-23|Complete|Done|3|2|2|2|3|2|2.33|||||||||1|3|3|1|2|3|2.17|||||||||2|2|2|2||||||1|3|2|1|1.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Yellow||Child: Severity of challenges|71.6||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|M|White||32|28277|Bachelors Degree|Single|Tech: Engineer|28117|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500914849|31|0|1|501345550|1|0|1|500323102|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|395241||4|3|45
500796255|BBBS of Greater Charlotte|Main Office|C|Active|2010-01-20|NaT|Followup|2013-01-20|2013-01-22|Complete|Done|3|2|1|1|1|3|1.83|||||||||4|4|4|4|4|4|4|||||||||3|3|3|3||||||5|3|3|2|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||3|2|2.5|||||2|2||||4|4||||Green|||85.8||3|3|1|1|M|White||18|No|Mother|28031|One Parent: Male|$20,000 to $24,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||60|28269|||Medical: Admin|28207|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500796529|1|0|1|501846438|1|0|1|500424314|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|395352||4|3|45
502875276|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-06|2013-06-06|Baseline|2012-01-26|2012-02-06|Complete|Done|4|3|3|3|4|3|3.33|||||||||3|3|3|3|2|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|2|2.5|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|16||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Enrollment|M|White||30|28031|Bachelors Degree|Single|Finance|28027|1|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502876679|31|0|1|502877270|1|0|1|500594084|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|395401|-1|4|3|44
500185601|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-28|2015-07-23|Followup|2013-01-28|2013-03-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|89.8||2|2|1|1|M|Black||20||Mother|28210|Other/Unknown|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28078|High School Graduate|Single|Finance: Accountant|28202|0|4|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500187235|31|0|1|501082220|1|0|1|500236473|2||-2||4|1|||-2||-2|6854|8|||7458|9|||1|395427||4|1|45
501516900|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-28|2015-08-27|Followup|2013-01-28|2013-03-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|78.9||1|1|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||39|28212|Bachelors Degree|Single|Medical: Healthcare Worker|28210|1|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500018987|501517192|31|0|2|501438601|31|0|2|500332399|2||-2||4|1|||-2||-2|6854|8|||7462|13|||1|395432||4|1|45
502340295|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-23|2012-03-16|Baseline|2012-01-26|2012-02-23|Complete|Done|3|2|2|2|2|2|2.17|||||||||3|3|3|2|3|3|2.83|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|||||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|0.7||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Single|Business: Marketing|28036|5|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502340731|31|0|1|502881673|1|0|1|500594127|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|395445|-1|4|3|44
502666840|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-17|2013-02-27|Baseline|2012-01-27|2012-02-17|Complete|Done|3|2|4|1|4|4|3|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|12.4||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$20,000 to $24,999||Yes|Arby's|Workplace Partner/Business|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||49|28173|Bachelors Degree|Single|Insurance|28210|21|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502667667|31|0|1|502872585|31|0|1|500594266|2||-2||4|3||500005291|-2||-2|3394|14|||7496|10|||1|395754|-1|4|3|44
502469903|BBBS of Greater Charlotte|Main Office|C|Active|2012-02-22|NaT|Baseline|2012-01-27|2012-02-18|Complete|Done|3|4|4|3|3|4|3.5|||||||||3|4|3|3|3|3|3.17|||||||||3|4|4|3.67||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||1|1||||4|4||||Green|||60.7||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$15,000 to $19,999|Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||34|28269|Bachelors Degree|Single|Business: Human Resources|28025|2|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500020910|502470350|31|0|1|502868874|31|0|1|500594396|2||-2||2|1|||-2||-2|0|5|||4748|14|1360|3|1|395896|-1|4|3|44
500261295|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-21|2017-03-09|Followup|2012-12-21|2013-02-28|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|134.6||1|1|1|1|M|White||20||Mother|28104|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||60|28270|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500261310|1|0|1|500188435|1|0|1|500073081|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|395950||4|1|45
502211307|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-03|2014-04-24|Followup|2013-02-03|2013-03-18|Declined|Done||||||||4|4|4|3|4|3|3.67|||||||||4|3|3|4|3|3|3.33||||||4|4|4|4|||||||4|4|4||||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4||||||3|||||2|2|||||||Yellow|Amachi|Volunteer: Time constraint|38.6||1|1|1|1|M|Black||16|Yes|Mother|28278|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||51|28214|Bachelors Degree|Single|Business: Sales|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502211737|31|0|1|502371462|1|0|1|500512414|2||-2||4|2|500000294|500000294|-2|500000294|-2|7016|11|||7496|10|||1|395953|177660|4|1|45
501536365|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-03|2014-07-17|Followup|2013-02-03|2013-02-01|Complete|Done|4|1|4|1|4|4|3|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|1|4|4|3.57||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|65.4||1|1|1|1|M|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Enrollment|M|Black||57|28105|Some College|Married|Retail: Sales|28105|10|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501536657|31|0|1|501443152|31|0|1|500336020|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|396299||4|3|45
502673798|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-30|2014-04-24|Followup|2013-01-30|2013-02-04|Complete|Done|2|2|3|2|3|3|2.5|4|1|1|3|4|4|2.83|-11.66|2|2|3|2|2|2|2.17|1|1|3|2|1|4|2|8.5|3|2|2|2.33|4|4|3|3.67|-36.51|1|4|4|4|3.25|5|5|3|3|4|-18.75|4|4|4|4|3|4|4|3.86|4|4|4|4|1|4|4|3.57|8.12|3|3|3|3|4|3|4|3.67|-18.26|3|2|2.5|2|1|1.5|66.67|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Time constraint|26.8||1|1|1|1|M|Black||17|No|Mother|28105|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|White||36|28173|Bachelors Degree|Separated|Business: Mgt, Admin|28110|15|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502674626|31|0|1|502860952|1|0|1|500590803|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|396641|389961|4|3|45
501201377|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-31|2016-08-26|Followup|2013-01-31|2013-02-04|Complete|Done|3|3|3|2|3|3|2.83|||||||||4|4|4|3|3|4|3.67|||||||||4|4|3|3.67||||||5|5|4|4|4.5|||||||4|4|4|3|4|3|3|3.57||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|90.8||1|1|1|1|F|Hispanic||18|No|Mother|28212|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community||Match Support|F|Hispanic||65|28269|Masters Degree|Single|Medical: Admin|28262|8|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500017777|501201651|3|0|2|501497622|3|0|2|500331903|2||-2||4|3|||-2||-2|7016|11|||7446|3|||1|398090||4|3|45
501347056|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2015-10-12|Followup|2012-12-12|2013-02-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|82||1|1|1|1|M|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28226|Bachelors Degree|Married|Tech: Engineer|28202|2|8|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|501347335|31|0|1|501217000|1|0|1|500322327|2||-2||4|2|||-2||-2|34|2|||7446|3|||1|398095||4|1|45
500185897|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-05|2014-01-31|Followup|2013-02-05|2013-03-06|Complete|Done|3|2|4|2|3|3|2.83|||||||||2|3|2|4|4|3|3|||||||||3|4|4|3.67||||||2|3|4|4|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|2|2|2.33||||||3|2|2.5|||||2|2||||4|4||||Red|Project Big|Child: Graduated|83.8||2|2|1|1|M|Black||21|No|Relative: Other|28208|Other Relative|Unknown||No||Self|General Community||Match Support|M|White||39|28277|Bachelors Degree|Single|Tech: Computer/Programmer||4|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500008321|500187458|31|0|1|500549520|1|0|1|500155451|2||500004641||4|3|500004640||-2||-2|0|10|||46|2|||1|398378||4|3|45
502225378|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-26|NaT|Followup|2013-01-26|2013-02-26|Complete|Done|4|4|4|2|1|4|3.17|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||73.6||1|1|1|1|M|White||14|No|Mother|28277|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||67|28277|Bachelors Degree|Divorced|Tech: Sales, Mktg||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|502225809|1|0|1|502245842|1|0|1|500509780|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|399169||4|3|45
502875276|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-06|2013-06-06|Followup|2013-02-06|2013-01-26|Complete|Done|3|1|1|1|1|1|1.33|4|3|3|3|4|3|3.33|-60.06|2|4|4|4|4|4|3.67|3|3|3|3|2|3|2.83|29.68|4|4|4|4|4|4|4|4|0|2|4|4|3|3.25|3|3|3|3|3|8.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|3|3|3|11|2|3|2.5|3|2|2.5|0|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Lost contact with child/agency|16||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Enrollment|M|White||30|28031|Bachelors Degree|Single|Finance|28027|1|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502876679|31|0|1|502877270|1|0|1|500594084|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|399365|395401|4|3|45
502824908|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-21|2015-07-22|Baseline|2012-02-06|2012-02-20|Complete|Done|3|2|3|2|3|3|2.67|||||||||3|4|4|2|2|3|3|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|41||1|1|1|1|F|Black||19|No|Mother|28226|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community||Match Support|F|White||34|28226|Bachelors Degree|Married|Unknown|29715|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502826191|31|0|2|502891382|1|0|2|500596373|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|399457|-1|4|3|44
501389722|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-06|2014-04-24|Followup|2013-02-06|2013-01-09|Complete|Early|1|2|4|1|3|3|2.33|||||||||1|3|4|2|1|4|2.5|||||||||3|3|3|3||||||3|4|2|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Green||Child: Graduated|62.5||1|1|1|1|F|White||21|No|Mother|28027|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||56|28027||Divorced|Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500012459|501390003|1|0|2|500787778|1|0|2|500337267|2||-2||4|1|||-2||-2|0|10|||46|2|||1|399898||4|3|45
501811395|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-10|NaT|Followup|2013-03-10|2013-02-12|Complete|Early|4|4|4|1|4|1|3|||||||||2|4|3|1|1|4|2.5|||||||||2|3|4|3||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|Cabarrus County||84.2||1|1|1|1|F|Black||15|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||60|28213||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501811730|31|0|2|500876892|31|0|2|500436702|2||500016307||2|1|500016374|500016374|-2|500016374|-2|6854|8|||2238|7|||1|399906||4|3|45
502753873|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-29|2013-02-22|Baseline|2012-02-07|2012-02-29|Complete|Done|3|3|3|3|4|4|3.33|||||||||3|2|3|3|2|3|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|11.8||2|2|1|1|F|Hispanic||14|No|Mother|28262|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||27|28269|Bachelors Degree|Single|Finance|28227|0|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|502751081|3|0|2|502896683|31|0|2|500596765|2||-2||4|2|||-2||-2|0|10|||46|2|||1|399995|-1|4|3|44
502875778|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-10|2013-03-29|Baseline|2012-02-08|2012-02-10|Complete|Done|3|4|4|2|4|4|3.5|||||||||4|1|4|4|2|4|3.17|||||||||4|4|4|4||||||3|5|2|2|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Feels incompatible with child/family|13.6||1|1|1|1|F|Black||18|Yes|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||44|28216|Associate Degree|Divorced|Finance: Banking||0|5|Charlotte Cares|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502877181|31|0|2|502885755|31|0|2|500597009|2||-2||4|3|500000294|500000294|-2||-2|0|10|||11246|6|||1|400385|-1|4|3|44
502859187|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-14|2012-05-31|Baseline|2012-02-08|2012-03-14|Complete|Done|2|2|4|2|4|4|3|||||||||2|3|3|3|3|4|3|||||||||4|4|4|4||||||4|5|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|2.6||2|2|2|2|F|Black||15|No|GrandMother|28205|Grandparents|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|White||28|28213|Bachelors Degree|Single|Medical: Nurse||0|4|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|500187987|31|0|2|502849360|1|0|2|500597086|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|400467|-1|4|3|44
501132052|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-08|2015-10-15|Followup|2013-02-08|2013-03-23|Complete|Done|3|1|4|1|4|4|2.83|||||||||1|3|4|4|4|4|3.33|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|44.2||2|3|1|2|F|Black||17||Mother|28213|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||35|85254|Bachelors Degree|Married|Medical: Admin|28217|2|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500018987|501076355|31|0|2|501356464|1|0|2|500597097|2||-2||4|1|||-2||-2|0|4|||7446|3|||1|400480||4|3|45
502317500|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-08|2015-07-31|Followup|2013-02-08|2013-03-07|Complete|Done|3|2|2|2|3|3|2.5|4|2|1|2|4|4|2.83|-11.66|2|3|3|3|3|3|2.83|2|3|4|2|2|4|2.83|0|4|4|3|3.67|4|4|4|4|-8.25|4|3|4|4|3.75|4|3|2|3|3|25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|3|2|2.67|3|4|3|3.33|-19.82|2|3|2.5|3|2|2.5|0|2|2|2|2|0|4|4|4|4|0|Red|Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|41.7||1|1|2|2|M|Black||15|No|Mother|28214|One Parent: Female|Unknown||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|M|White||33|28214|Associate Degree|Single|Law: Security Officer|28208|2|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502317931|31|0|1|502658498|1|0|1|500587614|2||-2||4|3|500004640, 500004901|500004640, 500004901|-2||-2|0|4|||7464|9|||1|400549|383492|4|3|45
502671406|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-14|2014-09-04|Baseline|2012-02-09|2012-02-13|Complete|Done|3|4|4|3|3|3|3.33|||||||||3|3|2|3||3||||||||||3|3|3|3||||||1|3|3|3|2.5|||||||4|4|4|4|2|4|4|3.71||||||||||3|4|4|3.67||||||3|1|2|||||1|1||||4|4||||Yellow||Volunteer: Infraction of match rules/agency policies|30.7||1|1|1|1|F|Black||19|No|Mother|28210|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||34|28226|PHD|Single|Medical: Healthcare Worker|28207|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502672234|31|0|2|502885637|31|0|2|500597397|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|400951|-1|4|3|44
500186071|BBBS of Greater Charlotte|Main Office|C|Completed|2004-01-05|2014-04-30|Followup|2013-01-05|2013-02-18|Complete|Done|4|3|3|2|3|4|3.17|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|123.8||1|1|1|1|M|White||21|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||40|28277|Masters Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187670|1|0|1|500189012|1|0|1|500037012|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|400968||4|3|45
500717519|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-08|2013-08-29|Followup|2012-12-08|2013-01-09|Complete|Done|3|2|3|2|3|3|2.67|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Child: Lost interest|80.7||1|1|2|2|M|Black||20||Mother|28205|One Parent: Female|$20,000 to $24,999|Y|No||School|General Community||Match Support|M|Black||37|28269|Bachelors Degree|Married|Education: Admin||0|0|Yahoo!|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011746|500717786|31|0|1|500188838|31|0|1|500145722|2||-2||4|2|||-2||-2|0|4|||32|2|||1|401183||4|3|45
502083429|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-11|2016-08-19|Followup|2013-02-11|2013-01-02|Complete|Early|4|4|4|3|4|4|3.83|4|2|4|3|2|4|3.17|20.82|3|1|3|3|3|3|2.67|4|4|4|1|4|4|3.5|-23.71|4|4|4|4|4|3|3|3.33|20.12|4|5|3|4|4|3|5|4|4|4|0|4|4|4|4|4|3|3|3.71|4|2|4|4|4|4|3|3.57|3.92|3|4|3|3.33|4|4|4|4|-16.75|4|3|3.5|3|3|3|16.67|1|1|2|2|-50|4|4|4|4|0|Red||Volunteer: Moved|54.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Cabarrus County|Match Support|F|Black||29|28027|Bachelors Degree|Single|Education: Teacher||1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|502083853|31|0|2|502653045|31|0|2|500590992|2||-2||4|3||500016374|-2|500016374|-2|7016|11|||7464|9|||1|401514|220254|4|3|45
500636617|BBBS of Greater Charlotte|Main Office|C|Completed|2007-01-10|2013-08-20|Followup|2013-01-10|2013-03-27|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|79.3||2|2|1|1|M|Black||17||Mother|28269|One Parent: Female|$20,000 to $24,999|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28262||Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500636863|31|0|1|500756919|31|0|1|500151137|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|401577||4|0|45
501222138|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2015-05-07|Followup|2012-04-30|2012-04-30|Complete|Done|4|2|3|1|2|4|2.67|||||||||2|2|3|2|2|3|2.33|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|60.2||2|2|2|3|F|Black||14|Yes|GrandMother|28227|Grandparents|Unknown||No||Self|General Community|Amachi|Enrollment|F|Black||53|28269|Some College|Married|Business: Sales|28227|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501222414|31|0|2|500189173|31|0|2|500447311|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|401596||4|3|45
502336272|BBBS of Greater Charlotte|Main Office|C|Completed|2011-01-07|2013-11-21|Followup|2013-01-07|2012-12-18|Complete|Early|1|4|4|2|1|3|2.5|||||||||4|1|1|4|4|1|2.5|||||||||1|1|1|1||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|34.5||2|2|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||31|28208|Bachelors Degree|Single|Business: Sales||0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502336707|31|0|2|502363052|31|0|2|500502396|2||-2||4|2|||-2||-2|6854|8|||7464|9|||1|401622||4|3|45
502472483|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2014-08-28|Followup|2013-02-28|2013-04-12|Blank|Done||||||||3|1|4|4|1|1|2.33|||||||||2|2|3|3|4|3|2.83||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|3|4|3|3.71||||||4|4|4|4|||||2|3|2.5||||1|1|||||||Red|Amachi|Volunteer: Time constraint|42||1|1|1|1|F|Black||18|Yes|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi|Match Support|F|White||33|28202|Bachelors Degree|Single|Education|28208|4|10|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013781|502472930|31|0|2|502453698|1|0|2|500518061|2||500003586||4|3|500000294|500000294|-2|500004640|-2|0|10|||7464|9|||1|401675|245268|4|3|45
501390344|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-26|NaT|Followup|2013-02-26|2013-02-07|Complete|Early|4|4|2|2|2|4|3|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|2|3|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi||96.6||1|1|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Single|Tech: Computer/Programmer||0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|501390617|31|0|1|501380163|1|0|1|500342682|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|401727||4|3|45
502859440|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-01|2014-04-21|Baseline|2012-02-13|2012-08-01|Complete|Done|3|2|3|1|3|3|2.5|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||1|1||||4|4||||Green||Volunteer: Time constraint|20.6||1|1|1|1|F|Hispanic|Mexican|15|No|Mother|28215|Two Parent|Unknown||Yes||School|General Community||Match Support|F|Multi-race (Hispanic & White)||30|28202|Bachelors Degree|Married|Finance: Banking|28255|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502860839|3|10|2|503046471|35|0|2|500623399|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|401855|-1|4|3|44
501735420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2015-08-13|Followup|2013-01-26|2013-02-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|66.5||2|2|2|2|F|Black||16||GrandMother|28215|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||41|28277|Bachelors Degree|Single|Business: Mgt, Admin||9|0|General|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500017732|501735760|31|0|2|500956022|1|0|2|500428818|2||-2||4|1|||-2||-2|6854|8|||6450|12|||1|401927||4|1|45
502551045|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-03-06|Baseline|2012-02-13|2012-02-20|Complete|Done|4|1|1|2|1|4|2.17|||||||||1|1|2|2|1|2|1.5|||||||||1|2|2|1.67||||||2|2|2|2|2|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|2|3||||||2|2|2|||||1|1||||4|4||||Yellow||Volunteer: Health|24.4||2|2|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||54|28031|Bachelors Degree|Married|Business: Mgt, Admin|28262|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502551498|31|0|2|502864071|1|0|2|500597976|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|401956|-1|4|3|44
501045214|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-30|2015-12-16|Followup|2013-11-30|2014-02-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|96.5||1|1|2|2|F|Black||20|No|Relative: Other|28269|Grandparents|$20,000 to $24,999||Yes||BBBS Board/Staff|General Community||Match Support|F|Black||35|28213|Masters Degree|Single|Business||4|0|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|277|60|598|500000170|500002335|501045484|31|0|2|500953330|31|0|2|500217682|2||-2||4|1|||-2|500014505, 500016394|-1|0|13|||46|2|||1|402076||4|0|45
502671406|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-14|2014-09-04|Followup|2013-02-14|2013-01-22|Complete|Early|1|2|4|4|4|4|3.17|3|4|4|3|3|3|3.33|-4.8|2|3|3|2|2|3|2.5|3|3|2|3||3|||3|3|3|3|3|3|3|3|0|3|4|3|3|3.25|1|3|3|3|2.5|30|4|4|4|4|4|4|3|3.86|4|4|4|4|2|4|4|3.71|4.04|3|3|3|3|3|4|4|3.67|-18.26|1|1|1|3|1|2|-50|1|1|1|1|0|4|4|4|4|0|Yellow||Volunteer: Infraction of match rules/agency policies|30.7||1|1|1|1|F|Black||19|No|Mother|28210|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||34|28226|PHD|Single|Medical: Healthcare Worker|28207|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502672234|31|0|2|502885637|31|0|2|500597397|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|402157|400951|4|3|45
500186905|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-10|2015-11-04|Followup|2013-02-10|2013-03-12|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|3|4|2|3|2.83|||||||||4|4|4|4||||||3|3|3|2|2.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||1|1|1|||||2|2||||4|4||||Red|Amachi|Child: Graduated|128.8||1|1|1|1|F|Black||19|Yes|Mother|28205|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|F|Black||50|28215|Some College|Single|Finance: Banking||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188151|31|0|2|500189677|31|0|2|500037790|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|402864||4|3|45
502136043|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-21|2013-06-06|Followup|2013-02-21|2013-03-13|Complete|Done|4|1|2|2|3|3|2.5|4|1|4|4|3|4|3.33|-24.92|1|3|4|3|3|4|3|3|4|2|1|3|3|2.67|12.36|4|4|4|4|4|4|4|4|0|4|3|4|4|3.75|3|5|5|4|4.25|-11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|4|4|4|3|4|3.5|14.29|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Moved|27.5||1|1|2|2|M|Black||19|No|GrandMother|28227|Other Relative|Unknown||Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500011746|502136472|31|0|1|502459922|1|0|1|500517447|2||-2||4|1|500005291|500005291|-2|500004640|-2|56|1|||7464|9|||1|403321|244354|4|3|45
502222545|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-03|2017-01-24|Followup|2012-08-03|2012-08-06|Complete|Done|3|1|2|1|1|1|1.5|||||||||2|3|3|3|3|3|2.83|||||||||3|3|2|2.67||||||2|4|3|4|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|2|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|77.7||1|1|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|F|White||37|28208|Masters Degree|Single|Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502222979|31|0|2|502196116|1|0|2|500462566|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|403481||4|3|45
502255210|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-27|NaT|Followup|2012-09-27|2012-12-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||77.6||1|1|1|1|M|Black||14|No|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||29|28210|Bachelors Degree|Married|Business: Mgt, Admin|97224|6|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|500910307|31|0|1|502255794|1|0|1|500470233|2||-2||2|1|||-2|500000294|-2|0|10|||7496|10|||1|403500||4|0|45
501796006|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-17|2013-03-21|Followup|2013-02-17|2013-03-05|Complete|Done|4|4|4|3|2|3|3.33|3|4|4|2|3|4|3.33|0|3|4|4|3|2|4|3.33|2|4|4|4|2|4|3.33|0|4|3|4|3.67|4|4|4|4|-8.25|5|5|5|4|4.75||3|3|5|||4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|4|3.67|4|4|3|3.67|0|2|3|2.5|4|2|3|-16.67|2|2|2|2|0|4|4||||Yellow||Volunteer: Time constraint|13.1||3|3|1|1|F|Black||17|No|Mother|28031|Two Parent|Unknown|Y|Yes||School|General Community||Match Support|F|White||37|28031|Masters Degree|Married|Finance: Banking|28202|7|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500015820|501489205|31|0|2|502469185|1|0|2|500595418|2||-2||4|2|||-2||-2|0|4|||7462|13|||1|403791|6008|4|3|45
500186990|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-17|2014-02-28|Followup|2013-02-17|2013-03-18|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|60.4||2|2|3|3|M|Black||19|Yes|Mother|28269|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||51|28269|Bachelors Degree|Married|Unknown|28202|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500188170|31|0|1|500189496|31|0|1|500339895|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|403873||4|1|45
501378357|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-13|NaT|Followup|2013-02-13|2013-04-12|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||97||1|1|2|2|M|Multi-race (Black & White)||18|No|Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Mgt, Admin|28215|10|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501378636|36|0|1|501174997|31|0|1|500339619|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|404239||4|1|45
502824908|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-21|2015-07-22|Followup|2013-02-21|2013-02-20|Complete|Done|3|2|3|1|2|4|2.5|3|2|3|2|3|3|2.67|-6.37|3|4|3|2|3|4|3.17|3|4|4|2|2|3|3|5.67|4|3|2|3|4|4|4|4|-25|4|3|3|4|3.5|5|5|4|4|4.5|-22.22|4|4|4|4|3|4|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|3|4|3.67|4|4|4|4|-8.25|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green||Child: Graduated|41||1|1|1|1|F|Black||19|No|Mother|28226|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community||Match Support|F|White||34|28226|Bachelors Degree|Married|Unknown|29715|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502826191|31|0|2|502891382|1|0|2|500596373|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|404544|399457|4|3|45
501185594|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-29|2016-06-15|Followup|2013-03-01|2013-04-18|Complete|Late|4|4|4|4|4|4|4|||||||||3|4|4|3|4|4|3.67|||||||||4|1|1|2||||||3|1|5|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green||Child: Graduated|99.5||1|1|1|1|M|Multi-race (Black & White)||19|No|Mother|28227|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Consultant|28226|0|8|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501153366|1|0|1|500248756|2||-2||4|1|||-2||-2|0|4|||7452|6|||1|404760||4|3|45
501254255|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-23|2017-02-28|Followup|2012-09-23|2012-09-20|Complete|Done|4|2|2|2|4|3|2.83|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|101.2||1|1|1|1|F|Black||14|No|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28205|Masters Degree|Single|Finance: Banking|28217|0|4|Yahoo!|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501254531|31|0|2|501356688|1|0|2|500282157|2||-2||4|1|||-2|500000294|-2|0|10|||32|2|||1|404894||4|3|45
502551045|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-03-06|Followup|2013-02-22|2013-02-15|Complete|Done|4|1|1|2|1|1|1.67|4|1|1|2|1|4|2.17|-23.04|1|2|3|2|2|2|2|1|1|2|2|1|2|1.5|33.33|3|3|3|3|1|2|2|1.67|79.64|1|3|2|5|2.75|2|2|2|2|2|37.5|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|4|3.86|0|3|4|2|3|3|4|2|3|0|2|3|2.5|2|2|2|25|1|1|1|1|0|4|4|4|4|0|Yellow||Volunteer: Health|24.4||2|2|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||54|28031|Bachelors Degree|Married|Business: Mgt, Admin|28262|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502551498|31|0|2|502864071|1|0|2|500597976|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|404959|401956|4|3|45
502469903|BBBS of Greater Charlotte|Main Office|C|Active|2012-02-22|NaT|Followup|2013-02-22|2013-01-14|Complete|Early|4|4|4|1|3|4|3.33|3|4|4|3|3|4|3.5|-4.86|2|4|4|4|2|4|3.33|3|4|3|3|3|3|3.17|5.05|4|4|4|4|3|4|4|3.67|8.99|3|4|4|4|3.75|4|4|3|3|3.5|7.14|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|2|2|2|2|1|1.5|33.33|2|2|1|1|100|4|4|4|4|0|Green|||60.7||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$15,000 to $19,999|Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||34|28269|Bachelors Degree|Single|Business: Human Resources|28025|2|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500020910|502470350|31|0|1|502868874|31|0|1|500594396|2||-2||2|1|||-2||-2|0|5|||4748|14|1360|3|1|404986|395896|4|3|45
502328599|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-10-31|Followup|2013-02-22|2013-03-06|Complete|Done|3|2|3|2|2|3|2.5|4|1|4|1|4|3|2.83|-11.66|3|4|3|3|3|3|3.17|2|4|4|2|2|4|3|5.67|3|3|3|3|2|2|2|2|50|4|4|4|4|4|4|3|4|5|4|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|2|2.5|2|4|3|-16.67|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Time constraint|32.3||1|1|1|1|M|Black||15|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||73|28226|Bachelors Degree|Widowed|Construction||7|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502329034|31|0|1|502732347|1|0|1|500594124|2||-2||4|3|||-2||-2|0|10|||131|1|||1|405142|376848|4|3|45
502860019|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-02-24|Followup|2013-02-22|2013-01-14|Complete|Early|4|2|1|1|3|3|2.33|3|3|4|3|3|4|3.33|-30.03|2|4|4|2|1|4|2.83|2|4|4|4|3|4|3.5|-19.14|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3|3|3|4|3.25|53.85|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|4|4|4|4|3|3.67|8.99|4|4|4|2|1|1.5|166.67|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Time constraint|24.1||1|1|1|1|F|Hispanic||19|No|Mother|28213|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|White||36|28205|Bachelors Degree||Tech: Engineer|28204|1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502861418|3|0|2|502873149|1|0|2|500596129|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|405323|390412|4|3|45
502002990|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-28|2013-08-29|Baseline|2012-02-23|2012-03-26|Complete|Done|4|4|1|4|4|4|3.5|||||||||1|1|4|4|2|4|2.67|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|4|3.5|||||1|1||||4|4||||Red||Volunteer: Infraction of match rules/agency policies|17.1||1|1|1|1|M|Black||14||Non-Relative: Other|28215|One Parent: Female|$10,000 to $14,999|Y|Yes|AARTF|Neighbor/Friend|General Community||Enrollment|M|Asian||32|28204|Bachelors Degree|Single|Finance: Banking||4|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502003389|31|0|1|502912865|4|0|1|500599902|2||500003586||4|3|||-2||-2|6855|8|||7496|10|||1|405498|-1|4|3|44
502876870|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-06|2013-01-31|Baseline|2012-02-23|2012-03-06|Complete|Done|3|3|4|1|4|4|3.17|||||||||3|4|4|4|1|4|3.33|||||||||4|4|4|4||||||5|3|4|5|4.25|||||||4|4|4|4|2|3|2|3.29||||||||||4|4|3|3.67||||||1|2|1.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|10.9||2|2|1|1|F|Black||16|No|GrandMother|28206|Grandparents|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|White||30|28205|Associate Degree|Single|Business: Mgt, Admin|28204|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502878273|31|0|2|502818822|1|0|2|500599930|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|405521|-1|4|3|44
502893765|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-08|2015-05-11|Baseline|2012-02-23|2012-03-08|Complete|Done|4|4|4|2|3|3|3.33|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|3|3||||||2|2|2|||||1|1||||4|4||||Green||Child: Graduated|38.1||1|1|1|1|F|Black||19|No|Mother|28213|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||32|28262|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502895172|31|0|2|502874079|31|0|2|500599963|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|405542|-1|4|3|44
501525308|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-16|2015-06-18|Followup|2013-02-16|2013-04-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|76||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28205|Some College|Married|Retail: Sales|28206|1|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|501525600|31|0|1|501536144|1|0|1|500335230|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|405606||4|1|45
502526973|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-19|2013-02-21|Baseline|2012-02-23|2012-07-19|Complete|Done|2|4|4|3|3|2|3|||||||||1|1|1|1|2|3|1.5|||||||||4|1|1|2||||||1|2|3|1|1.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|1|2|||||1|1||||4|4||||Green||Volunteer: Moved|7.1||1|1|1|1|M|Hispanic||19|No|Mother|28210|One Parent: Female|Less than $10,000||Yes||Relative|General Community||Match Support|M|Hispanic||27|28202|Bachelors Degree|Single|Finance|28255|0|11|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|502527426|3|0|1|503037794|3|0|1|500623286|2||-2||4|1|||-2||-2|0|3|||7447|3|||1|405610|-1|4|3|44
502926909|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-30|2013-08-15|Baseline|2012-02-27|2012-03-30|Complete|Done|3|2|4|2|3|4|3|||||||||4|4|3|4|4|1|3.33|||||||||4|3|4|3.67||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Red||Volunteer: Moved|16.5||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes|AARTF|BBBS Board/Staff|General Community||Match Support|M|White||42|28205|PHD|Divorced|Education: Teacher||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502928325|31|0|1|502880005|1|0|1|500600626|2||-2||4|3|||-2||-2|7294|13|||7464|9|||1|406712|-1|4|3|44
502875279|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-19|2014-12-17|Baseline|2012-02-27|2012-03-19|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|4|3|4|1|2|2.83|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4||||||||3|2|2.5|||||1|1||||4|4||||Red||Volunteer: Time constraint|33||2|2|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||32|28210|Bachelors Degree|Single|Business: Sales||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502876679|31|0|2|502864263|31|0|2|500600651|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|406736|-1|4|3|44
502506397|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-30|2016-11-01|Baseline|2012-02-28|2012-06-30|Complete|Done|2|1|2|2|3|3|2.17|||||||||3|3|4|3|2|4|3.17|||||||||3|2|2|2.33||||||5|4|3|2|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||1|3|3|2.33||||||2|4|3|||||1|1||||4|4||||Yellow||Child: Severity of challenges|52.1||1|1|1|1|F|White||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||33|28277|Bachelors Degree|Single|Consultant|28202|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502506846|1|0|2|503039829|1|0|2|500619509|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|407242|-1|4|3|44
502142129|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-04|2013-05-22|Baseline|2012-02-28|2012-04-04|Complete|Done|3|1|4|3|2|3|2.67|||||||||3|3|4|4|4|3|3.5|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||3|4|4|3|4|4|2|3.43||||||||||3|3|2|2.67||||||3|2|2.5|||||1|1||||4|4||||Red||Volunteer: Time constraint|13.6||1|1|1|1|F|Some Other Race||19|No|Father|28214|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||45|28209|Bachelors Degree|Single|Tech: Engineer|2494|14|0||Relative|Big|General Community||Match Support|277|60|598|500000170|500015820|502142558|41|0|2|502926748|1|0|2|500605216|2||-2||4|3|||-2||-2|0|10|||0|11|||1|407441|-1|4|3|44
502859604|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-26|2014-12-18|Baseline|2012-02-28|2012-03-26|Complete|Done|3|4|4|3|3|4|3.5|||||||||4|2|4|4|4|3|3.5|||||||||4|4|4|4||||||5|3|5|1|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||1|1||||4|4||||Green||Volunteer: Time constraint|32.8||1|1|1|1|F|Hispanic|Other Central American|19|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Hispanic||40|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502860998|3|14|2|502863229|3|0|2|500604130|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|407511|-1|4|3|44
501833026|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-02|2016-09-30|Followup|2013-03-02|2013-03-22|Complete|Done|4|4|4|2|4|4|3.67|2|4|4|3|1|3|2.83|29.68|2|4|4|2|2|4|3|2|1|3|2|3|2|2.17|38.25|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3|3|3.25|23.08|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|2|3|33.33|3|3|3|2|4|3|0|2|2|1|1|100|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|67||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28205|Masters Degree|Single|Education: Teacher|2122|1|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502451325|1|0|2|500518305|2||-2||4|2|500005291|500005291|-2|500000294|-2|0|10|||7464|9|||1|407901|157601|4|3|45
502057399|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2014-03-31|Followup|2013-02-28|2013-03-07|Declined|Done||||||||4|3|4|3|2|4|3.33|||||||||3|3|2|3|3|3|2.83||||||4|4|4|4|||||||4|5|5|4|4.5||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|1|2.5||||2|2|||||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|37||2|2|1|1|M|White||20|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||50|28078|Bachelors Degree|Single|Arts, Entertainment, Sports|28078|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502057823|1|0|1|502389976|1|0|1|500516780|2||-2||4|2|500005291|500005291|-2||-2|0|4|||7464|9|||1|408303|161076|4|1|45
501635933|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-19|2014-02-26|Baseline|2012-03-01|2012-03-19|Comprehension|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|23.3||1|1|1|1|M|Black||14|No|Mother|28202|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||29|28078|Bachelors Degree|Single|Finance|28205|1|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501636256|31|0|1|502887536|1|0|1|500601528|2||-2||4|3|||-2||-2|0|10|||7438|1|||1|408577|-1|4|2|44
502197486|BBBS of Greater Charlotte|Main Office|C|Active|2012-02-22|NaT|Followup|2013-02-22|2013-02-12|Complete|Done|4|2|1|1|4|3|2.5|||||||||2|4|3|1|2|4|2.67|||||||||4|4|4|4||||||5|3|4|2|3.5|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|3|3.67||||||1|2|1.5|||||2|2||||4|4||||Green|||60.7||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||30|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502197915|31|0|1|502870668|1|0|1|500597982|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|409359||4|3|45
502255223|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-11|NaT|Followup|2012-08-11|2012-08-22|Complete|Done|3|2|4|3|3|3|3|||||||||3|4|4|4|3|3|3.5|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||79.1||1|1|1|1|F|Hispanic||14|No|Mother|28212|One Parent: Female|Unknown|Y|No|Spanish Radio|Media|General Community||Match Support|F|White||33|28209||Single|Education: Teacher||0|0||High School Partner|Big|General Community||Match Support|277|60|598|500000170|500020753|502255655|3|0|2|501823103|1|0|2|500463922|2||-2||2|1|||-2||-2|7068|1|||0|4|||1|409436||4|3|45
502838495|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-24|2012-06-05|Baseline|2012-03-06|2012-04-24|Complete|Done|3|2|3|1|3|3|2.5|||||||||1|2|2|2|2|3|2|||||||||2|2|2|2||||||3|4|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||2|4|1|2.33||||||4|2|3|||||1|1||||4|4||||Green||Volunteer: Unrealistic expectations|1.4||1|1|1|1|F|Hispanic|Other Central American|16|No|Mother|28213|Grandparents|Unknown|Y|Yes||School|General Community||Match Support|F|Hispanic||38|28202||Single|Unknown||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502839787|3|14|2|502707985|3|0|2|500605723|2||-2||4|1|||-2||-2|0|4|||7462|13|||1|410062|-1|4|3|44
502859599|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2014-05-05|Baseline|2012-03-06|2012-04-30|Complete|Done|3|1|2|1|3|4|2.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|4|3.67||||||2|3|2.5|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|24.1||1|1|1|1|M|Hispanic|Other Central American|14|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|Hispanic|Other South American|35|28209|High School Graduate|Married|Business||0|1|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500017777|502860998|3|14|1|502864237|3|15|1|500610310|2||-2||4|1|||-2||-2|0|4|||17161|11|||1|410107|-1|4|3|44
502317496|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-12|2013-06-18|Baseline|2012-03-08|2012-04-12|Complete|Done|4|4|4|2|3|2|3.17|||||||||2|2|3|2|1|3|2.17|||||||||3|2|3|2.67||||||3|5|2|2|3|||||||4|1|4|3|3|4|4|3.29||||||||||3|4|3|3.33||||||1|1|1|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|14.2||1|1|1|1|M|Black||18|Yes|Mother|28214|One Parent: Female|Unknown||Yes||School|General Community|Amachi, Project Big|Match Support|M|Black||42|28214|Some College|Married|Business|28217|17|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502317931|31|0|1|502860968|31|0|1|500602986|2||500004641||4|3||500000294, 500004640|-2||-2|0|4|||7462|13|||1|411006|-1|4|3|44
502893765|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-08|2015-05-11|Followup|2013-03-08|2013-04-01|Complete|Done|3|4|4|4|3|4|3.67|4|4|4|2|3|3|3.33|10.21|2|4|4|4|2|3|3.17|3|3|3|3|3|3|3|5.67|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|2|2|3|3|2.5|30|4|4|4|3|4|4|1|3.43|4|4|4|4|4|4|3|3.86|-11.14|4|4|3|3.67|2|4|3|3|22.33|3|1|2|2|2|2|0|1|1|1|1|0|4|4|4|4|0|Green||Child: Graduated|38.1||1|1|1|1|F|Black||19|No|Mother|28213|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||32|28262|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502895172|31|0|2|502874079|31|0|2|500599963|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|411126|405542|4|3|45
502874566|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-24|2015-10-16|Baseline|2012-03-09|2012-05-24|Complete|Done|3|1|3|1|3|4|2.5|||||||||2|3|4|2|3|4|3|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2|||||||||Green||Volunteer: Moved|40.7||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|White||28|27235|Bachelors Degree||Business: Engineer||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502875969|3|10|2|502894480|1|0|2|500607372|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|411252|-1|4|3|44
501936316|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-28|2016-08-29|Followup|2013-01-28|2013-03-01|Complete|Done|3|2|2|2|3|3|2.5|3|3|3|2|2|2|2.5|0|4|4|3|2|2|3|3|3|3||3|3|3|||4|4|4|4|3|3|3|3|33.33|5|5|3|3|4|4|5|4|4|4.25|-5.88|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|1|1|2|2|-50|4|4||||Green||Child/Family: Lost contact with volunteer/agency|79||1|1|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||54|28203|||Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|501936714|31|0|1|501872326|1|0|1|500428557|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|411330|28181|4|3|45
502896719|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-01|2015-08-19|Baseline|2012-03-09|2012-06-01|Complete|Done|4|1|2|1||4||||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Yellow||Volunteer: Moved|38.6||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|F|White||27|28269|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|502898127|31|0|2|502959645|1|0|2|500614239|2||-2||4|2|||-2||-2|0|10|||46|2|||1|411397|-1|4|3|44
502236255|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-24|2014-11-30|Followup|2013-02-24|2013-02-04|Complete|Early|3|4|2|4|1|1|2.5|||||||||1|4|4|2|1|4|2.67|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|45.2||1|1|1|1|M|Black||14|No|Father|28214|Two Parent|Unknown||Yes||Relative|General Community||Match Support|M|White||64|28207|Masters Degree|Married|Education: Teacher||0|0|Radio|Media|Big|General Site|mentor2.0 2015|Enrollment|277|60|598|500000170|500013781|502236686|31|0|1|502436546|1|0|1|500518376|2||-2||4|3|||-2|500015184|-1|0|3|||131|1|||1|411646||4|3|45
502945480|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-29|NaT|Baseline|2012-03-12|2012-03-29|Complete|Done|1|4|3|1|4|4|2.83|||||||||1|4|3|3|2|2|2.5|||||||||4|4|4|4||||||5|5|3|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||1|3|2|||||2|2||||4|4||||Green|||59.6||1|1|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||54|28262|Bachelors Degree|Single|Business: Mgt, Admin||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502946906|31|0|2|502919780|31|0|2|500603409|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|411819|-1|4|3|44
500824037|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-15|NaT|Followup|2013-03-15|2013-03-11|Complete|Done|4|4|4|3|3|4|3.67|||||||||4|4|4|4|1|4|3.5|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|||120||1|1|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|F|White||34|28210|Bachelors Degree|Single|Education: Teacher|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500824306|31|0|2|500789337|1|0|2|500165956|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|412157||4|3|45
500577150|BBBS of Greater Charlotte|Main Office|C|Active|2011-03-22|NaT|Followup|2013-03-22|2013-03-06|Complete|Early|3|2|4|3|3|3|3|||||||||3|4|3|3|2|3|3|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||3|1|2|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI||71.8||4|5|1|2|F|Black||15||Aunt|28213|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||40|29715|||Customer Service||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500214349|31|0|2|501734288|1|0|2|500526894|2||500004641||2|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|412162||4|3|45
500570756|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-22|2013-02-19|Followup|2013-03-22|2013-02-19|Complete|Early|4|3|4|3|3|4|3.5|||||||||2|3|3|2|3|2|2.5|||||||||4|4|4|4||||||5|1|1|3|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Moved|23||4|5|1|2|F|Black||15||Aunt|28213|Two Parent|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||25|28202|||Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500214349|31|0|2|501865290|1|0|2|500526958|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|412245||4|3|45
502278985|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-01|NaT|Followup|2013-03-01|2013-03-18|Complete|Done|3|4|4|2|2|3|3|||||||||2|3|3|3|3|3|2.83|||||||||4|4|3|3.67||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|2|2.5|||||2|2||||3|3||||Green|Project Big||60.5||1|1|2|2|M|Black||14|No|Mother|28213|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||40|28269||Married|Business: Marketing||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502279417|31|0|1|500220237|31|0|1|500599107|2||-2||2|1|500004640||-2|500000294|-2|6854|8|||2238|7|||1|412566||4|3|45
501833031|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2015-11-04|Followup|2013-02-28|2013-03-22|Complete|Done|4|4|4|1|4|4|3.5|3|3|1|4|4|4|3.17|10.41|1|3|3|2|2|3|2.33|2|2|3|2|4|4|2.83|-17.67|4|4|4|4|4|4|4|4|0|2|2|2|2|2|4|4|4|4|4|-50|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|4|4|4|4|-8.25|1|3|2|4|2|3|-33.33|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Moved|56.2||1|1|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28205|Masters Degree|Single|Medical: Doctor, Provider|28277|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502427342|1|0|2|500518294|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|412627|157600|4|3|45
502681380|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-21|2014-12-18|Baseline|2012-03-14|2012-03-21|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|3|4|1|4|3.33|||||||||3|3|3|3||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||2|3|2.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|32.9||1|1|1|1|M|White||14|No|Mother|28075|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|M|White||29|28277|Bachelors Degree|Single|Insurance|28262|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502682208|1|0|1|502847991|1|0|1|500603939|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|412646|-1|4|3|44
501788776|BBBS of Greater Charlotte|Main Office|C|Active|2010-01-25|NaT|Followup|2013-01-25|2013-03-09|Complete|Done|2|2|2|2|3|2|2.17|||||||||2|2|2|2|2|2|2|||||||||4|2|2|2.67||||||2|3|2|2|2.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|3|3.33||||||2|2|2|||||2|2||||4|4||||Green|Amachi||85.7||1|1|1|1|M|Black||14|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||64|28117||Married|Business: Sales|28031|0|0|Alpha Kappa Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500020752|501789128|31|0|1|501698382|1|0|1|500418170|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||8697|14|||1|412899||4|3|45
500938154|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-12|NaT|Followup|2013-01-12|2013-01-17|Complete|Done|4|3|4|2|4|4|3.5|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||98.1||2|2|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||32|28208|Associate Degree|Single|Service: Restaurant|28211|4|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500938424|31|0|1|501446421|1|0|1|500323753|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|412905||4|3|45
502275241|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-21|2015-10-15|Followup|2013-03-21|2013-03-13|Complete|Done|3|3|4|3|3|3|3.17|4|3|3|3|4|3|3.33|-4.8|3|3|3|2|4|3|3|3|3|4|3|3|2|3|0|4|4|4|4|4|4|4|4|0|3|3|2|2|2.5|2|3|3|3|2.75|-9.09|4|4|4|4|3|4|3|3.71|4|4|4|4|4|||||3|4|3|3.33|3|3|3|3|11|4|2|3|3|3|3|0|2|2|2|2|0|4|4||||Green|Amachi|Child: Lost interest|54.8||1|1|1|1|F|Black||17|No|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||26|28031|Bachelors Degree|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|502275673|31|0|2|502394690|1|0|2|500521625|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7496|10|||1|413244|235273|4|3|45
502850780|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-06|2013-04-26|Baseline|2012-03-19|2012-04-06|Complete|Done|3|3|4|4|4|4|3.67|||||||||2|3|3|1|4|3|2.67|||||||||4|3|3|3.33||||||3|3|3|5|3.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|2|3.33||||||3|2|2.5|||||1|1||||4|4||||Red||Child/Family: Moved|12.6||1|1|1|1|M|Black||16|No|Mother|28105|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community||Match Support|M|White||54|28173|Some College|Married|Unemployed||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|502852142|31|0|1|502835253|1|0|1|500604783|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|414074|-1|4|3|44
502875279|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-19|2014-12-17|Followup|2013-03-19|2013-03-15|Complete|Done|3|4|4|1|4|4|3.33|3|2|2|2|3|3|2.5|33.2|4|4|4|4|1|4|3.5|3|4|3|4|1|2|2.83|23.67|4|4|4|4|4|4|4|4|0|5|4|4|5|4.5|3|3|4|5|3.75|20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4||||3|2|2.5|3|2|2.5|0|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Time constraint|33||2|2|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||32|28210|Bachelors Degree|Single|Business: Sales||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502876679|31|0|2|502864263|31|0|2|500600651|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|414115|406736|4|3|45
501635933|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-19|2014-02-26|Followup|2013-03-19|2013-04-12|Complete|Done|3|1|4|1|1|1|1.83|||||||||1|4|4|2|2|3|2.67|||||||||4|4|4|4||||||3|2|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Red||Volunteer: Time constraint|23.3||1|1|1|1|M|Black||14|No|Mother|28202|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||29|28078|Bachelors Degree|Single|Finance|28205|1|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501636256|31|0|1|502887536|1|0|1|500601528|2||-2||4|3|||-2||-2|0|10|||7438|1|||1|414169|408577|4|3|45
502671420|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-13|2013-04-04|Baseline|2012-03-19|2012-04-13|Complete|Done|3|4|3|2|3|3|3|||||||||4|3|3|3|3|4|3.33|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|4|3|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|11.7||1|1|1|1|M|Black||17|No|Mother|28210|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Multi-race (Black & White)||33|28277|Associate Degree|Married|Tech: Computer/Programmer||6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502672248|31|0|1|502938924|36|0|1|500604987|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|414321|-1|4|3|44
502183053|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-28|NaT|Baseline|2012-03-20|2012-06-28|Complete|Done|3|1|2|1|1|2|1.67|||||||||4|2|4|2|3|4|3.17|||||||||4|4|3|3.67||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|||56.6||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||46|28134|Bachelors Degree|Married|Finance|28105|1|6|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|502183482|31|0|1|503073638|31|0|1|500621039|2||-2||2|1|||-2|500014681|-2|0|10|||4748|14|633|1|1|414734|-1|4|3|44
502681380|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-21|2014-12-18|Followup|2013-03-21|2013-04-04|Complete|Done|3|3|3|2|3|4|3|3|4|4|4|3|4|3.67|-18.26|4|4|4|3|3|4|3.67|4|4|3|4|1|4|3.33|10.21|4|4|3|3.67|3|3|3|3|22.33|5|4|4|5|4.5|4|4|5|5|4.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|2|3|33.33|4|4|4|2|3|2.5|60|1|1|2|2|-50|4|4|4|4|0|Green||Volunteer: Lost contact with child/agency|32.9||1|1|1|1|M|White||14|No|Mother|28075|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|M|White||29|28277|Bachelors Degree|Single|Insurance|28262|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502682208|1|0|1|502847991|1|0|1|500603939|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|414962|412646|4|3|45
502700503|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-30|NaT|Baseline|2012-03-22|2012-03-30|Complete|Done|4|1|1|1|3|1|1.83|||||||||2|3|3|2|2|2|2.33|||||||||4|4|4|4||||||3|2|2|3|2.5|||||||4|4|4|4||4|3|||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||59.5||1|1|1|1|M|Black||14|No|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||36|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502701348|31|0|1|502931327|1|0|1|500605634|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|415426|-1|4|3|44
502926905|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-31|2014-09-18|Baseline|2012-03-22|2012-10-31|Complete|Done|2|4|4|4|4|4|3.67|||||||||2|3|3|2|2|3|2.5|||||||||4|3|3|3.33||||||2|3|3|2|2.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||3|4|3.5|||||2|2||||4|4||||Yellow||Volunteer: Feels incompatible with child/family|22.6||1|1|1|1|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||32|28216|Bachelors Degree|Single|Tech: Support, Writing|28117|1|9|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502928325|31|0|2|503096831|31|0|2|500635818|2||-2||4|2|||-2||-2|7294|13|||7438|1|||1|415449|-1|4|3|44
502874571|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-27|2013-07-29|Baseline|2012-03-22|2012-06-27|Complete|Done|3|2|3|2|2|4|2.67|||||||||2|4|3|3|4|3|3.17|||||||||4|4|4|4||||||5||4|3||||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||1|1||||4|4||||Red||Volunteer: Moved|13||1|1|2|2|F|Hispanic||17|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|F|White||30|28202|Bachelors Degree|Single|Tech: Management|28202|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|502875969|3|0|2|501375210|1|0|2|500617142|2||-2||4|3|||-2||-2|0|4|||7446|3|||1|415556|-1|4|3|44
502912141|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-05|2016-06-17|Baseline|2012-03-23|2012-04-05|Complete|Done|2|4|4|3|4|4|3.5|||||||||2|4|3|2|2|4|2.83|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4||3|||||||4|||||||1|1||||4|4||||Red||Volunteer: Moved|50.4||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Business: Marketing|28203|0|8|Other Church Partner|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|502913549|31|0|2|502932948|1|0|2|500605880|2||-2||4|3|||-2||-2|34|2|||7453|7|||1|415863|-1|4|3|44
502320003|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2014-09-24|Baseline|2012-03-26|2012-04-30|Complete|Done|4|2|4|4|3|4|3.5|||||||||2|3|4|1|2|4|2.67|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|1|2.5|||||2|2||||4|4||||Red||Volunteer: Moved|28.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||30|28216||Single|Tech: Research/Design||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502320438|31|0|2|502810883|31|0|2|500606071|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|416362|-1|4|3|44
502610186|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-26|NaT|Followup|2013-03-26|2013-03-24|Complete|Done|4|4|4|1|3|4|3.33|4|1|4|1|4|4|3|11|2|4|4|2|2|4|3|3|3|3|2|2|3|2.67|12.36|4|3|4|3.67|4|4|4|4|-8.25|4|3|4|3|3.5|2|4|2|4|3|16.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|3|3|3|33.33|2|2|2|3|3|3|-33.33|2|2|2|2|0|4|4|4|4|0|Green|||59.7||1|1|1|1|F|Black||16|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Asian||35|28210|Masters Degree|Married|Arts, Entertainment, Sports|28202|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|502610737|31|0|2|502913393|4|0|2|500601697|2||-2||2|1|||-2||-2|6854|8|||7671|13|||1|416418|388768|4|3|45
502859604|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-26|2014-12-18|Followup|2013-03-26|2013-04-12|Complete|Done|4|2|2|2|3|3|2.67|3|4|4|3|3|4|3.5|-23.71|2|4|4|2|2|3|2.83|4|2|4|4|4|3|3.5|-19.14|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|3|5|1|3.5|42.86|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|4|4|4|3|3|3|33.33|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Time constraint|32.8||1|1|1|1|F|Hispanic|Other Central American|19|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Hispanic||40|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502860998|3|14|2|502863229|3|0|2|500604130|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|416496|407511|4|3|45
502902269|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-26|2014-02-21|Baseline|2012-03-27|2013-01-26|Complete|Done|4|3|4|1|3|4|3.17|||||||||2|3|4|3|4|4|3.33|||||||||4|4|4|4||||||3|5|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child: Lost interest|12.8||1|1|3|3|M|Black||14|No|Mother|28215|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Enrollment|M|Black||31|28203|Juris Doctorate (JD)||Law: Lawyer|28203|1|0|Self|Self|Big|General Site|mentor2.0 2015|Match Support|277|60|598|500000170|500011349|502903679|31|0|1|501631588|31|0|1|500677452|2||-2||4|2|||-2|500015184|-1|0|10|||7464|9|||1|417037|-1|4|3|44
502431164|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-30|2015-10-12|Baseline|2012-03-27|2012-03-30|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|4|4|2|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Graduated|42.4||1|1|1|1|M|Black||19|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community||Match Support|M|White||59|28277|Masters Degree|Single|Tech: Computer/Programmer|28203|3|4|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502431607|31|0|1|502850528|1|0|1|500606503|2||-2||4|1|||-2||-2|0|5|||7439|1|||1|417125|-1|4|3|44
502002990|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-28|2013-08-29|Followup|2013-03-28|2013-04-02|Complete|Done|3|3|4|2|4|3|3.17|4|4|1|4|4|4|3.5|-9.43|2|3|3|2|2|3|2.5|1|1|4|4|2|4|2.67|-6.37|4|4|4|4|4|4|4|4|0|3|4|5|4|4|3|5|5|5|4.5|-11.11|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|4|3|3.33|0|2|2|2|3|4|3.5|-42.86|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Infraction of match rules/agency policies|17.1||1|1|1|1|M|Black||14||Non-Relative: Other|28215|One Parent: Female|$10,000 to $14,999|Y|Yes|AARTF|Neighbor/Friend|General Community||Enrollment|M|Asian||32|28204|Bachelors Degree|Single|Finance: Banking||4|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502003389|31|0|1|502912865|4|0|1|500599902|2||500003586||4|3|||-2||-2|6855|8|||7496|10|||1|417708|405498|4|3|45
502526965|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-03|NaT|Baseline|2012-03-28|2012-04-03|Complete|Done|4|3|3|4|4|4|3.67|||||||||2|4|2|3|2|3|2.67|||||||||4|4|4|4||||||3|4|3|5|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||59.4||1|1|1|1|M|Black||17|No|Mother|28278|Two Mothers|$50,000 to $59,999||No||Self|General Community||Match Support|M|White||32|28278|Bachelors Degree|Single|Medical|28208|3|5|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502527418|31|0|1|502881104|1|0|1|500606886|2||-2||2|1|||-2||-2|0|10|||17161|11|||1|417778|-1|4|3|44
502845758|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-19|2015-09-16|Baseline|2012-03-28|2012-04-19|Complete|Done|4|2|4|2|3|4|3.17|||||||||1|3|3|2|2|4|2.5|||||||||4|3|3|3.33||||||3|4|4|2|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|40.9||1|1|1|1|M|Black||15|No|Mother|28202|One Parent: Male|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28277||Single|Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502847118|31|0|1|502944923|1|0|1|500606912|2||-2||4|3|||-2||-2|34|2|||7464|9|||1|417837|-1|4|3|44
500948129|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-18|2016-06-30|Followup|2013-03-18|2013-03-17|Complete|Done|3|3|3|4|3|3|3.17|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|75.4||2|2|1|1|F|Black||18|No|Mother|28217|One Parent: Female|$25,000 to $29,999|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||40|28203|Some College|Living w/ Significant Other|Finance: Banking|28281|1|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501891556|1|0|2|500438403|2||500003586||4|1|500000294|500000294|-2||-2|34|2|||7464|9|||1|418045||4|3|45
500843863|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-21|2016-06-17|Followup|2013-02-21|2013-02-05|Complete|Early|3|4|4|4|4|3|3.67|||||||||2|3|4|2|2|3|2.67|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|1|2|||||2|2||||4|4||||Green|Amachi|Volunteer: Changed workplace/school partnership|99.8||2|2|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|No|TV|Media|General Community|Amachi|Match Support|F|Black||32|28269|Bachelors Degree|Single|Business: Marketing|28273|0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500844129|31|0|2|501078655|31|0|2|500241388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|56|1|||2238|7|||1|418046||4|3|45
502945480|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-29|NaT|Followup|2013-03-29|2013-03-26|Complete|Done|4|4|4|1|4|4|3.5|1|4|3|1|4|4|2.83|23.67|2|3|3|1|4|3|2.67|1|4|3|3|2|2|2.5|6.8|4|4|4|4|4|4|4|4|0|4|5|3|5|4.25|5|5|3|4|4.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|1|2.33|4|4|3|3.67|-36.51|3|3|3|1|3|2|50|2|2|2|2|0|4|4|4|4|0|Green|||59.6||1|1|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||54|28262|Bachelors Degree|Single|Business: Mgt, Admin||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502946906|31|0|2|502919780|31|0|2|500603409|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|418231|411819|4|3|45
502765606|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-03|2014-09-24|Baseline|2012-03-29|2012-04-03|Complete|Done|4|1|2|2|2|4|2.5|||||||||3|2|3|2|2|2|2.33|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||3|4|3|4|2|4|4|3.43||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Red||Volunteer: Moved|29.7||1|1|1|1|F|Black||19|No|Mother|28105|One Parent: Female|$15,000 to $19,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28209|Some College|Single|Finance: Accountant|28232|0|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502766519|31|0|2|502842142|31|0|2|500607132|2||-2||4|3|||-2||-2|6854|8|||7462|13|||1|418328|-1|4|3|44
500896361|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-14|2014-02-27|Followup|2013-01-14|2013-01-07|Complete|Done|3|4|4|4|4|3|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||1|1|1|1||||||4|4|4|||||2|2||||4|4||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|61.4||2|2|1|1|F|Black||20|Yes|Mother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28075||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500012459|500896631|31|0|2|501276501|31|0|2|500291021|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|418574||4|3|45
502926909|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-30|2013-08-15|Followup|2013-03-30|2013-03-20|Complete|Done|3|4|4|1|4|4|3.33|3|2|4|2|3|4|3|11|4|4|4|4|4|4|4|4|4|3|4|4|1|3.33|20.12|4|4|4|4|4|3|4|3.67|8.99|3|4|3|5|3.75|5|5|4|5|4.75|-21.05|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|3|2.5|4|2|3|-16.67|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Moved|16.5||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes|AARTF|BBBS Board/Staff|General Community||Match Support|M|White||42|28205|PHD|Divorced|Education: Teacher||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502928325|31|0|1|502880005|1|0|1|500600626|2||-2||4|3|||-2||-2|7294|13|||7464|9|||1|418615|406712|4|3|45
501295538|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-30|NaT|Followup|2013-03-30|2013-02-20|Complete|Early|4|3|3|4|3|3|3.33|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||59.5||2|2|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||31|28078|Bachelors Degree||Medical||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500740560|31|0|2|502897530|1|0|2|500603727|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|418627||4|3|45
502700503|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-30|NaT|Followup|2013-03-30|2013-03-27|Complete|Done|3|1|4|2|4|3|2.83|4|1|1|1|3|1|1.83|54.64|2|4|4|2|4|4|3.33|2|3|3|2|2|2|2.33|42.92|4|4|4|4|4|4|4|4|0|3|3|4|5|3.75|3|2|2|3|2.5|50|4|4|4|4|4|4|4|4|4|4|4|4||4|3|||4|4|4|4|4|4|4|4|0|4|1|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Green|||59.5||1|1|1|1|M|Black||14|No|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||36|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502701348|31|0|1|502931327|1|0|1|500605634|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|418635|415426|4|3|45
500185863|BBBS of Greater Charlotte|Main Office|C|Completed|2005-03-12|2014-05-15|Followup|2013-03-12|2013-04-24|Complete|Done|4|1|2|1|1|3|2|||||||||4|3|3|2|3|4|3.17|||||||||4|4|4|4||||||3|4|5|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|110.1||1|1|1|1|F|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||43|28202|Bachelors Degree|Married|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187435|31|0|2|500188915|1|0|2|500036915|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|418713||4|3|45
502431164|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-30|2015-10-12|Followup|2013-03-30|2013-04-10|Complete|Done|2|3|2|1|1|4|2.17|4|4|4|3|4|4|3.83|-43.34|4|3|3|4|2|4|3.33|4|4|4|4|4|4|4|-16.75|4|4|4|4|4|4|4|4|0|4|3|2|4|3.25|3|4|4|2|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|4|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Green||Child: Graduated|42.4||1|1|1|1|M|Black||19|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community||Match Support|M|White||59|28277|Masters Degree|Single|Tech: Computer/Programmer|28203|3|4|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502431607|31|0|1|502850528|1|0|1|500606503|2||-2||4|1|||-2||-2|0|5|||7439|1|||1|418717|417125|4|3|45
500186206|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-24|2013-09-30|Followup|2013-02-24|2013-04-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Moved|103.2||1|1|1|1|M|Black||20||GrandMother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||44|28214|PHD|Married|Medical: Doctor, Provider||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|500187812|31|0|1|500189157|31|0|1|500037157|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|418719||4|1|45
502866475|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-23|NaT|Baseline|2012-03-30|2012-05-23|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|2|4|4|3.5|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Green|||57.8||1|1|1|1|M|Black||16|No|Mother|28270|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|M|White||29|28203|Bachelors Degree||Finance: Accountant||1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502867876|31|0|1|502961396|1|0|1|500614954|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|418831|-1|4|3|44
502319984|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-03-24|Baseline|2012-03-30|2012-04-30|Complete|Done|3|3|4|4|4|4|3.67|||||||||2|4|3|2|2|4|2.83|||||||||4|4|4|4||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Red||Volunteer: Time constraint|34.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Bachelors Degree|Single|Finance|28216|3|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502320419|31|0|1|502290677|1|0|1|500607367|2||-2||4|3||500005291|-2||-2|6854|8|||17161|11|||1|418895|-1|4|3|44
502319972|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-08-19|Baseline|2012-03-30|2012-04-30|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow||Volunteer: Moved|39.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Less than $10,000||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||32|28214|Bachelors Degree|Married|Self-Employed, Entrepreneur|29715|0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502320407|31|0|1|502911091|1|0|1|500607368|2||-2||4|2||500005291|-2||-2|6854|8|||7464|9|||1|418896|-1|4|3|44
500892914|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-16|2014-09-11|Followup|2013-02-16|2013-02-18|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|3|3|2|2|3|2.5|||||||||4|1|3|2.67||||||3|3|4|2|3|||||||3|4|4|4|3|4|4|3.71||||||||||4|4|4|4||||||3|1|2|||||1|1||||4|4||||Red|Amachi|Child: Graduated|54.8||2|2|1|1|M|Black||20|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Sales|28269|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500893173|31|0|1|501964388|1|0|1|500429157|2||500003586||4|3|500000294|500000294|-2||-2|0|5|||7464|9|||1|419037||4|3|45
502828137|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-06-29|Baseline|2012-04-01|2012-04-30|Complete|Done|3|1|1|3|1|1|1.67|||||||||1|2|2|2|1|3|1.83|||||||||4|4|4|4||||||2|2|4|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child/Family: Moved|37.9||1|1|1|1|F|Multi-Race (None of the above)||16|No|Father|28214|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher|28078|0|8|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502829415|7|0|2|502446364|31|0|2|500607445|2||-2||4|1|||-2|500004640|-2|0|10|||7464|9|||1|419338|-1|4|3|44
502828131|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-03-31|Baseline|2012-04-01|2012-04-30|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|4|3|3|4|3|3.17|||||||||4|4|4|4||||||4|5|4|2|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|3|1|2.67||||||3|3|3|||||1|1||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|35||1|1|1|1|F|Multi-Race (None of the above)||17|No|Father|28214|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|White||33|28216|Bachelors Degree|Single|Business: Sales|28270|2|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502829415|7|0|2|502881454|1|0|2|500607446|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|419339|-1|4|3|44
502868925|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-25|2014-09-24|Baseline|2012-04-02|2012-04-25|Complete|Done|3|1|2|1|3|3|2.17|||||||||2|4|4|1|2|3|2.67|||||||||4|3|3|3.33||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|29||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||35|28262|Bachelors Degree|Divorced|Finance: Banking||2|6|Charlotte Cares|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502870324|31|0|2|502885744|31|0|2|500607510|2||-2||4|3|||-2||-2|0|4|||11246|6|||1|419518|-1|4|3|44
502030263|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2013-03-31|2013-04-12|Complete|Done|4|1|2|2|3|3|2.5|||||||||3|3|4|2|2|4|3|||||||||4|4|4|4||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||83.5||1|1|1|1|M|White||15|No|Mother|29710|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community||Match Support|M|White||38|28210|||Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502030662|1|0|1|501923553|1|0|1|500438867|2||-2||2|1|||-2||-2|6855|8|||7464|9|||1|419539||4|3|45
502828146|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2014-05-30|Baseline|2012-04-02|2012-04-30|Complete|Done|2|2|3|2|2|1|2|||||||||2|2|3|2|2|2|2.17|||||||||4|4|4|4||||||2|2|3|2|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|25||1|1|1|1|M|Black||17|No|Father|28214|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|Black||37|28278|Bachelors Degree|Single|Unknown||0|0|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502829415|31|0|1|502860825|31|0|1|500607619|2||-2||4|3|||-2||-2|0|10|||9229|13|||1|419662|-1|4|3|44
502765606|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-03|2014-09-24|Followup|2013-04-03|2013-05-14|Complete|Done|3|2|3|2|3|3|2.67|4|1|2|2|2|4|2.5|6.8|2|3|3|3|3|3|2.83|3|2|3|2|2|2|2.33|21.46|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|3|4|3|3.25|-7.69|3|4|3|4|3|4|4|3.57|3|4|3|4|2|4|4|3.43|4.08|4|4|3|3.67|3|4|4|3.67|0|2|3|2.5|3|2|2.5|0|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Moved|29.7||1|1|1|1|F|Black||19|No|Mother|28105|One Parent: Female|$15,000 to $19,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28209|Some College|Single|Finance: Accountant|28232|0|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502766519|31|0|2|502842142|31|0|2|500607132|2||-2||4|3|||-2||-2|6854|8|||7462|13|||1|419820|418328|4|3|45
502526965|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-03|NaT|Followup|2013-04-03|2013-05-14|Complete|Done|4|3|4|2|4|4|3.5|4|3|3|4|4|4|3.67|-4.63|4|4|3|4|4|4|3.83|2|4|2|3|2|3|2.67|43.45|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|3|5|3.75|6.67|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|3|3.67|4|4|3|3.67|0|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green|||59.4||1|1|1|1|M|Black||17|No|Mother|28278|Two Mothers|$50,000 to $59,999||No||Self|General Community||Match Support|M|White||32|28278|Bachelors Degree|Single|Medical|28208|3|5|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502527418|31|0|1|502881104|1|0|1|500606886|2||-2||2|1|||-2||-2|0|10|||17161|11|||1|420185|417778|4|3|45
502083450|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-05|2013-10-16|Followup|2013-04-05|2013-06-20|Expired|Late||||||||4|4|4|4|3|4|3.83|||||||||4|2|3|2|4|3|3||||||4|4|4|4|||||||3|4|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Yellow||Volunteer: Time constraint|18.4||2|2|3|3|M|Black||16|No|Mother|28027|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||49|28027|Bachelors Degree|Married|Transport: Driver|28208|6|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|277|60|598|500000170|500002335|502083874|31|0|1|500863980|31|0|1|500605881|2||-2||4|2||500005291|-2|500014505, 500014506|-1|7016|11|||7671|13|||1|420797|39542|4|0|45
502941572|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-16|2013-04-22|Baseline|2012-04-05|2012-04-16|Complete|Done|4|2|2|1|3|3|2.5|||||||||2|3|3|3|2|3|2.67|||||||||3|3|3|3||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|Amachi|Child/Family: Moved|12.2||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community|Amachi|Match Support|F|White||44|28269|PHD|Single|Medical|64506|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502942998|31|0|2|502884011|1|0|2|500608269|2||-2||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|420804|-1|4|3|44
502710796|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-13|NaT|Baseline|2012-04-05|2012-04-13|Complete|Done|4|1|2|1|4|4|2.67|||||||||1|1|3|1|1|4|1.83|||||||||3|4|3|3.33||||||3|4|4|2|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2||||4|4||||Green|Project Big||59.1||1|1|1|1|M|Black||17|No|GrandMother|28208|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|Project Big|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502711683|31|0|1|502926804|1|0|1|500608316|2||500004641||2|1|500004640|500004640|-2||-2|6854|8|||7464|9|||1|420876|-1|4|3|44
502912141|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-05|2016-06-17|Followup|2013-04-05|2013-04-01|Complete|Done|3|4|4|4|4|4|3.83|2|4|4|3|4|4|3.5|9.43|4|4|4|4|2|4|3.67|2|4|3|2|2|4|2.83|29.68|4|4|4|4|4|4|4|4|0|5|5|5|4|4.75|3|4|5|5|4.25|11.76|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|4|4|4||3|||3|3|3|4||||1|1|1|1|0|4|4|4|4|0|Red||Volunteer: Moved|50.4||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Business: Marketing|28203|0|8|Other Church Partner|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|502913549|31|0|2|502932948|1|0|2|500605880|2||-2||4|3|||-2||-2|34|2|||7453|7|||1|420990|415863|4|3|45
502809446|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-12|2016-06-20|Baseline|2012-04-05|2012-04-12|Complete|Done|4|4|4|4|3|4|3.83|||||||||2|4|4|3|4|4|3.5|||||||||3|4|4|3.67||||||4|3|5|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|2|3.33||||||4|4|4|||||1|1||||4|4||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|50.3||1|1|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Multi-race (Black & White)||33|28269|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502810724|31|0|2|502909383|36|0|2|500608444|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7462|13|||1|421044|-1|4|3|44
502850780|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-06|2013-04-26|Followup|2013-04-06|2013-04-12|Declined|Done||||||||3|3|4|4|4|4|3.67|||||||||2|3|3|1|4|3|2.67||||||4|3|3|3.33|||||||3|3|3|5|3.5||||||||||4|4|4|4|4|4|2|3.71||||||4|4|2|3.33|||||3|2|2.5||||1|1||||4|4||Red||Child/Family: Moved|12.6||1|1|1|1|M|Black||16|No|Mother|28105|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community||Match Support|M|White||54|28173|Some College|Married|Unemployed||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|502852142|31|0|1|502835253|1|0|1|500604783|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|421218|414074|4|1|45
501011735|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-11|2015-03-05|Followup|2013-04-11|2013-04-01|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|3|4|3|3.5|||||||||4|4|4|4||||||5|3|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Yellow|2010-2012 OJJDP JJI|Child: Lost interest|46.8||3|3|1|1|F|Black||17||Mother|28215|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28215|High School Graduate|Married|Finance: Banking|28255|13|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500012459|500417756|31|0|2|502473442|31|0|2|500528270|2||-2||4|2|500005291|500005291|-2||-2|0|10|||7446|3|||1|421619||4|3|45
502931305|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-27|2012-07-31|Baseline|2012-04-09|2012-04-27|Complete|Done|3|3|4|2|4|4|3.33|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|4|3|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Family structure changed|3.1||1|1|2|2|M|Black||16|No|Mother|28214|One Parent: Female|$100,000 to $124,999||No||Self|General Community||Match Support|M|White||31|28269|Masters Degree|Single|Insurance|28262|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008629|502932726|31|0|1|502500246|1|0|1|500608719|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|421713|-1|4|3|44
501252806|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-25|NaT|Followup|2012-11-25|2013-01-09|Complete|Done|4|3|3|3|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||99.6||1|1|1|1|M|Black||13|No|Mother|28078|One Parent: Female|Unknown||No||Relative|General Community||Match Support|M|Black||45|28262|Bachelors Degree|Married|Business: Mgt, Admin||0|6|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|501253082|31|0|1|501320197|31|0|1|500310204|2||-2||2|1|||-2||-2|0|3|||6247|12|||1|422040||4|3|45
500887862|BBBS of Greater Charlotte|Main Office|C|Active|2011-04-13|NaT|Followup|2013-04-13|2013-04-08|Complete|Done|4|4|4|4|4|3|3.83|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|3|4|5|4.25|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Cabarrus County||71.1||2|2|2|2|F|Black||18|Yes|Mother|28025|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|F|Black||43|28027||Divorced|Finance: Banking||0|7|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500888132|31|0|2|500923430|31|0|2|500530980|2||500016307||2|1|500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|422576||4|3|45
502902247|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-11|NaT|Baseline|2012-04-11|2012-07-11|Complete|Done|2|4|4|2||2||||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||1|1||||4|4||||Green|||56.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||30|28203|Bachelors Degree|Single|Business: Marketing|28117|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502903657|31|0|2|502801082|1|0|2|500619356|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|422744|-1|4|3|44
502846423|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-07|2013-02-28|Baseline|2012-04-11|2012-05-07|Complete|Done|2|4|4|4|4|4|3.67|||||||||3|4|4|2|2|4|3.17|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|9.8||1|1|1|1|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Some Other Race||40|28205|Bachelors Degree|Married|Construction|28031|8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|502847784|31|0|2|502877894|41|0|2|500609448|2||-2||4|2|||-2||-2|0|4|||7496|10|||1|422860|-1|4|3|44
502539860|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-15|2014-02-10|Followup|2013-04-15|2013-04-30|Complete|Done|3|2|2|1|4|3|2.5|3|2|1|1|1|4|2|25|4|3|1|3|3|4|3|2|3|3|3|2|3|2.67|12.36|4|4|4|4|2|2|2|2|100|4|4|5|5|4.5|3|2|1|1|1.75|157.14|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|3|3.33|20.12|4|4|4|||||2|2|1|1|100|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|33.9||1|1|1|1|M|Hispanic||17|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Hispanic||33|28270|Associate Degree|Married|Business: Sales||9|0|Other|BBBS Board/Staff|Big|General Community|Project Big|Match Support|277|60|598|500000170|500017777|502540313|3|0|1|502498837|3|0|1|500529729|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||7671|13|||1|422872|264531|4|3|45
502966254|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-04|2015-03-18|Baseline|2012-04-12|2012-05-04|Complete|Done|2|3|2|4|2|3|2.67|||||||||2|4|3|2|2|3|2.67|||||||||4|3|4|3.67||||||3|4|2|2|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|34.4||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community||Match Support|F|Black||48|28217|Bachelors Degree|Divorced|Medical: Admin|28232|11|5|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|500784955|31|0|2|502895517|31|0|2|500609631|2||-2||4|2|||-2||-2|0|10|||7438|1|||1|423139|-1|4|3|44
501376745|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-01|2016-01-11|Followup|2013-04-01|2013-04-04|Complete|Done|4|2|4|2|3|3|3|||||||||3|4|4|4|3|3|3.5|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green||Volunteer: Time constraint|81.3||1|1|3|4|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28269|||Business: Marketing||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|501377024|31|0|2|500725077|31|0|2|500350905|2||-2||4|1|||-2||-2|6854|8|||46|2|||1|423249||4|3|45
502317496|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-12|2013-06-18|Followup|2013-04-12|2013-06-17|Declined|Late||||||||4|4|4|2|3|2|3.17|||||||||2|2|3|2|1|3|2.17||||||3|2|3|2.67|||||||3|5|2|2|3||||||||||4|1|4|3|3|4|4|3.29||||||3|4|3|3.33|||||1|1|1||||2|2||||4|4||Red||Volunteer: Lost contact with child/agency|14.2||1|1|1|1|M|Black||18|Yes|Mother|28214|One Parent: Female|Unknown||Yes||School|General Community|Amachi, Project Big|Match Support|M|Black||42|28214|Some College|Married|Business|28217|17|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502317931|31|0|1|502860968|31|0|1|500602986|2||500004641||4|3||500000294, 500004640|-2||-2|0|4|||7462|13|||1|423259|411006|4|1|45
502809446|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-12|2016-06-20|Followup|2013-04-12|2013-05-14|Complete|Done|4|4|4|4|4|4|4|4|4|4|4|3|4|3.83|4.44|4|4|4|4|4|4|4|2|4|4|3|4|4|3.5|14.29|4|4|4|4|3|4|4|3.67|8.99|4|5|5|4|4.5|4|3|5|4|4|12.5|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|3|3.71|4.04|4|4|3|3.67|4|4|2|3.33|10.21|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|50.3||1|1|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Multi-race (Black & White)||33|28269|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502810724|31|0|2|502909383|36|0|2|500608444|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7462|13|||1|423300|421044|4|3|45
501340097|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-23|2016-09-19|Followup|2013-03-23|2013-03-20|Complete|Done|3|4|4|2|4|3|3.33|||||||||2|4|3|1|4|3|2.83|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|2|2.67||||||2|1|1.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|77.9||2|2|1|1|M|Multi-race (Black & Hispanic)||17|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Hispanic||28|28277|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340376|38|0|1|501934966|3|0|1|500440292|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|423512||4|3|45
500997880|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-19|2016-07-29|Followup|2013-02-19|2013-03-04|Complete|Done|3|4|4|4|3|4|3.67|||||||||2|4|3|4|2|3|3|||||||||4|3|4|3.67||||||3|5|3|3|3.5|||||||3|3|4|4|4|3|3|3.43||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green||Child: Graduated|101.3||1|1|1|1|M|Black||18|No|Mother|28204|Two Parent|$40,000 to $44,999||Yes||Self|General Community||Match Support|M|White||33|28202|Bachelors Degree|Married|Business: Marketing||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500998153|31|0|1|500990660|1|0|1|500237316|2||-2||4|1|||-2||-2|0|10|||46|2|||1|423627||4|3|45
502710796|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-13|NaT|Followup|2013-04-13|2013-05-14|Complete|Done|4|3|4|3|4|4|3.67|4|1|2|1|4|4|2.67|37.45|3|4|3|4|3|4|3.5|1|1|3|1|1|4|1.83|91.26|4|4|4|4|3|4|3|3.33|20.12|3|4|4|3|3.5|3|4|4|2|3.25|7.69|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|3|3.67|0|2|3|2.5|1|4|2.5|0|2|2|2|2|0|4|4|4|4|0|Green|Project Big||59.1||1|1|1|1|M|Black||17|No|GrandMother|28208|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|Project Big|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502711683|31|0|1|502926804|1|0|1|500608316|2||500004641||2|1|500004640|500004640|-2||-2|6854|8|||7464|9|||1|423643|420876|4|3|45
500961015|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-11|2014-10-02|Followup|2013-04-11|2013-04-03|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|4|3|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|77.7||1|1|1|1|M|Black||20|Yes|Mother|28227|Two Parent|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||43|28104||Married|Tech: Computer/Programmer|29607|10|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500013781|500934638|31|0|1|501210561|31|0|1|500257073|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||17161|11|||1|424090||4|3|45
500546821|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-21|2015-09-15|Followup|2013-02-21|2013-01-09|Complete|Early|4|4|4|4|4|4|4|||||||||2|4|4|2|4|3|3.17|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Child: Graduated|102.8||1|1|3|3|M|Black||20|No|Mother|28083|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||52|28025||Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500012459|500547073|31|0|1|500790181|31|0|1|500159910|2||-2||4|1|||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|424234||4|3|45
501526664|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-25|2013-02-19|Followup|2013-02-25|2013-02-19|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|3|3|4|3|4|3.33|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Yellow|Amachi|Volunteer: Moved|47.8||1|1|1|1|F|White||15|Yes|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|F|White||35|28269|Bachelors Degree|Single|Business: Sales|33609|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|501526956|1|0|2|501233757|1|0|2|500332719|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7496|10|||1|424247||4|3|45
501247269|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-21|NaT|Followup|2013-02-21|2013-01-09|Complete|Early|3|1|1|1|1|1|1.33|||||||||1|1|4|1|1|4|2|||||||||2|2|2|2||||||3|2|2|2|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI, Cabarrus County||72.8||2|2|1|1|F|White||15|No|Father|28025|One Parent: Male|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|White||43|28027|Associate Degree|Married|Student: College||4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500341682|1|0|2|501914025|1|0|2|500515263|2||500016307||2|1|500005291, 500016374|500016374|-2|500016374|-2|0|10|||7496|10|||1|424267||4|3|45
502941572|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-16|2013-04-22|Followup|2013-04-16|2013-04-22|Declined|Done||||||||4|2|2|1|3|3|2.5|||||||||2|3|3|3|2|3|2.67||||||3|3|3|3|||||||4|3|4|5|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|2|2.5||||1|1||||4|4||Green|Amachi|Child/Family: Moved|12.2||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community|Amachi|Match Support|F|White||44|28269|PHD|Single|Medical|64506|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502942998|31|0|2|502884011|1|0|2|500608269|2||-2||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|424329|420804|4|1|45
501314104|BBBS of Greater Charlotte|Main Office|C|Active|2008-12-04|NaT|Followup|2012-12-04|2013-01-15|Complete|Done|4|3|4|1|1|4|2.83|||||||||2|4|4|3|4|4|3.5|||||||||4|4|4|4||||||5|3|4|1|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|4|3.5|||||2|2||||4|4||||Yellow|||99.4||1|1|1|1|M|Black||13|No|Mother|28217|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28134|Bachelors Degree|Single|Business: Mgt, Admin||6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501314382|31|0|1|501170940|1|0|1|500315948|2||-2||2|2|||-2||-2|0|10|||7464|9|||1|424468||4|3|45
502896701|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2013-04-29|Baseline|2012-04-18|2012-04-30|Complete|Done|4|1|3|3|3|3|2.83|||||||||2|3|2|3|3|3|2.67|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|12||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|$40,000 to $44,999||No||Self|General Community||Match Support|M|White||64|28216|Juris Doctorate (JD)|Divorced|Law: Lawyer||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502898109|31|0|1|502888938|1|0|1|500610476|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|425053|-1|4|3|44
502478428|BBBS of Greater Charlotte|Main Office|C|Active|2011-04-28|NaT|Followup|2013-04-28|2013-04-24|Complete|Done|4|4|4|4|4|4|4|4|4|1|4|4|4|3.5|14.29|4|4|4|4|4|4|4|4|2|4|2|4|4|3.33|20.12|4|4|4|4|4|4|4|4|0|4|5|4|4|4.25|4|5|5|5|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|2|3|2.5|2|4|3|-16.67|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||70.6||1|1|1|1|M|White||16|No|Mother|28277|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||54|28205|Some College|Separated|Self-Employed, Entrepreneur|28214|29|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502478875|1|0|1|502555822|1|0|1|500533009|2||-2||2|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|425602|270021|4|3|45
502885468|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-30|NaT|Baseline|2012-04-19|2012-04-30|Complete|Done|4|4|4|4|1|4|3.5|||||||||4|4|4|1||3||||||||||1|4|1|2||||||3|3|2|1|2.25|||||||2|1|3|4|4|4|4|3.14||||||||||1|1|1|1||||||1|2|1.5|||||1|1||||4|4||||Green|||58.5||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Black||47|28227|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502886874|31|0|1|502954219|31|0|1|500610806|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|425685|-1|4|3|44
502845758|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-19|2015-09-16|Followup|2013-04-19|2013-06-03|Declined|Done||||||||4|2|4|2|3|4|3.17|||||||||1|3|3|2|2|4|2.5||||||4|3|3|3.33|||||||3|4|4|2|3.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|1|1.5||||1|1||||4|4||Red||Volunteer: Lost contact with child/agency|40.9||1|1|1|1|M|Black||15|No|Mother|28202|One Parent: Male|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28277||Single|Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502847118|31|0|1|502944923|1|0|1|500606912|2||-2||4|3|||-2||-2|34|2|||7464|9|||1|425782|417837|4|1|45
500765381|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-26|2015-10-20|Followup|2013-02-26|2013-04-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|79.7||1|1|1|1|M|Black||16|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|10019|Bachelors Degree|Single|Business: Marketing|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500739190|31|0|1|501579025|1|0|1|500342803|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|426159||4|1|45
501015965|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-29|2013-10-09|Followup|2013-04-29|2013-04-24|Complete|Done|4|3|4|3|4|4|3.67|||||||||3|3|4|3|2|4|3.17|||||||||4|4|3|3.67||||||5|3|4|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||3|2|3|2.67||||||4|4|4|||||2|2||||4|4||||Yellow|Amachi|Child: Lost interest|41.4||2|2|2|2|F|Black||17|Yes|Mother|28208|One Parent: Female|Less than $10,000||Yes||Self|General Community|Amachi|Match Support|F|Black||60|28269|Bachelors Degree|Married|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|500189376|31|0|2|500447721|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|426856||4|3|45
500361200|BBBS of Greater Charlotte|Main Office|C|Active|2006-03-21|NaT|Followup|2013-03-21|2013-04-29|Complete|Done|2|2|3|2|2|3|2.33|||||||||2|3|3|1|3|3|2.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Cabarrus County||131.8||2|2|1|1|F|White||17|No|Mother|28027|Two Parent|Unknown||No||Relative|General Community|Cabarrus County|Match Support|F|White||32|28115|Bachelors Degree|Single|Human Services: Social Worker||0|0|other|College Partner|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500361450|1|0|2|500368628|1|0|2|500085591|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|3|||7670|5|||1|426936||4|3|45
500799303|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-27|2016-08-19|Followup|2013-03-27|2013-03-21|Complete|Done|3|4|4|2|2|4|3.17|||||||||2|4|3|3|3|3|3|||||||||3|3|3|3||||||2|4|4|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|112.8||1|1|1|1|M|White||19|No|Mother|28081|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||46|28202||Single|Business: Sales||0|4|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500799571|1|0|1|500798390|1|0|1|500167062|2||-2||4|3||500016374|-2|500016374|-2|34|2|||7464|9|||1|426941||4|3|45
501074345|BBBS of Greater Charlotte|Main Office|C|Active|2008-03-31|NaT|Followup|2013-03-31|2013-03-25|Complete|Done|4|1|4|1|1|4|2.5|||||||||4|1|4|4|4|4|3.5|||||||||4|4|4|4||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Green|Amachi, Cabarrus County||107.5||1|1|1|1|M|White||16|Yes|GrandMother|28025|Grandparents|Unknown||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|White||46|28027|Bachelors Degree|Divorced|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501074618|1|0|1|501158523|1|0|1|500250038|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|5635|9|||46|2|||1|426942||4|3|45
502570188|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Followup|2013-04-30|2013-04-30|Complete|Done|4|4|4|3|4|4|3.83|4|3|3|2|4|4|3.33|15.02|4|4|3|4|4|4|3.83|2|4|4|2|3|4|3.17|20.82|4|4|4|4|4|4|4|4|0|5|4|4|4|4.25|5|5|5|4|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|3|3.33|4|4|4|4|-16.75|4|4|4|2|2|2|100|2|2|2|2|0|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|69.8||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||56|28226|Masters Degree|Married|Medical: Nurse|28217|34|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570642|31|0|2|502366830|1|0|2|500533448|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||10326|3|||1|427002|271777|4|3|45
502255156|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-24|NaT|Followup|2013-04-24|2013-07-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||58.7||2|2|1|1|F|Black||14|Yes|Relative: Other|28227|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||35|28277|Masters Degree|Single|Education: Admin||8|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|502255582|31|0|2|502946412|1|0|2|500608992|2||500003586||2|1|500000294|500000294|-2||-2|0|5|||7462|13|||1|427231||4|0|45
502868925|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-25|2014-09-24|Followup|2013-04-25|2013-06-17|Declined|Late||||||||3|1|2|1|3|3|2.17|||||||||2|4|4|1|2|3|2.67||||||4|3|3|3.33|||||||3|4|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|3|2.5||||2|2||||4|4||Red||Child/Family: Lost contact with volunteer/agency|29||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||35|28262|Bachelors Degree|Divorced|Finance: Banking||2|6|Charlotte Cares|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502870324|31|0|2|502885744|31|0|2|500607510|2||-2||4|3|||-2||-2|0|4|||11246|6|||1|427848|419518|4|1|45
502255150|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-14|NaT|Followup|2013-02-14|2013-01-15|Complete|Early|4|1|1|2|4|4|2.67|1|2|1|1|1|4|1.67|59.88|1|3|2|1|3|3|2.17|1|4|3|1|1|3|2.17|0|4|4|4|4|4|4|4|4|0|1|5|5|1|3|2|3|3|2|2.5|20|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|2|1|1|1.33|4|4|3|3.67|-63.76|2|2|2|1|1|1|100|2|2|2|2|0|4|4||||Green|Amachi||73||1|1|1|1|F|Black||17|Yes|Relative: Other|28227|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||34|28212|Masters Degree|Single|Education: Teacher|28216|6|3|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020752|502255582|31|0|2|502392989|1|0|2|500512287|2||500003586||2|1|500000294|500000294|-2|500000294, 500004640|-2|0|5|||7464|9|||1|429730|235505|4|3|45
500392419|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-06|2013-08-29|Followup|2013-03-06|2013-04-12|Complete|Done|3|2|2|2|3|4|2.67|||||||||2|2|3|2|2|4|2.5|||||||||4|4|4|4||||||5|4|4|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Yellow||Child/Family: Moved|77.8||2|2|1|1|F|Black||21||Father|28105|One Parent: Male|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||32|28277||Single|Business: Sales||0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500392669|31|0|2|500746900|1|0|2|500162012|2||-2||4|2|||-2||-2|6855|8|||7464|9|||1|429755||4|3|45
502320003|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2014-09-24|Followup|2013-04-30|2013-06-14|Complete|Done|4|3|3|2|4|4|3.33|4|2|4|4|3|4|3.5|-4.86|3|4|4|4|4|4|3.83|2|3|4|1|2|4|2.67|43.45|4|4|4|4|4|4|4|4|0|5|4|4|4|4.25|4|3|5|4|4|6.25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|4|3|3.5|4|1|2.5|40|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Moved|28.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||30|28216||Single|Tech: Research/Design||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502320438|31|0|2|502810883|31|0|2|500606071|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|429766|416362|4|3|45
502319984|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-03-24|Followup|2013-04-30|2013-06-17|Declined|Late||||||||3|3|4|4|4|4|3.67|||||||||2|4|3|2|2|4|2.83||||||4|4|4|4|||||||3|3|4|4|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|3|3.5||||2|2||||4|4||Red||Volunteer: Time constraint|34.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Bachelors Degree|Single|Finance|28216|3|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502320419|31|0|1|502290677|1|0|1|500607367|2||-2||4|3||500005291|-2||-2|6854|8|||17161|11|||1|429774|418895|4|1|45
502885468|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-30|NaT|Followup|2013-04-30|2013-04-29|Complete|Done|3|4|4|2|4|4|3.5|4|4|4|4|1|4|3.5|0|2|4|4|2|4|4|3.33|4|4|4|1||3|||4|4|4|4|1|4|1|2|100|4|3|5|3|3.75|3|3|2|1|2.25|66.67|4|4|4|4|4|4|4|4|2|1|3|4|4|4|4|3.14|27.39|4|4|4|4|1|1|1|1|300|2|1|1.5|1|2|1.5|0|2|2|1|1|100|4|4|4|4|0|Green|||58.5||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Black||47|28227|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502886874|31|0|1|502954219|31|0|1|500610806|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|429792|425685|4|3|45
502319972|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-08-19|Followup|2013-04-30|2013-06-17|Declined|Late||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|3|4|4|3.83||||||4|4|4|4|||||||4|4|3|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4||||1|1||||4|4||Yellow||Volunteer: Moved|39.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Less than $10,000||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||32|28214|Bachelors Degree|Married|Self-Employed, Entrepreneur|29715|0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502320407|31|0|1|502911091|1|0|1|500607368|2||-2||4|2||500005291|-2||-2|6854|8|||7464|9|||1|429795|418896|4|1|45
502859599|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2014-05-05|Followup|2013-04-30|2013-04-30|Complete|Done|4|1|4|4|4|3|3.33|3|1|2|1|3|4|2.33|42.92|2|3|3|2|2|3|2.5|4|4|4|4|4|4|4|-37.5|4|3|3|3.33|4|4|4|4|-16.75|4|4|4|4|4|5|4|4|5|4.5|-11.11|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|3|4|3.67|8.99|4|4|4|2|3|2.5|60|2|2|1|1|100|3|3|4|4|-25|Green||Volunteer: Lost contact with child/agency|24.1||1|1|1|1|M|Hispanic|Other Central American|14|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|Hispanic|Other South American|35|28209|High School Graduate|Married|Business||0|1|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500017777|502860998|3|14|1|502864237|3|15|1|500610310|2||-2||4|1|||-2||-2|0|4|||17161|11|||1|429888|410107|4|3|45
500814240|BBBS of Greater Charlotte|Main Office|C|Active|2008-04-24|NaT|Followup|2013-04-24|2013-04-22|Complete|Done|1|2|3|3|2|3|2.33|||||||||3|2|4|3|2|4|3|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||106.7||1|1|1|1|M|Black||18|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||46|28215|Bachelors Degree|Single|Business: Mgt, Admin|28226|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500814509|31|0|1|500981509|31|0|1|500248568|2||500003586||2|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|430160||4|3|45
501222138|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2015-05-07|Followup|2013-04-30|2013-04-24|Complete|Done|3|1|4|4|4|4|3.33|||||||||2|4|3|2|4|3|3|||||||||4|3|4|3.67||||||2|2|4|5|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|2|2.5|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|60.2||2|2|2|3|F|Black||14|Yes|GrandMother|28227|Grandparents|Unknown||No||Self|General Community|Amachi|Enrollment|F|Black||53|28269|Some College|Married|Business: Sales|28227|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501222414|31|0|2|500189173|31|0|2|500447311|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|430314||4|3|45
501160887|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2013-05-14|Followup|2013-04-30|2013-04-24|Complete|Done|4|3|4|3|4|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|3|4|4|4|4|4|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|36.5||2|2|1|1|F|Black||14|Yes|Mother|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Enrollment|F|White||58|28226|||Education: Teacher Asst/Aid|28203|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|501016235|31|0|2|501615415|1|0|2|500447312|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|430318||4|3|45
502828137|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-06-29|Followup|2013-04-30|2013-06-14|Comprehension|Done||||||||3|1|1|3|1|1|1.67|||||||||1|2|2|2|1|3|1.83||||||4|4|4|4|||||||2|2|4|2|2.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Green||Child/Family: Moved|37.9||1|1|1|1|F|Multi-Race (None of the above)||16|No|Father|28214|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher|28078|0|8|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502829415|7|0|2|502446364|31|0|2|500607445|2||-2||4|1|||-2|500004640|-2|0|10|||7464|9|||1|430602|419338|4|2|45
502828131|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-03-31|Followup|2014-04-30|2014-06-14|Complete|Done|4|2|3|3|3|3|3|4|4|4|3|4|4|3.83|-21.67|2|3|3|3|3|3|2.83|2|4|3|3|4|3|3.17|-10.73|4|3|3|3.33|4|4|4|4|-16.75|3|3|3|3|3|4|5|4|2|3.75|-20|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|4|3|1|2.67|37.45|1|2|1.5|3|3|3|-50|2|2|1|1|100|4|4|4|4|0|Red||Child/Family: Lost contact with volunteer/agency|35||1|1|1|1|F|Multi-Race (None of the above)||17|No|Father|28214|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|White||33|28216|Bachelors Degree|Single|Business: Sales|28270|2|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502829415|7|0|2|502881454|1|0|2|500607446|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|430607|419339|4|3|45
502828146|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2014-05-30|Followup|2013-04-30|2013-05-09|Declined|Done||||||||2|2|3|2|2|1|2|||||||||2|2|3|2|2|2|2.17||||||4|4|4|4|||||||2|2|3|2|2.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Red||Volunteer: Lost contact with child/agency|25||1|1|1|1|M|Black||17|No|Father|28214|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|Black||37|28278|Bachelors Degree|Single|Unknown||0|0|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502829415|31|0|1|502860825|31|0|1|500607619|2||-2||4|3|||-2||-2|0|10|||9229|13|||1|430611|419662|4|1|45
501662033|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-03|2014-03-20|Followup|2013-03-03|2013-04-30|Complete|Late|3|2|2|4|3|3|2.83|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|3|2|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|24.5||2|2|4|4|F|Black||13|No|Mother|28215|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Enrollment|F|Black||38|28219||Single|Finance: Banking|28273|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501090456|31|0|2|500459674|31|0|2|500597964|2||-2||4|1|||-2|500000294|-2|0|10|||2238|7|||1|430648||4|3|45
502307585|BBBS of Greater Charlotte|Main Office|C|Active|2011-03-21|NaT|Followup|2013-03-21|2013-04-12|Complete|Done|4|2|2|2|3|3|2.67|4|1|2|1|1|1|1.67|59.88|3|2|3|3|3|2|2.67|2|2|4|1|2|3|2.33|14.59|3|3|3|3|4|4|4|4|-25|3|4|5|5|4.25|4|5|5|5|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|3|3|3|16.67|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi||71.9||1|1|1|1|F|Black||17|Yes|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||53|28031||Divorced|Medical: Admin|28207|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500020910|502308017|31|0|2|501519450|1|0|2|500521250|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|4|||7446|3|||1|431139|251051|4|3|45
500781988|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-16|2013-09-04|Followup|2013-02-16|2013-05-03|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|78.6||1|1|1|1|M|White||21||Mother|28027||Unknown||No||Self|General Community||Match Support|M|White||71|28083|Some College|Married|Business: Mgt, Admin|28027|13|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500002335|500782256|1|0|1|500773716|1|0|1|500160560|2||-2||4|1|||-2||-2|0|10|||46|2|||1|431241||4|0|45
501631547|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2016-07-29|Followup|2013-03-31|2013-03-27|Complete|Done|3|3|3|3|3|3|3|||||||||2|4|3|1|1|3|2.33|||||||||4|4|4|4||||||4|3|3|1|2.75|||||||3|4|4|4|3|4|3|3.57||||||||||1|4|2|2.33||||||3|2|2.5|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child: Graduated|64||2|2|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||38|28277|Bachelors Degree|Single|Arts, Entertainment, Sports|28203|3|6|UnitedMethodistChrch|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|501631870|31|0|1|502170945|1|0|1|500528464|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||8529|7|||1|431424||4|3|45
501868918|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-27|2014-05-22|Followup|2013-05-27|2013-05-23|Complete|Done|3|4|4|4|2|3|3.33|3|3|3|4|3|3|3.17|5.05|4|4|4|4|4|4|4|3|4|4|2|3|3|3.17|26.18|4|3|3|3.33|4|4|3|3.67|-9.26|3|4|5|3|3.75|3|3|5|5|4|-6.25|4|4|4|4|4|4|3|3.86|3|4|3|3|4|3|2|3.14|22.93|2|4|2|2.67|3|4|3|3.33|-19.82|2|2|2|2|3|2.5|-20|2|2|1|1|100|4|4||||Green||Child: Graduated|47.8||1|1|1|1|M|Black||20|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||35|27612|Juris Doctorate (JD)|Living w/ Significant Other|Law|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|501869291|31|0|1|501921115|1|0|1|500454496|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|431428|128915|4|3|45
501868921|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2016-07-29|Followup|2013-03-31|2013-04-18|Complete|Done|3|3|4|4|3|4|3.5|3|1|1|1|1|2|1.5|133.33|3|4|3|4|2|3|3.17|3|2|4|4|4|4|3.5|-9.43|4|2|2|2.67|4|3|3|3.33|-19.82|3|5|4|5|4.25|4|5|5|4|4.5|-5.56|4|4|3|3|2|2|2|2.86|4|4|4|4|3|3|3|3.57|-19.89|3|3|2|2.67|2|4|3|3|-11|2|3|2.5|2|1|1.5|66.67|2|2|1|1|100|4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Moved|64||2|2|2|2|F|Black||19|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28211||Married|Finance: Banking|28255|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501869291|31|0|2|501382633|1|0|2|500524206|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|431431|4527|4|3|45
501247286|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-14|2016-11-08|Followup|2013-05-14|2013-05-13|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|101.8||1|1|1|1|M|White||15|No|Father|28025|One Parent: Male|Unknown||No||Self|General Community|Cabarrus County|Enrollment|M|White||49|27103|Masters Degree|Single|Education: Teacher|27282|0|0|Other|Service Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500341682|1|0|1|501247141|1|0|1|500264655|2||-2||4|1||500016374|-2|500016374|-2|0|10|||7452|6|||1|431629||4|3|45
502961272|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-21|2014-01-29|Baseline|2012-05-02|2012-05-21|Complete|Done|4|2|3|3|2|2|2.67|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||4|2|2|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||2|2|4|2.67||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Child/Family: Moved|20.3||1|1|1|1|F|White||17|Yes|Mother|28205|Grandparents|$25,000 to $29,999||Yes||Self|General Community|Amachi|Match Support|F|White||62|28299|Some College|Divorced|Business: Sales||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502962447|1|0|2|503009515|1|0|2|500614268|2||-2||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|431654|-1|4|3|44
501811385|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-23|2016-08-19|Followup|2013-03-23|2013-03-12|Complete|Done|4|4|4|3|3|4|3.67|||||||||4|4|4|1|2|4|3.17|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI, Cabarrus County|Child: Graduated|64.9||2|2|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||43|28075|Bachelors Degree|Married|Business: Mgt, Admin||7|0|Recruitment Event|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501811730|31|0|2|502460013|31|0|2|500524684|2||-2||4|3|500005291, 500016374|500016374|-2|500016374|-2|6854|8|||7459|10|||1|431739||4|3|45
502530227|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2014-10-20|Followup|2013-05-04|2013-06-07|Complete|Done|3|3|3|1|3|3|2.67|4|1|1|2|4|4|2.67|0|3|4|4|4|4|4|3.83|2|4|4|2|3|4|3.17|20.82|4|4|4|4|4|4|4|4|0|4|4|4|4|4|5|5|4|5|4.75|-15.79|4|4|4|4|4|4|4|4|4|4|4|3|4|3|4|3.71|7.82|4|4|4|4|3|4|3|3.33|20.12|4|3|3.5|2|4|3|16.67|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|41.6||1|1|1|1|F|Hispanic||15|No|Mother|28213|One Parent: Female|$10,000 to $14,999||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||30|28210|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502530676|3|0|2|502531485|3|0|2|500532078|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|432130|268895|4|3|45
501575257|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-18|2013-09-24|Followup|2013-03-18|2013-04-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|54.2||1|1|1|1|M|Black||15|No|Mother|28079|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||38|28079||Married|Law: Police Officer|28211|5|0|Recruitment Event|Self|Big|General Community||Enrollment|277|60|598|500000170|500004169|501575553|31|0|1|501234758|1|0|1|500348757|2||-2||4|3|||-2||-2|0|10|||7458|9|||1|432496||4|1|45
501621811|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-16|2017-03-09|Followup|2013-03-16|2013-02-12|Complete|Early|3|4|4|1|3|4|3.17|||||||||1|3|3|2|2|3|2.33|||||||||4|4|4|4||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|4|3.5|||||2|2||||4|4||||Yellow|Project Big|Child/Family: Lost contact with volunteer/agency|95.8||1|1|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||36|28269||Married|Self-Employed, Entrepreneur|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501622131|31|0|2|501621016|31|0|2|500344465|2||-2||4|2|500004640||-2||-2|0|10|||7464|9|||1|432497||4|3|45
502637403|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-24|2014-03-31|Baseline|2012-05-04|2012-05-24|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|2|3|4|3.33|||||||||4|3|3|3.33||||||4|3|4|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|22.2||1|1|1|1|F|Black||15|Yes|Mother|28278|One Parent: Female|$30,000 to $34,999||No||School|General Community|Amachi|Match Support|F|White||24|28105|Some College||Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|502638098|31|0|2|502883455|1|0|2|500613355|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|4|||46|2|||1|432517|-1|4|3|44
500740296|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-04|NaT|Followup|2013-05-04|2013-04-30|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|||58.4||2|2|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Therapist/Counselor|General Community||Match Support|F|Asian||32|28216|Bachelors Degree|Single|Business: Mgt, Admin|28208|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500740560|31|0|2|502893901|4|0|2|500611525|2||-2||2|2|||-2||-2|0|5|||7464|9|||1|432563||4|3|45
502866443|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-14|2014-09-23|Baseline|2012-05-04|2012-06-14|Complete|Done|4|1|2|1|3|4|2.5|||||||||1|3|3|1|2|4|2.33|||||||||4|2|4|3.33||||||5|3|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|1|2.5|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|27.3||1|1|1|1|F|Black||14|No|Mother|28262|One Parent: Female|$30,000 to $34,999|Y|No||Self|General Community||Match Support|F|Black||38|28212|Some College|Single|Business: Mgt, Admin|28270|7|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502867844|31|0|2|502920462|31|0|2|500613414|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|432716|-1|4|3|44
502966254|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-04|2015-03-18|Followup|2013-05-04|2013-05-28|Complete|Done|3|2|4|4|2|4|3.17|2|3|2|4|2|3|2.67|18.73|2|4|3|2|3|3|2.83|2|4|3|2|2|3|2.67|5.99|4|4|4|4|4|3|4|3.67|8.99|3|5|3|5|4|3|4|2|2|2.75|45.45|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|1|1.5|4|4|4|-62.5|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Lost contact with child/agency|34.4||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community||Match Support|F|Black||48|28217|Bachelors Degree|Divorced|Medical: Admin|28232|11|5|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|500784955|31|0|2|502895517|31|0|2|500609631|2||-2||4|2|||-2||-2|0|10|||7438|1|||1|432717|423139|4|3|45
502997008|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-30|2013-07-17|Baseline|2012-05-07|2012-05-30|Complete|Done|2|2|2|2|2|2|2|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|5|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Yellow||Volunteer: Unrealistic expectations|13.6||2|2|1|1|F|Black||17|No|Mother|28226|Two Parent|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||31|28273|Juris Doctorate (JD)|Single|Law: Lawyer||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|502998473|31|0|2|502908444|31|0|2|500613594|2||-2||4|2|||-2||-2|34|2|||7464|9|||1|433513|-1|4|3|44
500727291|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-17|2016-07-29|Followup|2013-05-17|2013-05-09|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|110.4||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|Black||46|28269|||Human Services: Non-Profit||0|0|BBBS National Site|Web Link|Big|General Community|VOL - Adjudicated, VOL - Cultural Comp, VOL - PreMatch|Match Support|277|60|598|500000170|500008321|500727558|31|0|1|500857838|31|0|1|500176403|2||-2||4|1|||-2|500007913, 500007920, 500011311|-2|0|10|||46|2|||1|433548||4|3|45
502469110|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-11|2014-03-03|Followup|2013-05-11|2013-06-07|Complete|Done|4|2|3|2|3|3|2.83|3|3|3|2|4|3|3|-5.67|4|4|3|3|3|4|3.5|2|4|3|2|2|3|2.67|31.09|4|4|4|4|4|4|4|4|0|5|5|5|5|5|2|5|3|4|3.5|42.86|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|4|3.5|4|3|3.5|0|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Moved|33.7||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||35|28269|Associate Degree|Married|Arts, Entertainment, Sports|28262|3|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502469557|31|0|1|502564995|31|0|1|500535534|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7496|10|||1|433590|277903|4|3|45
502596391|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-12|2013-08-20|Followup|2013-06-12|2013-07-14|Complete|Done|4|2|4|3|4|4|3.5|3|4|4|4|4|4|3.83|-8.62|4|4|4|3|3|3|3.5|3|4|3|4|4|3|3.5|0|4|4|4|4|4|2|2|2.67|49.81|4|4|5|5|4.5|2|3|5|3|3.25|38.46|4|4|4|4|4|4|4|4|4|4|4|3|1|3|2|3|33.33|4|4|4|4|3|4|2|3|33.33|4|2|3|1|4|2.5|20|2|2|2|2|0|4|4|4|4|0|Yellow|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|26.3||1|1|2|2|F|Black||16|No|Mother|28208|Two Mothers|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502596909|31|0|2|502485670|31|0|2|500540403|2||500004641||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7462|13|1204|3|1|433619|284319|4|3|45
501143674|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-08|2016-08-05|Followup|2013-05-08|2013-06-19|Complete|Done|3|2|3|2|2|3|2.5|3|4|3|3|1|3|2.83|-11.66|2|3|4|3|2|4|3|2|2|2|3|2|4|2.5|20|4|4|4|4|2|3|3|2.67|49.81|4|4|4|4|4|2|4|3|3|3|33.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|3|3|3|2|2|2|50|2|2|2|2|0|4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|50.9||3|3|1|1|F|Black||16||Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||28|28211|Bachelors Degree|Single|Human Services||2|0|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|277|60|598|500000170|500008321|501143948|31|0|2|502958999|1|0|2|500612879|2||500004641||4|2|||-2||-2|0|10|||132|8|||1|433788|17126|4|3|45
502908460|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-07|2014-09-04|Baseline|2012-05-08|2012-06-07|Complete|Done|4|4|1|3|4|4|3.33|||||||||2|2|2|2|1|3|2|||||||||4|2|2|2.67||||||1|5|3|3|3|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|3|3.67||||||4|1|2.5|||||1|1||||4|4||||Yellow||Volunteer: Lost contact with child/agency|26.9||1|1|1|1|F|Hispanic||18|No|Mother|28227|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||40|28079|Bachelors Degree|Single|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502909871|3|0|2|502938939|1|0|2|500616222|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|434253|-1|4|3|44
501390345|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-08|NaT|Followup|2013-05-08|2013-05-01|Complete|Done|4|2|2|2|2|3|2.5|||||||||2|2|4|2|2|3|2.5|||||||||4|4|4|4||||||2|3|4|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|Amachi||58.3||2|2|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||35|28206|Bachelors Degree|Single|Business: Sales|28117|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501390617|31|0|1|502966998|1|0|1|500609269|2||-2||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|434353||4|3|45
502863776|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-31|NaT|Baseline|2012-05-09|2012-07-31|Complete|Done|2|2|3|4|3|4|3|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||3|5|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||1|1|1|||||1|1||||4|4||||Green|||55.5||1|1|1|1|F|Black||14|No|Mother|28031|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Mgt, Admin|28078|1|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502865175|31|0|2|503029273|1|0|2|500622877|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|434619|-1|4|3|44
501434147|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2013-03-31|2013-04-12|Complete|Done|4|1|2|2|4|4|2.83|3|1|4|3|1|3|2.5|13.2|3|3|4|3|3|2|3|2|4|4|4|4|4|3.67|-18.26|4|4|4|4|4|4|4|4|0|5|4|3|3|3.75|4|5|2|5|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4||||Green|||83.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||26|28215|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501434432|31|0|1|501926474|31|0|1|500441566|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|435423|29966|4|3|45
501506214|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-28|2016-06-23|Followup|2013-03-28|2013-04-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|86.9||1|1|1|1|M|Black||19|No|Mother|28105|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||55|28173|||Unknown|28203|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501506506|31|0|1|501588885|31|0|1|500351462|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|436390||4|1|45
501626199|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-26|2013-09-30|Followup|2013-03-26|2013-04-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|54.2||1|1|1|1|F|Black||21|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||33|28203|Masters Degree|Single|Finance: Accountant|28211|1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|501622822|31|0|2|501293622|1|0|2|500351814|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|436991||4|1|45
501626218|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-24|2014-12-18|Followup|2013-03-24|2013-04-18|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|3|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|68.8||1|1|1|1|F|Black||20|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||30|11215|Bachelors Degree|Single|Consultant|11215|0|5|other|College Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501622822|31|0|2|501587214|31|0|2|500350222|2||-2||4|1|||-2|500000294|-2|0|10|||7670|5|||1|436993||4|3|45
502259046|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-25|2013-09-16|Followup|2013-05-25|2013-05-22|Complete|Done|4|4|4|4|4|4|4|2|3|4|3|3|4|3.17|26.18|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|5|5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|2|2|1|1|100|4|4||||Yellow||Volunteer: Time constraint|27.8||1|1|1|1|F|White||17|No|Mother|28025|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Enrollment|F|White||64|28083|High School Graduate|Married|Finance: Banking||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502259478|1|0|2|502502361|1|0|2|500537239|2||||4|2|||-2||-2|6854|8|||7464|9|||1|437584|285946|4|3|45
500544921|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2013-08-29|Followup|2013-03-31|2013-04-12|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi|Child: Lost interest|29||2|2|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$15,000 to $19,999|Y|No|TV|Media|General Community|Project Big AND Amachi|Match Support|M|White||31|28211|Bachelors Degree|Married|Finance: Banking|28202|0|2|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011746|500545173|31|0|1|502079132|1|0|1|500523387|2||500004772||4|3|500000294, 500004640, 500004901|500004901|-2||-2|56|1|||7464|9|||1|438054||4|3|45
502997211|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-01|2013-09-05|Baseline|2012-05-15|2012-06-01|Complete|Done|3|1|3|4|4|4|3.17|||||||||1|3|3|3|2|4|2.67|||||||||4|4|3|3.67||||||3|3|2|2|2.5|||||||4|1|4|4|3|4|4|3.43||||||||||4|3|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|15.1||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|F|White||27|28105|Some College||Student: College||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011349|502998689|31|0|2|502926434|1|0|2|500614826|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|438072|-1|4|3|44
502494753|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-14|2013-10-22|Followup|2013-04-14|2013-04-30|Complete|Done|4|3|2|2|3|3|2.83|4|3|3|1|4|3|3|-5.67|2|3|3|2|2|3|2.5|2|3|2|3|1|4|2.5|0|4|4|4|4|4|4|4|4|0|3|2|3|3|2.75|1|4|3|5|3.25|-15.38|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|3|3.33|1|4|4|3|11|4|3|3.5|4|2|3|16.67|2|2|1|1|100|4|4||||Yellow|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|30.3||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28212|Masters Degree|Single|Business|28105|5|8|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500011746|502495202|31|0|2|502481799|31|0|2|500529173|2||500004772||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|4|||7438|1|||1|438844|263617|4|3|45
501919423|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-24|NaT|Followup|2013-03-24|2013-06-08|Expired|Late||||||||4|4|4|4|4|4|4|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||4|5|4|3|4||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|3|3.5||||1|1|||||||Green|Project Big||83.7||1|1|1|1|M|Multi-race (Black & Hispanic)||17|No|Mother|28214|One Parent: Female|Unknown||No|TV|Media|General Community|Project Big|Match Support|M|White||34|28164|Masters Degree||Finance|28210|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501919819|38|0|1|502034798|1|0|1|500442066|2||500004641||2|1|500004640|500004640|-2||-2|56|1|||7464|9|||1|438969|36152|4|0|45
501716720|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-02|2017-02-06|Followup|2013-03-02|2013-05-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Cabarrus County|Child/Family: Lost contact with volunteer/agency|83.2||1|1|1|1|M|Black||15|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||52|28075||Married|Medical: Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501716992|31|0|1|501878786|31|0|1|500435676|2||500016307||4|3|500016374|500016374|-2|500016374|-2|6854|8|||7464|9|||1|439501||4|0|45
502552438|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-02|2017-02-23|Followup|2013-06-02|2013-06-24|Complete|Done|4|2|2|1|4|3|2.67|4|3|4|1|3|4|3.17|-15.77|4|4|3|2|4|3|3.33|4|4|4|2|4|3|3.5|-4.86|4|4|4|4|4|4|4|4|0|5|5|4|4|4.5|5|4|4|5|4.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|4|4|4|2|4|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|68.8||1|1|1|1|M|Black||16|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||36|28205|Masters Degree|Living w/ Significant Other|Journalist/Media|28202|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502552891|31|0|1|502549491|1|0|1|500538826|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||7464|9|||1|439798|292098|4|3|45
502495501|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-20|NaT|Followup|2013-05-20|2013-06-07|Complete|Done|3|1|3|2|1|4|2.33|3|1|4|2|2|2|2.33|0|4|3|4|4|4|4|3.83|2|3|3|1|2|3|2.33|64.38|4|4|4|4|4|4|4|4|0|4|3|3|3|3.25|5|3|2|3|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|3|4|3.67|4|4|3|3.67|0|4|4|4|2|1|1.5|166.67|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||69.9||1|1|1|1|M|White||15|No|Mother|28226|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||55|28210|Bachelors Degree|Married|Finance|28203|1|6|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500018851|502495950|1|0|1|502508181|1|0|1|500531873|2||-2||2|1|500005291|500005291|-2|500005291|-2|0|10|||7464|9|||1|439808|268809|4|3|45
502920377|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-29|2017-02-28|Baseline|2012-05-17|2012-06-29|Complete|Done|3|2|2|2|2|3|2.33|||||||||2|3|2|3|3|3|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|||||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|56||1|1|1|1|F|Black||14|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||31|28211|Bachelors Degree|Single|Real Estate: Realtor|19137|2|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502921794|31|0|2|502942994|1|0|2|500620441|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|439883|-1|4|3|44
502225262|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-10|2013-02-28|Followup|2012-08-10|2012-09-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|30.7||2|2|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown|Y|Yes|AARTF|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||33|28204|Bachelors Degree|Single|Education: Teacher||0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502225693|31|0|2|502244560|31|0|2|500463849|2||500003586||4|2|500000294|500000294|-2|500000294|-2|6855|8|||7496|10|||1|440265||4|1|45
500186141|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-02|2014-04-30|Followup|2013-04-02|2013-05-14|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|3|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green||Child: Graduated|72.9||3|3|1|1|F|Black||20|No|Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||45|28269|Bachelors Degree|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|500187731|31|0|2|501046739|31|0|2|500254296|2||-2||4|1|||-2|500000294|-2|0|10|||46|2|||1|440939||4|3|45
502961272|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-21|2014-01-29|Followup|2013-05-21|2013-07-22|Complete|Late|4|2|2|2|3|2|2.5|4|2|3|3|2|2|2.67|-6.37|2|3|3|3|2|3|2.67|2|4|3|3|2|3|2.83|-5.65|4|4|4|4|4|4|4|4|0|4|4|4|2|3.5|4|2|2|3|2.75|27.27|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|2|2|4|2.67|24.72|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Yellow|Amachi|Child/Family: Moved|20.3||1|1|1|1|F|White||17|Yes|Mother|28205|Grandparents|$25,000 to $29,999||Yes||Self|General Community|Amachi|Match Support|F|White||62|28299|Some College|Divorced|Business: Sales||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502962447|1|0|2|503009515|1|0|2|500614268|2||-2||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|441191|431654|4|3|45
500724632|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-07|NaT|Followup|2013-03-07|2013-05-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||120.3||1|1|1|1|F|Black||17||Mother|28213|One Parent: Female|Less than $10,000|Y|No||School|General Community||Match Support|F|Black||32|28214|Bachelors Degree|Married|Architect|28270|0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|500724899|31|0|2|500803551|31|0|2|500164708|2||-2||2|1|||-2||-2|0|4|||46|2|||1|442008||4|0|45
502570183|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Followup|2013-04-30|2013-04-30|Complete|Done|3|2|3|2|3|3|2.67|3|3|4|3|4|3|3.33|-19.82|1|3|2|3|3|2|2.33|4|4|4|4|4|3|3.83|-39.16|4|4|4|4|4|4|3|3.67|8.99|5|5|4|4|4.5|3|3|4|3|3.25|38.46|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|2|2|0|3|3||||Green|Amachi, Project Big, Project Big AND Amachi|Agency: Challenges with program/partnership|69.8||1|1|1|1|F|Black||17|Yes|Mother|28206|Other/Unknown|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||61|28134|Bachelors Degree|Married|Medical: Admin||33|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570637|31|0|2|502570153|31|0|2|500534090|2||500004772||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|442234|273709|4|3|45
502303088|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2016-08-29|Followup|2013-06-27|2013-07-24|Complete|Done|3|4|4|4|3|4|3.67|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|Project Big|Volunteer: Time constraint|62.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community|Project Big|Enrollment|F|Black||33|28215|Bachelors Degree|Single|Human Services: Social Worker|28217|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017777|502303520|31|0|2|502445797|31|0|2|500533193|2||-2||4|1|500004640|500004640|-2|500000294, 500004640|-2|6854|8|||7464|9|||1|442241||4|3|45
502530223|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2013-05-21|Followup|2013-04-29|2013-04-30|Declined|Done||||||||3|2|1|1|2|2|1.83|||||||||1|3|2|1|2|2|1.83||||||3|4|4|3.67|||||||3|2|4|4|3.25||||||||||4|4|4|4|4|4|4|4||||||3|4|4|3.67|||||4|4|4||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|24.7||1|1|1|1|M|Hispanic||16||Mother|28213|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||44|28078|Masters Degree|Married|Business|28036|8|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502530676|3|0|1|502501248|3|0|1|500533054|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|442247|269200|4|1|45
500850236|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-04|2013-09-16|Followup|2013-04-04|2013-04-12|Complete|Done|3|2|2|2|3|3|2.5|||||||||1|4|4|2|2|3|2.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green||Child: Graduated|77.4||1|1|2|2|M|Black||21|No|Mother|28205|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|Black||37|28262|Bachelors Degree|Single|Real Estate: Realtor||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|500850505|31|0|1|500189198|31|0|1|500169235|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|442250||4|3|45
502578459|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-23|NaT|Baseline|2012-05-22|2012-07-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Cabarrus County||55.8||1|1|1|1|M|Black||18|No|Mother|28025|One Parent: Female|$35,000 to $39,999||Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||48|28269|Some College|Married|Tech: Management|28204|10|0|AA Task Force|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502578962|31|0|1|502869485|31|0|1|500615803|2||500016307||2|2|500016374|500016374|-2|500016374|-2|6854|8|||9229|13|||1|442607|-1|4|1|44
502287066|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-03|2014-09-04|Followup|2013-05-03|2013-06-07|Complete|Done|4|2|4|2|4|3|3.17|||||||||4|4|4|4|2|3|3.5|||||||||4|3|4|3.67||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|40.1||2|2|1|1|M|Black||15||GrandMother|28227|One Parent: Female|Unknown|Y|Yes|AARTF|BBBS Board/Staff|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28215|Associate Degree|Married|Medical: Nurse||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502287498|31|0|1|502501212|1|0|1|500532817|2||-2||4|1|500005291|500005291|-2||-2|7294|13|||7464|9|||1|442794||4|3|45
502866475|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-23|NaT|Followup|2013-05-23|2013-06-13|Complete|Done|3|2|3|2|3|2|2.5|4|4|4|4|4|4|4|-37.5|4|3|4|4|4|4|3.83|3|4|4|2|4|4|3.5|9.43|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|3|3|4|3.75|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Green|||57.8||1|1|1|1|M|Black||16|No|Mother|28270|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|M|White||29|28203|Bachelors Degree||Finance: Accountant||1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502867876|31|0|1|502961396|1|0|1|500614954|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|443332|418831|4|3|45
502868923|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-27|2015-10-30|Followup|2013-01-27|2013-02-09|Complete|Done|4|3|3|2|3|4|3.17|||||||||2|4|3|3|4|3|3.17|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Volunteer: Moved|45.1||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Black||28|28262|Bachelors Degree|Single|Finance: Banking||0|0|AA Task Force|Special Event|Big|General Community||Match Support|277|60|598|500000170|500008321|502870324|31|0|2|502832013|31|0|2|500591320|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||11098|8|||1|444190||4|3|45
502637403|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-24|2014-03-31|Followup|2013-05-24|2013-06-25|Declined|Done||||||||4|4|4|4|4|4|4|||||||||3|4|4|2|3|4|3.33||||||4|3|3|3.33|||||||4|3|4|5|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Green|Amachi|Child/Family: Lost contact with volunteer/agency|22.2||1|1|1|1|F|Black||15|Yes|Mother|28278|One Parent: Female|$30,000 to $34,999||No||School|General Community|Amachi|Match Support|F|White||24|28105|Some College||Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|502638098|31|0|2|502883455|1|0|2|500613355|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|4|||46|2|||1|444242|432517|4|1|45
500186245|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-24|NaT|Followup|2013-05-24|2013-06-10|Complete|Done|4|3|4|2|3|4|3.33|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||4|5|3|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|1|2.33||||||2|1|1.5|||||2|2||||4|4||||Green|Amachi||57.7||2|3|1|1|M|Black||16|Yes|Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|M|White||34|28203|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500187840|31|0|1|502989318|1|0|1|500614903|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|444762||4|3|45
502874566|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-24|2015-10-16|Followup|2013-05-24|2013-05-17|Complete|Done|4|4|4|4|3|4|3.83|3|1|3|1|3|4|2.5|53.2|4|4|4|2|4|4|3.67|2|3|4|2|3|4|3|22.33|4|4|4|4|4|4|4|4|0|5|5|5|5|5|4|4|5|5|4.5|11.11|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|2|4|3|4|4|4|-25|2|2|2|2|0|4|4||||Green||Volunteer: Moved|40.7||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|White||28|27235|Bachelors Degree||Business: Engineer||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502875969|3|10|2|502894480|1|0|2|500607372|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|444854|411252|4|3|45
500186798|BBBS of Greater Charlotte|Main Office|C|Completed|2005-03-30|2015-10-20|Followup|2013-03-30|2013-04-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Time constraints|126.7||1|2|1|2|F|Multi-Race (None of the above)||19|No|Father|28208|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||45|28226|Bachelors Degree||Business: Human Resources||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500187961|7|0|2|500189825|1|0|2|500038158|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|445403||4|1|45
502393980|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-25|NaT|Followup|2013-05-25|2013-06-25|Complete|Done|3|2|2|1|3|3|2.33|3|1|1|1|3|3|2|16.5|2|2|3|2|2|2|2.17|2|3|2|2|2|3|2.33|-6.87|4|4|4|4|4|4|4|4|0|3|3|3|3|3|2|3|5|5|3.75|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|2|3|2|2.33|1|4|1|2|16.5|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green|Amachi||57.7||2|2|1|1|F|Multi-race (Black & White)||16|Yes|Aunt|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28078|Associate Degree|Married|Tech: Support, Writing|28210|2|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502394418|36|0|2|502928199|31|0|2|500613992|2||500003586||2|1|500000294|500005291|-2||-2|0|5|||7462|13|||1|445432|254548|4|3|45
502632678|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-08|2012-09-14|Baseline|2012-05-25|2012-06-07|Complete|Done|4|3|3|3|3|3|3.17|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||5|2|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||1|1||||4|4||||Yellow||Child: Family structure changed|3.2||1|1|1|1|M|Black|Other African|17|No|Mother|28212|One Parent: Female|$20,000 to $24,999|Y|Yes||Relative|General Community||Match Support|M|Black||54|28269|Masters Degree|Single|Tech: Computer/Programmer|28212|5|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500001281|502633334|31|31|1|503007956|31|0|1|500616542|2||-2||4|2|||-2||-2|0|3|||7462|13|||1|445569|-1|4|3|44
502980965|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-18|2013-01-09|Baseline|2012-05-29|2012-06-18|Complete|Done|2|1|1||3|4||||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Red||Volunteer: Time constraint|6.7||2|2|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||40|28209|Bachelors Degree|Single|Finance: Banking|28255|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|502982410|31|0|2|503007163|1|0|2|500618600|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|447655|-1|4|3|44
502997008|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-30|2013-07-17|Followup|2013-05-30|2013-06-06|Declined|Done||||||||2|2|2|2|2|2|2|||||||||2|3|3|3|3|3|2.83||||||4|4|4|4|||||||3|5|4|3|3.75||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||4|4|4||||1|1||||4|4||Yellow||Volunteer: Unrealistic expectations|13.6||2|2|1|1|F|Black||17|No|Mother|28226|Two Parent|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||31|28273|Juris Doctorate (JD)|Single|Law: Lawyer||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500004169|502998473|31|0|2|502908444|31|0|2|500613594|2||-2||4|2|||-2||-2|34|2|||7464|9|||1|448618|433513|4|1|45
501599416|BBBS of Greater Charlotte|Main Office|C|Active|2009-04-28|NaT|Followup|2013-04-28|2013-05-22|Complete|Done|4|4|4|4|2|4|3.67|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|||94.6||1|1|1|1|M|White||14|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||46|28078|Masters Degree|Single|Retail: Mgt|28207|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501599736|1|0|1|500188567|1|0|1|500357914|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|449652||4|3|45
502180719|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-04|2014-03-20|Followup|2013-06-04|2013-06-03|Complete|Done|4|4|4|3|4|4|3.83|4|2|4|4|4|4|3.67|4.36|4|4|4|3|3|4|3.67|2|4|4|4|4|4|3.67|0|4|4|4|4|3|4|4|3.67|8.99|5|3|4|5|4.25|5|4|4|5|4.5|-5.56|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|3|3|3|2|2|2|50|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|45.5||2|2|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|Black||42|28273|Masters Degree|Divorced|Business: Marketing||1|6|Michael Baisden|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|502181148|31|0|2|502184470|31|0|2|500454904|2||500004772||4|1|500000294, 500004640, 500004901|500000294|-2|500000294|-2|7016|11|||11146|1|||1|450500|134611|4|3|45
500186955|BBBS of Greater Charlotte|Main Office|C|Completed|2004-05-21|2014-02-19|Followup|2013-05-21|2013-05-21|Complete|Done|4|3|4|3|4|4|3.67|||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Lost contact with child/agency|117||1|1|1|1|F|Black||18|No|Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||55|28226|||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|2|500189726|1|0|2|500037840|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|450789||4|3|45
502896719|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-01|2015-08-19|Followup|2013-06-01|2013-06-25|Complete|Done|3|2|3||4|4||4|1|2|1||4|||2|4|4|3|3|4|3.33|2|4|4|2|1|4|2.83|17.67|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|4|5|5|4.75|5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|4|4|4|4|-8.25|3|4|3.5|2|3|2.5|40|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Moved|38.6||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|F|White||27|28269|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|502898127|31|0|2|502959645|1|0|2|500614239|2||-2||4|2|||-2||-2|0|10|||46|2|||1|451498|411397|4|3|45
502997211|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-01|2013-09-05|Followup|2013-06-01|2013-08-16|Expired|Late||||||||3|1|3|4|4|4|3.17|||||||||1|3|3|3|2|4|2.67||||||4|4|3|3.67|||||||3|3|2|2|2.5||||||||||4|1|4|4|3|4|4|3.43||||||4|3|4|3.67|||||1|2|1.5||||2|2||||4|4||Yellow||Child/Family: Feels incompatible with volunteer|15.1||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|F|White||27|28105|Some College||Student: College||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011349|502998689|31|0|2|502926434|1|0|2|500614826|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|451803|438072|4|0|45
502485856|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-02|2013-08-20|Followup|2013-06-02|2013-06-07|Declined|Done|4|||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Moved|26.6||2|2|1|1|F|Hispanic|Other South American|13|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Hispanic||63|28227|Bachelors Degree|Married|Education: Teacher||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|502486303|3|15|2|502253272|3|0|2|500537140|2||-2||4|2|||-2||-2|0|10|||7462|13|||1|453118||4|1|45
502972004|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-29|2012-11-15|Baseline|2012-06-04|2012-06-29|Complete|Done|3|3|3|2|3|4|3|||||||||4|3|3|2|3|4|3.17|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|4.6||1|1|1|1|F|Black||15|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||57|28273|Masters Degree|Single|Business|28210|5|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500001281|502973441|31|0|2|502908172|31|0|2|500617689|2||-2||4|3|||-2||-2|7294|13|||7462|13|||1|453294|-1|4|3|44
502589865|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-29|Followup|2013-06-30|2013-08-08|Complete|Done|3|4|3|1|4|3|3|1|4|2|3|1|1|2|50|4|4|4|2|2|4|3.33|3|1|3|4|4|4|3.17|5.05|4|4|4|4|4|4|4|4|0|3|3|4|3|3.25|5|5|5|5|5|-35|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|3|3.33|20.12|4|3|3.5|1|1|1|250|2|2|2|2|0|4|4|4|4|0|Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|52||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Black||40|28037|Bachelors Degree|Married|Medical: Doctor, Provider||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502590381|31|0|1|502625828|31|0|1|500544108|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|454126|291589|4|3|45
503005868|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-24|2017-02-26|Baseline|2012-06-06|2012-07-20|Complete|Done|2|2|2|1|2|3|2|||||||||2|2|3|2|2|3|2.33|||||||||4|4|4|4||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child: Lost interest|55.1||1|1|1|1|M|Multi-race (Black & Hispanic)||15||Mother|28270|One Parent: Female|$25,000 to $29,999|Y|No||Therapist/Counselor|General Community||Match Support|M|White||51|28173|Bachelors Degree|Married|Consultant|28173|1|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020753|503007379|38|0|1|502935610|1|0|1|500623124|2||-2||4|3|||-2||-2|0|5|||7671|13|||1|456253|-1|4|3|44
500740295|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2013-06-12|2013-06-05|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Volunteer: Feels incompatible with child/family|85||1|1|1|1|M|Black||18||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|White||55|28216|Bachelors Degree|Divorced|Tech: Engineer||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500794907|1|0|1|500179696|2||-2||4|2|||-2||-2|0|5|||46|2|||1|456291||4|3|45
500740293|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2013-06-12|2013-06-05|Complete|Done|4|4|4|2|3|3|3.33|||||||||4|4|4|1|2|4|3.17|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||1|1||||4|4||||Yellow||Child: Lost interest|85||1|1|1|1|M|Black||19||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|Black||39|28216||Single|Transport: Pilot||3|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500876177|31|0|1|500179697|2||-2||4|2|||-2||-2|0|5|||6450|12|||1|456295||4|3|45
502270499|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-25|NaT|Followup|2013-05-25|2013-06-25|Complete|Done|4|3|3|2|3|4|3.17|4|2|1|1|3|4|2.5|26.8|4|4|4|4|4|4|4|2|4|4|2|1|3|2.67|49.81|4|4|4|4|4|4|4|4|0|4|4|5|4|4.25|3|4|3|4|3.5|21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|3|3|3|4|4|4|-25|2|2|2|2|0|4|4||||Green|Amachi||69.7||2|2|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||34|28203|Masters Degree|Single|Business: Mgt, Admin|28273|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502231230|31|0|2|502510107|1|0|2|500536754|2||500003586||2|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|456380|218599|4|3|45
503013779|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-10|2013-08-14|Baseline|2012-06-07|2012-07-10|Complete|Done|3|2|2|3|2|3|2.5|||||||||1|2|3|1|1|2|1.67|||||||||3|3|3|3||||||2|2|2|3|2.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Time constraint|13.1||2|2|1|1|F|Multi-race (Black & White)||17|No|Mother|28134|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|Asian||30|28270|Bachelors Degree|Married|Education|28211|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|503724588|36|0|2|502993965|4|0|2|500618402|2||-2||4|3|||-2||-2|0|10|||7462|13|||1|456670|-1|4|3|44
502908460|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-07|2014-09-04|Followup|2013-06-07|2013-06-07|Complete|Done|4|2|3|2|2|3|2.67|4|4|1|3|4|4|3.33|-19.82|3|3|4|4|4|4|3.67|2|2|2|2|1|3|2|83.5|4|4|4|4|4|2|2|2.67|49.81|5|4|4|4|4.25|1|5|3|3|3|41.67|4|4|4|4|4|4|4|4|4|4|4|4|3|4|2|3.57|12.04|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|1|2.5|60|2|2|1|1|100|2|2|4|4|-50|Yellow||Volunteer: Lost contact with child/agency|26.9||1|1|1|1|F|Hispanic||18|No|Mother|28227|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||40|28079|Bachelors Degree|Single|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502909871|3|0|2|502938939|1|0|2|500616222|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|456864|434253|4|3|45
502527168|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-19|2016-08-29|Baseline|2012-06-07|2012-06-19|Complete|Done|2|4|3|3|3|3|3|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|4|3.33||||||4|3|3.5|||||2|2||||4|4||||Red||Child: Graduated|50.3||1|1|2|2|M|Hispanic|Mexican|19|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502527621|3|10|1|501646021|3|0|1|500618440|2||-2||4|3||500005291|-2||-2|2203|12|||7464|9|||1|456875|-1|4|3|44
501765404|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-20|2013-08-29|Followup|2013-04-20|2013-04-30|Complete|Done|3|4|4|1|3|3|3|3|3|3|1|4|3|2.83|6.01|3|3|3|4|4|4|3.5|2|3|3|2|3|3|2.67|31.09|4|4|4|4|4|4|4|4|0|4|3|3|3|3.25|3|5|5|4|4.25|-23.53|4|4|4|4|4|4|4|4|4|4|4|3|2|3|1|3|33.33|4|4|4|4|4|3|4|3.67|8.99|4|4|4|4|3|3.5|14.29|2|2|1|1|100|4|4||||Yellow||Volunteer: Lost contact with child/agency|40.3||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Multi-race (Black & White)||28|28262||Single|Student: College|28262|3|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500011746|501765751|31|0|1|501958658|36|0|1|500443642|2||-2||4|2|||-2||-2|0|10|||9221|5|||1|457381|36416|4|3|45
503021552|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-19|2015-10-22|Baseline|2012-06-08|2012-06-18|Complete|Done|3|1|1|4|3|4|2.67|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4||||||||||||4|4|3|3.67||||||2|3|2.5|||||2|2||||4|4||||Yellow||Volunteer: Moved|40.1||1|1|1|1|F|Black||14|No|Mother|28270|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Multi-Race (None of the above)||28|28215|Some College|Single|Insurance||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503023091|31|0|2|502951522|7|0|2|500618601|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|457665|-1|4|3|44
502008563|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-02|2013-07-29|Followup|2013-06-02|2013-06-24|Complete|Done|3|2|3|1|3|4|2.67|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Moved|37.9||2|2|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||31|28210|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502008962|31|0|1|502053340|1|0|1|500453826|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|457686||4|3|45
501142903|BBBS of Greater Charlotte|Main Office|C|Active|2008-06-05|NaT|Followup|2013-06-05|2013-06-11|Complete|Done|4|2|4|4|4|4|3.67|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||105.3||1|1|1|1|M|Black||14|Yes|GrandMother|28208|One Parent: Female|Less than $10,000||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|M|White||53|28204|Juris Doctorate (JD)|Married|Law: Lawyer|28244|16|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501143177|31|0|1|501236825|1|0|1|500268808|2||500003586||2|1|500000294|500000294|-2|500000294|-2|7294|13|||2238|7|||1|457775||4|3|45
501755470|BBBS of Greater Charlotte|Main Office|C|Active|2010-06-30|NaT|Followup|2012-06-30|2012-07-24|Complete|Done|4|1|4|1|4|4|3|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||5|5|2|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||80.5||2|2|2|2|F|Black||13|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|501755813|31|0|2|502038804|31|0|2|500456645|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|457881||4|3|45
502102857|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-25|2013-06-18|Followup|2013-03-25|2013-06-09|Expired|Late||||||||4|4|3|1|4|4|3.33|||||||||3|4|3|3|1|4|3||||||4|4|2|3.33|||||||4|4|5|1|3.5||||||||||4|4|4|4|2|4|3|3.57||||||4|4|4|4|||||3|2|2.5||||2|2|||||||Red|2010-2012 OJJDP JJI|Volunteer: Moved|26.8||2|2|1|1|M|Black||18|No|Mother|28278|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||38|28273|Bachelors Degree|Married|Insurance|28202|2|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502103284|31|0|1|502464465|31|0|1|500526162|2||-2||4|3|500005291|500005291|-2|500000294, 500004640|-2|0|4|||7446|3|||1|457934|40474|4|0|45
500968246|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-29|2015-04-30|Followup|2014-04-29|2014-06-12|Complete|Done|3|2|4|2|3|4|3|||||||||2|4|3|3|3|3|3|||||||||4|4|3|3.67||||||1|2|4|4|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|84||1|1|1|1|M|Black||19|No|Aunt|28269|One Parent: Female|$10,000 to $14,999|Y|No||Therapist/Counselor|General Community||Match Support|M|Black||35|28213|Bachelors Degree|Single|Business: Sales||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500968516|31|0|1|501179573|31|0|1|500251681|2||-2||4|1|||-2||-2|0|5|||46|2|||1|458058||4|3|45
500186645|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-03|2016-01-06|Followup|2013-06-03|2013-07-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|139.1||1|1|1|1|M|Black||18|Yes|Mother|28208|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28256|High School Graduate|Married|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500018987|500188043|31|0|1|500189545|31|0|2|500037636|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|458067||4|1|45
501253965|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-11|2016-05-17|Followup|2013-06-11|2013-07-22|Complete|Done|4|4|4|1|4|4|3.5|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||3|4|2|3|3|||||||4|1|4|4|3|4|4|3.43||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Time constraint|47.2||3|3|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|Y|No||Self|General Community|Amachi|Enrollment|F|Black||34|28215|Some College|Single|Customer Service||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503287812|31|0|2|502985911|31|0|2|500613577|2||-2||4|1||500000294|-2||-2|0|10|||7464|9|||1|458764||4|3|45
502551092|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-20|2015-10-29|Followup|2013-05-20|2013-06-07|Declined|Done||||||||3|3|4|1|4|4|3.17|||||||||2|4|3|1|2|4|2.67||||||4|4|4|4|||||||3|4|5|3|3.75||||||||||4|4|4|4|4|4|2|3.71||||||3|4|4|3.67|||||4|2|3||||1|1||||4|4||Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|53.3||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||42|28210||Single|Business: Human Resources||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|502551545|31|0|2|502366844|1|0|2|500536172|2||-2||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||10326|3|460|3|1|458827|280274|4|1|45
502173445|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-23|2013-09-26|Followup|2013-05-23|2013-07-08|Declined|Late||||||||4|4|4|3|4|4|3.83|||||||||2|4|3|3|4|3|3.17||||||4|3|4|3.67|||||||5|4|4|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|3|3.5||||2|2|||||||Red|Amachi|Volunteer: Lost contact with child/agency|28.2||1|1|1|1|F|Black||19|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Service Organization|General Community|Amachi|Match Support|F|White||28|28206|Bachelors Degree|Single|Education: Teacher||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502173869|31|0|2|502266833|1|0|2|500532710|2||500003586||4|3|500000294|500000294|-2||-2|0|11|||7464|9|||1|459164|270032|4|1|45
500186702|BBBS of Greater Charlotte|Main Office|C|Completed|2004-04-28|2014-11-25|Followup|2013-04-28|2013-04-24|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|1|4|3.5|||||||||4|4|4|4||||||3|5|3|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|126.9||1|2|1|2|F|Black||20|Yes|GrandMother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||57|28212|Some College|Married|Unknown||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|RTBM|277|60|598|500000170|500017732|500188150|31|0|2|500189528|31|0|2|500038225|2||500003586||4|1|500000294|500000294|-2|500015184|-1|0|10|||7462|13|||1|459488||4|3|45
502990571|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-25|2013-05-21|Baseline|2012-06-13|2012-06-25|Complete|Done|3|3|2|1|2|1|2|||||||||3|3|4|3|4|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Yellow||Volunteer: Time constraint|10.8||2|2|1|1|F|Multi-race (Black & Hispanic)||15|Yes|Mother|28217|Two Parent|$35,000 to $39,999||Yes||Self|General Community||Match Support|F|Black||29|28217|Bachelors Degree|Single|Business||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502992028|38|0|2|503004889|31|0|2|500619186|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|460382|-1|4|3|44
502566108|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-24|2014-09-08|Followup|2013-05-24|2013-06-13|Complete|Done|4|1|2|1|2|3|2.17|3|2|4|1|3|4|2.83|-23.32|2|3|4|3|3|3|3|2|3|3|2|2|3|2.5|20|4|3|3|3.33|4|3|4|3.67|-9.26|4|4|4|4|4|4|1|4|4|3.25|23.08|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|1|1|1|1|4|3|4|3.67|-72.75|4|4|4|3|4|3.5|14.29|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|39.5||1|1|1|1|F|Hispanic||17|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||33|28209||Single|Student: College||0|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502566562|3|0|2|502562271|1|0|2|500535933|2||-2||4|1|500005291|500005291|-2|500005291|-2|0|4|||7464|9|||1|460594|279328|4|3|45
502866443|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-14|2014-09-23|Followup|2013-06-14|2013-06-30|Complete|Done|3|1|2|1|3|3|2.17|4|1|2|1|3|4|2.5|-13.2|2|3|3|2|2|3|2.5|1|3|3|1|2|4|2.33|7.3|4|4|4|4|4|2|4|3.33|20.12|3|3|4|3|3.25|5|3|5|4|4.25|-23.53|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|4|3.67|4|4|4|4|-8.25|3|4|3.5|4|1|2.5|40|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|27.3||1|1|1|1|F|Black||14|No|Mother|28262|One Parent: Female|$30,000 to $34,999|Y|No||Self|General Community||Match Support|F|Black||38|28212|Some College|Single|Business: Mgt, Admin|28270|7|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502867844|31|0|2|502920462|31|0|2|500613414|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|461081|432716|4|3|45
500545470|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-01-25|Followup|2013-04-30|2013-06-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|104.9||1|1|1|1|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||34|29708|Bachelors Degree|Single|Self-Employed, Entrepreneur|29708|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501750989|31|0|1|500815012|1|0|1|500173957|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|3|||2238|7|||1|461486||4|1|45
502700505|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-27|NaT|Baseline|2012-06-15|2012-06-27|Complete|Done|4|3|3|3|4|4|3.5|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|2|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||3|3||||||||3|3|3|||||2|2||||4|4||||Green|||56.6||1|1|1|1|M|Black||17|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Black||41|28210|Bachelors Degree|Separated|Arts, Entertainment, Sports|28202|2|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502701350|31|0|1|503029324|31|0|1|500619505|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|461562|-1|4|3|44
502477677|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-29|2013-08-22|Followup|2012-07-29|2012-07-23|Complete|Done|3|2|2|2|3|3|2.5|||||||||1|4|4|1|1|3|2.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||3|3||||Red||Volunteer: Lost contact with child/agency|24.8||1|1|1|1|M|Black||13|No|Mother|28273|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||31|28217|Bachelors Degree|Single|Business: Engineer|28273|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|502478124|31|0|1|502621765|31|0|1|500545314|2||-2||4|3|||-2||-2|0|5|||7496|10|||1|461950||4|3|45
501722052|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-11|2015-01-30|Followup|2013-05-11|2013-06-05|Complete|Done|3|1|2|2|2|3|2.17|||||||||2|3|4|2|4|3|3|||||||||3|4|4|3.67||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|2|2|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|56.7||2|2|1|1|F|White||13|Yes|GrandMother|28083|Grandparents|Unknown||No||Self|General Community||Enrollment|F|White||40|28027||Single|Customer Service|28027|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501227925|1|0|2|502030533|1|0|2|500450450|2||-2||4|1|500000294||-2||-2|0|10|||7464|9|12|3|1|462346||4|3|45
502435258|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-12|2014-10-30|Followup|2013-01-12|2013-01-08|Complete|Done|4|4|4|4|4|4|4|||||||||1|3|2|2|1|3|2|||||||||3|3|3|3||||||2|5|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|33.6||2|2|1|1|F|Black||13|No|Relative: Other|28081|Other Relative|Unknown|Y|Yes||Self|General Community||Enrollment|F|Black||31|28025|Bachelors Degree|Single|Child/Day Care Worker|28027|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|502435701|31|0|2|502670193|31|0|2|500589905|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|462432||4|3|45
501626226|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-30|2017-03-14|Followup|2013-06-30|2013-06-25|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|80.5||2|2|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||33|28203|High School Graduate|Single|Retail: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501622822|31|0|2|502036832|1|0|2|500457771|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|462595||4|3|45
500896018|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-03|2014-08-14|Followup|2013-07-03|2013-07-08|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|2|2.67||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|73.4||1|1|1|1|F|Black||20|Yes|Mother|28027|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||40|28027|Bachelors Degree|Separated|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500896288|31|0|2|501225232|31|0|2|500269506|2||-2||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|462687||4|3|45
500271303|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-30|2015-08-03|Followup|2013-04-30|2013-04-30|Complete|Done|4|4|4|4|4|4|4|||||||||1|4|4|1|1|3|2.33|||||||||4|4|4|4||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|75.1||2|2|1|1|F|Black||17|Yes|Mother|28227|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|White||31|28204|Bachelors Degree|Single|Business: Engineer|28269|0|2|TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500271368|31|0|2|501291358|1|0|2|500354049|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||130|1|||1|462743||4|3|45
501597169|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-06|2016-05-31|Followup|2013-04-06|2013-03-27|Complete|Done|4|3|4|2|4|4|3.5|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|2|3||||||4|4|4|||||2|2||||4|4||||Green||Agency: Challenges with program/partnership|85.8||1|1|1|1|M|Black||13||Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||54|28262|High School Graduate|Married|Disabled||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501597489|31|0|1|501563612|31|0|1|500352827|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|462984||4|3|45
500378354|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-01|NaT|Followup|2013-05-01|2013-04-29|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||106.5||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$40,000 to $44,999||No|Big|Neighbor/Friend|General Community||Match Support|M|White||36|28270|Juris Doctorate (JD)|Married|Law: Lawyer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500378596|31|0|1|501181060|1|0|1|500264206|2||-2||2|1|||-2||-2|6854|8|||46|2|||1|463257||4|3|45
502527168|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-19|2016-08-29|Followup|2013-06-19|2013-06-24|Complete|Done|3|2|3|2|3|3|2.67|2|4|3|3|3|3|3|-11|2|2|3|3|1|4|2.5|2|4|3|2|3|3|2.83|-11.66|4|4|4|4|4|4|4|4|0|4|4|3|3|3.5|4|4|3|4|3.75|-6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3|4|3.33|20.12|3|4|3.5|4|3|3.5|0|2|2|2|2|0|4|4|4|4|0|Red||Child: Graduated|50.3||1|1|2|2|M|Hispanic|Mexican|19|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502527621|3|10|1|501646021|3|0|1|500618440|2||-2||4|3||500005291|-2||-2|2203|12|||7464|9|||1|463362|456875|4|3|45
502570396|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-08|Followup|2013-06-30|2013-07-15|Complete|Done|4|3|1|2|4|4|3|3|4|4|4|4|4|3.83|-21.67|2|3|3|3|3|2|2.67|4|4|3|4|2|3|3.33|-19.82|3|3|3|3|4|4|4|4|-25|3|2|3|3|2.75|3|5|3|3|3.5|-21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|1|3|2|100|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|51.3||1|1|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28078|Bachelors Degree|Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018987|502570850|38|0|2|502545897|31|0|2|500539251|2||-2||4|1|500005291|500005291|-2||-2|34|2|||46|2|||1|463458|296321|4|3|45
502980958|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-17|NaT|Baseline|2012-06-19|2012-07-17|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|3|3|3|3|3|3|||||||||4|3|4|3.67||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||56||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Sales|28273|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502982410|31|0|1|503008664|1|0|1|500620394|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|463519|-1|4|3|44
503021552|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-19|2015-10-22|Followup|2013-06-19|2013-08-02|Declined|Done||||||||3|1|1|4|3|4|2.67|||||||||2|4|4|4|2|4|3.33||||||4|4|4|4|||||||3|4|3|4|3.5||||||||||4|4|4|4|4|4||||||||4|4|3|3.67|||||2|3|2.5||||2|2||||4|4||Yellow||Volunteer: Moved|40.1||1|1|1|1|F|Black||14|No|Mother|28270|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Multi-Race (None of the above)||28|28215|Some College|Single|Insurance||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503023091|31|0|2|502951522|7|0|2|500618601|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|463634|457665|4|1|45
501212047|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-07|NaT|Followup|2013-05-07|2013-05-14|Complete|Done|4|3|3|2|4|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||106.3||1|1|1|1|F|White||18|No|Father|28207|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||33|28226||Single|Human Services: Non-Profit|28205|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501212321|1|0|2|501242250|1|0|2|500264889|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|463668||4|3|45
501213488|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-19|NaT|Followup|2013-05-19|2013-06-17|Complete|Done|4|3|4|3|4|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||105.9||1|1|1|1|F|White||14|No|Father|28207|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Finance: Banking|28255|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|501213764|1|0|2|501225276|1|0|2|500262655|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|463669||4|3|45
502513881|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-21|2014-09-22|Followup|2013-06-21|2013-06-24|Complete|Done|3|2|2|1|4|3|2.5|||||||||2|2|4|3|3|3|2.83|||||||||3|3|3|3||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|2|3|2.67||||||4|3|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|27||2|2|3|3|F|Hispanic||14|No|Mother|28262|One Parent: Female|Unknown||No||School|General Community||Enrollment|F|Black||49|28213|Juris Doctorate (JD)|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502514330|3|0|2|502393006|31|0|2|500615307|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|464296||4|3|45
502863781|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-31|2015-01-30|Baseline|2012-06-22|2012-07-31|Complete|Done|3|4|3|2|3|4|3.17|||||||||2|4|3|2|1|2|2.33|||||||||4|4|4|4||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Red||Volunteer: Time constraint|30||1|1|1|1|M|Black||18|No|Mother|28031|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|M|White||26|28031|High School Graduate|Single|Personal Trainer/Coach|28117|0|4|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502865175|31|0|1|503002010|1|0|1|500621061|2||-2||4|3|||-2||-2|0|10|||17161|11|||1|465050|-1|4|3|44
502853025|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-11|2013-05-28|Baseline|2012-06-25|2012-07-09|Complete|Done|2|3|4|3|2|3|2.83|||||||||2|2|4|4|3|4|3.17|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|4|3|||||1|1||||4|4||||Green||Child: Lost interest|10.5||1|1|1|1|F|Hispanic|Mexican|17|No|Mother|28205|Two Parent|Unknown|Y|Yes||School|General Community||Match Support|F|Hispanic||40|28277|Some College|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502854420|3|10|2|503009880|3|0|2|500621608|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|465941|-1|4|3|44
502530688|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-25|2016-05-20|Followup|2013-06-25|2013-07-24|Complete|Done|3|3|4|1|4|4|3.17|4|3|2|2|4|4|3.17|0|2|3|3|2|3|2|2.5|3|4|4|2|3|4|3.33|-24.92|4|4|4|4|4|4|4|4|0|3|3|3|4|3.25|3|2|4|3|3|8.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|2|1|1.5|2|2|2|-25|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Time constraint|46.8||2|2|3|3|M|Black||17||Mother|28210|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28277|Bachelors Degree|Married|Business||0|0|Michael Baisden|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502531141|31|0|1|502166996|31|0|1|500621632|2||-2||4|2||500005291|-2||-2|0|3|||11272|1|||1|466035|279295|4|3|45
500783100|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-08-29|Followup|2013-04-30|2013-04-30|Declined|Done|4|1|2|||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|112||1|1|1|1|M|Black||16||Mother|28206|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||36|28203|||Retail: Sales|28226|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|500783368|31|0|1|500777047|1|0|1|500174449|2||-2||4|2|||-2||-2|0|10|||46|2|||1|466271||4|1|45
501721761|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-25|2015-07-27|Followup|2013-06-25|2013-07-22|Complete|Done|3|4|1|1|2|4|2.5|||||||||2|3|2|2|4|3|2.67|||||||||3|4|3|3.33||||||4|3|2|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|37||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|M|White||31|28210|Bachelors Degree|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501722098|31|0|1|503023854|1|0|1|500618753|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|466285||4|3|45
502569117|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-31|NaT|Followup|2013-05-31|2013-07-25|Declined|Late||||||||4|2|4|1|3|4|3|||||||||2|4|4|3|4|4|3.5||||||4|4|4|4|||||||5|4|5|3|4.25||||||||||4|4|4|4|4|4|3|3.86||||||4|3|2|3|||||2|2|2||||1|1||||4|4||Green|Amachi, 2010-2012 OJJDP JJI||69.5||1|1|1|1|F|Black||15|Yes|Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||40|28269|Masters Degree|Single|Tech: Engineer|77058|6|6|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500017732|502569571|31|0|2|502538689|31|0|2|500536957|2||500003586||2|1|500000294, 500005291|500005291|-2||-2|0|10|||17161|11|||1|466855|284793|4|1|45
502700505|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-27|NaT|Followup|2013-06-27|2013-06-25|Complete|Done|1|4|4|4|4|4|3.5|4|3|3|3|4|4|3.5|0|3|4|3|4|3|4|3.5|2|3|3|2|2|3|2.5|40|4|4|4|4|4|4|4|4|0|4|3|2|5|3.5|3|2|2|3|2.5|40|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3||||3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Green|||56.6||1|1|1|1|M|Black||17|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Black||41|28210|Bachelors Degree|Separated|Arts, Entertainment, Sports|28202|2|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502701350|31|0|1|503029324|31|0|1|500619505|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|467339|461562|4|3|45
502137546|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2015-10-20|Followup|2013-04-29|2013-04-30|Complete|Done|4|3|3|1|3|3|2.83|4|4|2|2|4|4|3.33|-15.02|4|4|4|4|4|4|4|2|4|3|2|2|3|2.67|49.81|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|5|4|4|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|3|4|3.5|14.29|2|2|2|2|0|4|4||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|53.7||1|2|1|2|F|Black||16||Mother|28213|Other/Unknown|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28262|||Business: Mgt, Admin|75234|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502137975|31|0|2|501641708|31|0|2|500520728|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|467587|36419|4|3|45
502552443|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-08|2014-12-30|Followup|2013-06-08|2013-06-07|Complete|Done|4|2|3|2|3|3|2.83|4|4|4|2|3|4|3.5|-19.14|2|3|3|3|4|3|3|4|4|4|4|2|4|3.67|-18.26|4|4|4|4|4|4|4|4|0|4|5|4|4|4.25|5|4|4|5|4.5|-5.56|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|4|4|3|4|3|3.33|20.12|4|3|3.5|2|2|2|75|2|2||||4|4||||Green|Project Big|Child: Graduated|42.7||1|1|1|1|F|Multi-race (Black & Hispanic)||20|No|GrandMother|28208|Grandparents|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28209|Bachelors Degree|Single|Medical|28209|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502552891|38|0|2|502471967|1|0|2|500537261|2||-2||4|1|500004640|500004640, 500005291|-2||-2|0|4|||7496|10|||1|467606|286064|4|3|45
502183053|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-28|NaT|Followup|2013-06-28|2013-06-18|Complete|Done|3|1|2|1|1|4|2|3|1|2|1|1|2|1.67|19.76|4|4|4|2|4|4|3.67|4|2|4|2|3|4|3.17|15.77|4|4|4|4|4|4|3|3.67|8.99|4|5|5|4|4.5|4|4|4|4|4|12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|4|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Green|||56.6||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||46|28134|Bachelors Degree|Married|Finance|28105|1|6|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|502183482|31|0|1|503073638|31|0|1|500621039|2||-2||2|1|||-2|500014681|-2|0|10|||4748|14|633|1|1|467899|414734|4|3|45
501662021|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-14|2014-02-21|Baseline|2012-06-28|2012-08-14|Complete|Done|3|1|4|1|1|3|2.17|||||||||2|4|4|4|4|3|3.5|||||||||4|4|3|3.67||||||5|4|3|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|1|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|18.3||2|2|1|1|M|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|Black||50|28269|Some College|Divorced|Retired||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500011349|501090456|31|0|1|502902255|31|0|1|500627357|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|468082|-1|4|3|44
502185074|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-12|2016-08-02|Followup|2013-05-12|2013-07-10|Declined|Late||||||||1|2|1|4|1|1|1.67|||||||||3|1|3|1|1|1|1.67||||||4|4|4|4|||||||3|2|4|5|3.5||||||||||4|4|4|4|4|4|4|4||||||2|3|2|2.33|||||2|2|2||||2|2|||||||Green|2010-2012 OJJDP JJI|Child: Graduated|62.7||2|2|1|1|F|Black||18|No|GrandMother|28208|Grandparents|Unknown||Yes|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||68|28262|Bachelors Degree|Living w/ Significant Other|Business: Clerical||2|0|Relative|Relative|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017732|502185503|31|0|2|502490418|31|0|2|500533846|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|5635|9|||17161|11|||1|468476|159621|4|1|45
502537477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-12|2016-07-14|Followup|2013-05-12|2013-07-10|Declined|Late||||||||3|2|1|1|3|3|2.17|||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||3|5|4|4|4||||||||||4|4|4|4|3|4|3|3.71||||||2|3|2|2.33|||||2|4|3||||2|2||||4|4||Green|Project Big, 2010-2012 OJJDP JJI|Child: Graduated|62.1||1|1|3|4|F|Black||19||Mother|28208|Two Parent|$15,000 to $19,999||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||48|28214|Bachelors Degree|Single|Tech: Management|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Project Big|Enrollment|277|60|598|500000170|500017732|502537922|31|0|2|500189507|31|0|2|500535475|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2|500000294, 500004640|-2|0|4|||2238|7|||1|468477|277756|4|1|45
502920377|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-29|2017-02-28|Followup|2013-06-29|2013-08-24|Declined|Late||||||||3|2|2|2|2|3|2.33|||||||||2|3|2|3|3|3|2.67||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||3||||||2|2||||4|4||Green||Volunteer: Lost contact with child/agency|56||1|1|1|1|F|Black||14|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||31|28211|Bachelors Degree|Single|Real Estate: Realtor|19137|2|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502921794|31|0|2|502942994|1|0|2|500620441|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|468652|439883|4|1|45
502506397|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-30|2016-11-01|Followup|2013-06-30|2013-07-22|Complete|Done|2|2|3|1|3|4|2.5|2|1|2|2|3|3|2.17|15.21|2|3|4|3|2|3|2.83|3|3|4|3|2|4|3.17|-10.73|3|2|2|2.33|3|2|2|2.33|0|4|3|3|2|3|5|4|3|2|3.5|-14.29|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|1|2|1|1.33|1|3|3|2.33|-42.92|1|3|2|2|4|3|-33.33|2|2|1|1|100|4|4|4|4|0|Yellow||Child: Severity of challenges|52.1||1|1|1|1|F|White||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||33|28277|Bachelors Degree|Single|Consultant|28202|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502506846|1|0|2|503039829|1|0|2|500619509|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|469118|407242|4|3|45
501157075|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-30|2016-01-21|Followup|2013-06-30|2013-07-22|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|3|3|2|3|3|||||||||4|4|4|4||||||4|3|2|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child: Lost interest|42.7||3|4|1|1|F|Black||17||Relative: Other|28206|Grandparents|Unknown||Yes||School|General Community|Amachi|Match Support|F|Black||37|28215|Masters Degree|Single|Human Services: Social Worker||2|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020752|501157349|31|0|2|502978065|31|0|2|500619009|2||-2||4|2||500000294|-2||-2|0|4|||7464|9|||1|469129||4|3|45
502402515|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-17|2015-12-28|Followup|2013-05-17|2013-06-05|Complete|Done|3|1|4|1|3|4|2.67|3|1|3|1|1|4|2.17|23.04|2|4|3|3|3|3|3|1|4|3|1|3|4|2.67|12.36|4|4|4|4|4|4|4|4|0|3|2|2|2|2.25|3|2|2|2|2.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|3|4|3.5|4|3|3.5|0|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|55.4||1|1|1|1|M|Black||16|No|Mother|28215|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28215||Single|Law: Police Officer||14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502402953|31|0|1|502537081|31|0|1|500535130|2||-2||4|1|500005291|500005291|-2||-2|34|2|||7464|9|||1|469331|276236|4|3|45
502549830|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-30|NaT|Followup|2013-06-30|2013-07-14|Complete|Done|1|2|4|1|4|3|2.5|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|2|2|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||68.5||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|Amachi, Project Big, Project Big AND Amachi|Match Support|M|Black||25|28211||Single|Transport: Driver||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|1|502462453|31|0|1|500538768|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-1||-2|0|4|||7464|9|||1|469429||4|3|45
502549829|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-30|NaT|Followup|2013-06-30|2013-06-24|Complete|Done|3|4|4|4|1|1|2.83|3|1|2|1|2|2|1.83|54.64|1|3|2|1|1|2|1.67|2|3|2|2|2|2|2.17|-23.04|4|4|4|4|3|2|2|2.33|71.67|2|2|3|3|2.5|3|2|2|3|2.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|2|2|1|1|100|4|4||||Green|Amachi, Project Big, Project Big AND Amachi||68.5||1|1|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|Amachi, PERL 2014-2016, Project Big, Project Big AND Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Business: Engineer|30357|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|1|502594393|31|0|1|500541795|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901, 500014681|-1||-2|0|4|||7464|9|||1|469436|283404|4|3|45
501129794|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-14|2015-10-29|Followup|2013-06-14|2013-07-14|Complete|Done|4|1|2|1|3|3|2.33|||||||||3|3|3|2|3|4|3|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|52.5||1|2|1|2|M|Black||14||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|F|Black||45|28273|Masters Degree|Single|Tech: Research/Design||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500017777|501130068|31|0|1|500922570|31|0|2|500540937|2||-2||4|1|||-2||-2|0|4|||46|2|||1|469573||4|3|45
502045258|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-25|2016-08-29|Followup|2013-06-25|2013-08-08|Complete|Done|3|3|3|3|3|3|3|4|2|4|1|4|4|3.17|-5.36|3|4|4|3|3|3|3.33|4|4|4|4|4|4|4|-16.75|4|4|4|4|4|4|4|4|0|5|3|4|4|4|5|5|5|5|5|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|4|3|3.5|4|3|3.5|0|2|2|2|2|0|4|4||||Green||Volunteer: Lost contact with child/agency|74.2||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28262|Bachelors Degree|Single|Medical: Nurse|28262|4|9|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502190790|31|0|2|500457916|2||-2||4|1|||-2||-2|0|10|||6247|12|||1|469584|148107|4|3|45
502590651|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2013-08-22|Followup|2013-06-30|2013-08-08|Declined|Done||||||||4|3|4|2|4|4|3.5|||||||||2|4|3|1|2|4|2.67||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||4|3|3.5||||1|1||||4|4||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Time constraint|25.8||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||36|28205|Bachelors Degree|Single|Business: Marketing|28117|7|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011746|502591168|31|0|2|502589724|1|0|2|500542166|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|469598|294373|4|1|45
502570185|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2014-05-15|Followup|2013-06-30|2013-08-28|Complete|Late|4|4|2|2|2|3|2.83|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|34.5||1|1|1|1|F|Black||14|No|Mother|28206|Other/Unknown|Unknown||Yes||Relative|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||58|28226|Masters Degree|Single|Tech: Management|28078|0|2|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|277|60|598|500000170|500017777|502570639|31|0|2|502191626|31|0|2|500542078|2||500004641||4|2|500000294, 500004640, 500004901, 500005291|500004640, 500005291|-2|500004640|-2|0|3|459|3|46|2|||1|470146||4|3|45
502802219|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-30|2014-02-27|Baseline|2012-07-06|2012-07-27|Complete|Done|3|1|1|1|2|2|1.67|||||||||3|4|4|3|2|4|3.33|||||||||3|3|2|2.67||||||4|4|4|4|4|||||||4|4|4|4|4|4|2|3.71||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|19||1|1|1|1|M|White||17|No|Mother|28209|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|M|White||35|28212|Some College|Single|Tech: Computer/Programmer|28212|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502803493|1|0|1|503060158|1|0|1|500623104|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|470627|-1|4|3|44
502605248|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-07|2014-02-27|Baseline|2012-07-06|2012-08-07|Complete|Done|2|2|3|2|2|3|2.33|||||||||2|4|1|4|2|3|2.67|||||||||4|4|4|4||||||4|2|5|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|18.7||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|Unknown||Yes||Relative|General Community|Project Big|Enrollment|M|White||36|28205|Masters Degree|Single|Finance: Banking||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502137975|31|0|1|503049689|1|0|1|500623109|2||-2||4|1||500004640|-2||-2|0|3|||7496|10|||1|470640|-1|4|3|44
502743091|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-18|2014-09-04|Baseline|2012-07-09|2012-07-18|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|3|2|3|3|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4|||||1|1||||4|4||||Yellow||Volunteer: Lost contact with child/agency|25.6||1|1|1|1|M|Black||19|No|Mother|28215|One Parent: Female|$30,000 to $34,999|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||39|28203|Bachelors Degree|Single|Unemployed||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502743998|31|0|1|503079983|1|0|1|500623169|2||-2||4|2||500005291|-2||-2|6854|8|||7496|10|||1|470985|-1|4|3|44
500186952|BBBS of Greater Charlotte|Main Office|C|Active|2004-07-15|NaT|Followup|2013-07-15|2013-07-09|Complete|Done|4|4|2|4|4|4|3.67|||||||||1|2|3|1|2|3|2|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green|Amachi||152||1|1|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||73|28203||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|500188132|31|0|2|500189723|1|0|2|500037836|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|471006||4|3|45
502045254|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-08|2015-10-09|Followup|2013-06-08|2013-06-07|Complete|Done|4|2|2|2|3|3|2.67|2|4|4|4|3|4|3.5|-23.71|1|3|3|2|3|3|2.5|2|4|3|2|2|3|2.67|-6.37|4|4|4|4|4|4|4|4|0|4|4|3|4|3.75|2|4|3|3|3|25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|2|3|33.33|4|4|4|3|3|3|33.33|2|2|1|1|100|3|3||||Yellow||Child: Graduated|64||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502171015|31|0|2|500454926|2||-2||4|2|||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1|471028|134736|4|3|45
501185592|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-23|2016-03-03|Followup|2013-06-23|2013-06-26|Complete|Done|3|4|4|4|4|3|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Family structure changed|92.3|Y|1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||45|28211||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501255830|1|0|1|500270254|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|471081||4|3|45
500186277|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2014-07-16|Followup|2013-07-08|2013-09-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Moved|60.3||3|4|2|3|F|Black||18||Mother|28206|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||39|28210|Bachelors Degree|Married|Business: Sales||8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500187876|31|0|2|500188587|1|0|2|500373187|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|471178||4|0|45
500243491|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-10|NaT|Followup|2013-07-10|2013-07-10|Complete|Done|1|4|4|4|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||56.2||4|4|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|F|Black||47|28269|Bachelors Degree|Single|Law: Paralegal|28202|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188056|31|0|2|502919490|31|0|2|500619145|2||-2||2|1||500000294|-2||-2|0|4|||7464|9|||1|471354||4|3|45
503013779|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-10|2013-08-14|Followup|2013-07-10|2013-08-08|Declined|Done||||||||3|2|2|3|2|3|2.5|||||||||1|2|3|1|1|2|1.67||||||3|3|3|3|||||||2|2|2|3|2.25||||||||||4|4|4|4|4|4|4|4||||||3|3|2|2.67|||||3|3|3||||2|2||||4|4||Red||Volunteer: Time constraint|13.1||2|2|1|1|F|Multi-race (Black & White)||17|No|Mother|28134|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|Asian||30|28270|Bachelors Degree|Married|Education|28211|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500011746|503724588|36|0|2|502993965|4|0|2|500618402|2||-2||4|3|||-2||-2|0|10|||7462|13|||1|471468|456670|4|1|45
502939293|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-24|2013-11-21|Baseline|2012-07-11|2012-09-24|Complete|Done|4|1|4|1|4|4|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|5|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|13.9||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|F|White||48|28269|Bachelors Degree|Single|Finance: Banking||18|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502940718|31|0|2|502855925|1|0|2|500632744|2||-2||4|3|||-2||-2|0|4|||131|1|||1|472079|-1|4|3|44
500408135|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-25|2015-01-30|Followup|2013-05-25|2013-06-30|Complete|Done|3|3|3|3|4|3|3.17|||||||||3|4|3|3|3|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|104.2||1|1|4|4|F|Black||19|Yes|Mother|28083|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500008321|500408385|31|0|2|500189709|31|0|2|500099932|2||500003586||4|1|500000294|500000294|-2|500000294, 500016374|-2|6854|8|||2230|7|||1|472090||4|3|45
502902247|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-11|NaT|Followup|2013-07-11|2013-08-21|Complete|Done|2|2|4|2|3|2|2.5|2|4|4|2||2|||3|4|3|4|4|4|3.67|3|4|3|3|3|3|3.17|15.77|4|4|4|4|4|4|4|4|0|4|5|4|5|4.5|4|5|3|5|4.25|5.88|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|4|3.67|3|4|3|3.33|10.21|3|3|3|3|3|3|0|2|2|1|1|100|4|4|4|4|0|Green|||56.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||30|28203|Bachelors Degree|Single|Business: Marketing|28117|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502903657|31|0|2|502801082|1|0|2|500619356|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|472131|422744|4|3|45
502067798|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-09|NaT|Followup|2013-07-09|2013-07-10|Complete|Done|4|4|4|4|4|4|4|4|1|1|1|1|4|2|100|2|4|3|2|4|3|3|2|3|4|1|1|4|2.5|20|4|4|4|4|4|4|4|4|0|4|4|5|4|4.25|1|4|5|2|3|41.67|4|4|4|4|4|4|3|3.86|3|4|4|4|2|4|3|3.43|12.54|4|4|4|4|2|2|3|2.33|71.67|3|3|3|2|4|3|0|2|2|2|2|0|4|4||||Green|||80.2||1|1|1|1|M|Black||17|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||52|28270|Bachelors Degree|Married|Business: Mgt, Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|0|1|502062408|1|0|1|500459576|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|472168|154145|4|3|45
502761850|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-18|2013-07-22|Baseline|2012-07-12|2012-07-18|Complete|Done|4|2|2|1|3|3|2.5|||||||||3|3|4|1|4|4|3.17|||||||||4|3|4|3.67||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Yellow||Volunteer: Moved|12.1||2|2|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||26|28212|Some College|Single|Military||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500012459|502762654|31|0|2|502925181|31|0|2|500623917|2||-2||4|2||500016374|-2||-2|0|10|||7496|10|||1|472351|-1|4|3|44
502728289|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-04|2017-03-09|Followup|2012-11-04|2013-01-09|Complete|Late|3|3|3|2|3|3|2.83|||||||||3|3|3|2|4|3|3|||||||||4|2|2|2.67||||||2|3|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child/Family: Moved|64.1||1|1|1|1|F|Hispanic||13|No|Mother|28278|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community||Match Support|F|White||32|28211||Married|Finance||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|502729186|3|0|2|502339145|1|0|2|500565493|2||-2||4|1|||-2|500000294|-2|0|3|||7496|10|||1|472960||4|3|45
502721278|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-12|NaT|Followup|2012-10-12|2012-10-02|Complete|Done|4|4|4|1|2|3|3|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Amachi, Cabarrus County||65.1||1|1|1|1|M|White||13|Yes|Mother|28025|One Parent: Female|Unknown||Yes||School|General Community|Cabarrus County|Match Support|M|White||47|28025||Single|Tech: Support, Writing|28026|0|2|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501938680|1|0|1|502701096|1|0|1|500560499|2||500003586||2|1|500000294, 500016374|500016374|-2|500016374|-2|0|4|||7464|9|||1|473193||4|3|45
501611456|BBBS of Greater Charlotte|Main Office|C|Active|2010-05-28|NaT|Followup|2013-05-28|2013-06-11|Complete|Done|4|2|4|1|3|4|3|||||||||1|3|3|3|1|3|2.33|||||||||4|4|4|4||||||3|3|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|3|3|3.33||||||2|4|3|||||2|2||||4|4||||Green|||81.6||1|1|1|1|M|Black||15|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black|Other African|32|28262||Married|Law: Police Officer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501611776|31|0|1|501876475|31|31|1|500450969|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|473310||4|3|45
500910040|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2014-05-08|Followup|2013-05-29|2013-07-25|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|59.3||1|1|1|1|M|White||21|No|Mother|28270|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||31|28209|||Human Services: Non-Profit|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|500910310|1|0|1|501600417|1|0|1|500363806|2||||4|3|||-2||-2|0|10|||7464|9|||1|473313||4|1|45
500771746|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2016-06-15|Followup|2013-05-29|2013-08-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Child: Graduated|84.6||3|4|1|2|F|Black||19||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||37|28012|Some College|Married|Finance: Banking|28208|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500772014|31|0|2|500996153|1|0|2|500366437|2||500004641||4|1|500004640||-2||-2|0|4|||7464|9|||1|473314||4|0|45
500186682|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2015-07-22|Followup|2013-07-20|2013-07-21|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|96.1||3|4|1|1|M|Black||20|Yes|Mother|28227|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|M|Black||57|28262||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|500887363|31|0|1|500184396|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|473343||4|3|45
502700500|BBBS of Greater Charlotte|Main Office|C|Active|2012-01-13|NaT|Followup|2013-01-13|2013-01-07|Complete|Done|4|2|1|3|2|1|2.17|||||||||1|3|3|3|2|4|2.67|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||4|1|2.5|||||2|2||||4|4||||Green|||62.1||1|1|1|1|M|Black||13|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|White||30|28202|Bachelors Degree|Single|Business: Sales|28212|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502701345|31|0|1|502824634|1|0|1|500589524|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|473532||4|3|45
502566369|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-17|NaT|Followup|2013-07-17|2013-07-10|Complete|Done|3|4|4|4|4|4|3.83|3|1|4|2|4|4|3|27.67|4|4|4|4|4|4|4|4|4|4|1|3|4|3.33|20.12|4|3|4|3.67|4|4|4|4|-8.25|5|5|5|5|5|3|5|4|5|4.25|17.65|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Green|||56||2|2|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||49|28215|Bachelors Degree|Married|Business: Mgt, Admin|28277|13|0|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|502566823|31|0|2|503065299|1|0|2|500622859|2||-2||2|1|||-2||-2|0|10|||7439|1|||1|473646|275023|4|3|45
502980958|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-17|NaT|Followup|2013-07-17|2013-07-12|Complete|Done|4|3|4|2|4|4|3.5|3|2|3|3|3|3|2.83|23.67|3|3|3|2|3|3|2.83|3|3|3|3|3|3|3|-5.67|3|4|4|3.67|4|3|4|3.67|0|3|4|3|4|3.5|4|4|3|3|3.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|1|1.5|3|3|3|-50|2|2|2|2|0|4|4|4|4|0|Green|||56||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Sales|28273|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502982410|31|0|1|503008664|1|0|1|500620394|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|473650|463519|4|3|45
502551048|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-19|2015-01-15|Followup|2012-10-19|2012-12-19|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Moved|38.9||1|1|2|2|F|Hispanic||13|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Enrollment|F|Black||52|30080|Bachelors Degree|Single|Consultant|2451|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502551498|3|0|2|501472128|31|0|2|500554178|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|473933||4|1|45
502591898|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-18|NaT|Followup|2013-07-18|2013-08-28|Complete|Done|4|1|4|2|3|2|2.67|3|3|4|2|3|4|3.17|-15.77|4|3|3|4|3|3|3.33|4|3|4|2|4|4|3.5|-4.86|4|4|3|3.67|4|4|4|4|-8.25|5|4|5|5|4.75|5|5|4|5|4.75|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|||55.9||2|2|1|1|F|Black||16|No|Mother|28214|Two Parent|$40,000 to $44,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28210|Masters Degree|Single|Medical: Healthcare Worker||1|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|502592415|31|0|2|503002003|31|0|2|500620503|2||-2||2|1||500004640, 500005291|-2||-2|0|4|||7496|10|||1|473958|294647|4|3|45
502907527|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-23|2014-11-21|Baseline|2012-07-18|2012-08-23|Complete|Done|4|1|4|1|4|4|3|||||||||4|4|4|4|1|4|3.5|||||||||4|4|4|4||||||3|5|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Moved|26.9||1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community|Amachi|Match Support|M|White||55|28202|Associate Degree|Married|Business||30|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502908938|31|0|1|502996593|1|0|1|500624606|2||-2||4|2||500000294|-2||-2|0|10|||7464|9|||1|473967|-1|4|3|44
502743091|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-18|2014-09-04|Followup|2013-07-18|2013-08-28|Complete|Done|4|4|4|3|3|3|3.5|4|4|4|4|4|4|4|-12.5|4|3|3|4|4|3|3.5|2|4|4|3|2|3|3|16.67|4|4|4|4|4|4|4|4|0|4|3|3|3|3.25|2|3|3|3|2.75|18.18|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3|3|3|33.33|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Lost contact with child/agency|25.6||1|1|1|1|M|Black||19|No|Mother|28215|One Parent: Female|$30,000 to $34,999|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||39|28203|Bachelors Degree|Single|Unemployed||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502743998|31|0|1|503079983|1|0|1|500623169|2||-2||4|2||500005291|-2||-2|6854|8|||7496|10|||1|473970|470985|4|3|45
503044619|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-03|2016-09-15|Baseline|2012-07-18|2012-08-03|Complete|Done|3|1|4|1|2|2|2.17|||||||||4|4|4|4|4|4|4|||||||||3|2|4|3||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2||||4|4||||Green||Child/Family: Moved|49.4||1|1|1|1|M|Black||15|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance: Banking|28202|0|7|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020910|503046265|31|0|1|503021454|1|0|1|500624634|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|474027|-1|4|3|44
502763968|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2016-09-08|Followup|2013-04-30|2013-06-12|Complete|Done|4|1|1|1|4|4|2.5|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red||Volunteer: Moved|52.3||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Enrollment|M|White||38|28206|Bachelors Degree|Divorced|Business: Mgt, Admin|28164|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502764880|31|0|1|502939016|1|0|1|500608284|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|474426||4|3|45
502912138|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-27|2013-06-28|Followup|2013-04-27|2013-04-22|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red||Volunteer: Moved|14||3|3|2|2|M|Black||13|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||33|28078|Bachelors Degree|Single|Business: Marketing|28036|5|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502913549|31|0|1|502881673|1|0|1|500610045|2||-2||4|3|||-2||-2|34|2|||7464|9|||1|474432||4|3|45
502839019|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-24|2016-01-28|Baseline|2012-07-19|2013-01-24|Complete|Done|4|3|4|4|4|4|3.83|||||||||3|4|3|2|4|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|3|2|3||||||3|3|3|||||1|1||||4|4||||Green||Volunteer: Moved|36.1||1|1|1|1|M|Black||17|No|Mother|28210|One Parent: Female|$40,000 to $44,999|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||32|28203|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502840311|31|0|1|502432390|31|0|1|500674451|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|474477|-1|4|3|44
501645192|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-21|2016-08-19|Followup|2013-07-21|2013-07-29|Complete|Done|3|3|4|3|2|3|3|||||||||4|4|4|2|3|3|3.33|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|85||1|1|2|2|M|Hispanic||19|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501645515|3|0|1|501519306|1|0|1|500374818|2||-2||4|3||500016374|-2|500016374|-2|0|10|||7464|9|||1|475331||4|3|45
500186956|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-21|2015-03-04|Followup|2013-06-21|2013-08-05|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|128.4||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28203|Bachelors Degree|Married|Law: Lawyer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|500189727|1|0|1|500037841|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|475336||4|1|45
500185647|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-09|2013-10-31|Followup|2013-07-09|2013-08-14|Complete|Done|3|3|3|3|4|4|3.33|||||||||3|4|4|4|3|4|3.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|123.8||1|2|1|2|F|Black||21|Yes|Mother|28217|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||38|28269|Bachelors Degree|Married|Unknown|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187284|31|0|2|500188649|31|0|2|500038124|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|475338||4|3|45
501716763|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-07|2016-11-11|Followup|2013-05-07|2013-07-22|Expired|Late||||||||1|1|1|1|1|1|1|||||||||2|1|2|2|3|2|2||||||3|3|3|3|||||||2|3|2|2|2.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||1|1|||||||Red||Child/Family: Lost contact with volunteer/agency|78.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Amachi, Cabarrus County|Match Support|F|Black||39|28269||Single|Self-Employed, Entrepreneur|28027|7|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501716992|31|0|2|502112513|31|0|2|500449029|2||-2||4|3||500000294, 500016374|-2|500016374|-2|6854|8|||7458|9|||1|475372|30228|4|0|45
502477677|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-29|2013-08-22|Followup|2013-07-29|2013-08-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|24.8||1|1|1|1|M|Black||13|No|Mother|28273|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||31|28217|Bachelors Degree|Single|Business: Engineer|28273|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|502478124|31|0|1|502621765|31|0|1|500545314|2||-2||4|3|||-2||-2|0|5|||7496|10|||1|475446||4|1|45
500896588|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2016-06-15|Followup|2013-07-20|2013-07-22|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|3|3|3|4|3|3|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|3|3|3.71||||||||||2|3|2|2.33||||||4|3|3.5|||||2|2||||4|4||||Green||Child: Graduated|106.9||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28273|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||36|28269|Masters Degree|Married|Education|28205|6|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|500896858|3|15|2|500924445|1|0|2|500183434|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|475449||4|3|45
501402710|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-19|2015-06-17|Followup|2013-06-19|2013-07-25|Complete|Done|2|2|3|3|3|3|2.67|||||||||2|3|3|3|2|3|2.67|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Moved|71.9||1|1|1|1|M|Black||18|No|Mother|30058|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28215||Married|Consultant|28285|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501402995|31|0|1|501728845|1|0|1|500368860|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|475451||4|3|45
502637589|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-19|2014-06-09|Followup|2013-07-19|2013-07-12|Complete|Done|2|4|2|1|4|4|2.83|4|2|2|1|2|4|2.5|13.2|1|4|3|2|3|4|2.83|1|4|3|3|1|1|2.17|30.41|3|4|3|3.33|4|4|4|4|-16.75|4|5|4|5|4.5|2|3|2|5|3|50|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|3|3.5|3|3|3|16.67|2|2|2|2|0|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Moved|34.7||1|1|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||30|28203|Masters Degree|Single|Business: Marketing|28203|0|10|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|502638284|31|0|2|502619035|1|0|2|500545174|2||-2||4|1|500005291|500005291|-2||-2|6854|8|||131|1|||1|475452|317220|4|3|45
500835156|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2016-11-10|Followup|2013-07-10|2013-09-03|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|100||1|2|1|2|M|Black||17||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Multi-Race (None of the above)||38|29710|Bachelors Degree|Single|Architect||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500835425|31|0|1|500466903|7|0|1|500277232|2||-2||4|1|||-2||-2|0|4|||46|2|||1|475455||4|1|45
502578459|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-23|NaT|Followup|2013-07-23|2013-07-25|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|Cabarrus County||55.8||1|1|1|1|M|Black||18|No|Mother|28025|One Parent: Female|$35,000 to $39,999||Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||48|28269|Some College|Married|Tech: Management|28204|10|0|AA Task Force|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502578962|31|0|1|502869485|31|0|1|500615803|2||500016307||2|2|500016374|500016374|-2|500016374|-2|6854|8|||9229|13|||1|475576|442607|4|3|45
501755470|BBBS of Greater Charlotte|Main Office|C|Active|2010-06-30|NaT|Followup|2013-06-30|2013-07-10|Complete|Done|4|3|4|3|4|4|3.67|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||2|2|1|1.67||||||4|3|3.5|||||2|2||||4|4||||Green|||80.5||2|2|2|2|F|Black||13|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|501755813|31|0|2|502038804|31|0|2|500456645|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|475959||4|3|45
500934908|BBBS of Greater Charlotte|Main Office|C|Active|2010-06-18|NaT|Followup|2013-06-18|2013-06-18|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||2|5|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi||80.9||2|2|1|1|M|Black||16|Yes|Aunt|28216|One Parent: Female|Less than $10,000|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||34|20175|Bachelors Degree|Single|Business: Sales|28211|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|500935173|31|0|1|502107314|1|0|1|500456443|2||500003586||2|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|475963||4|3|45
503005868|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-24|2017-02-26|Followup|2013-07-24|2013-07-24|Complete|Done|2|1|2|1|2|3|1.83|2|2|2|1|2|3|2|-8.5|1|2|3|1|1|3|1.83|2|2|3|2|2|3|2.33|-21.46|4|4|4|4|4|4|4|4|0|3|5|2|3|3.25|2|3|3|2|2.5|30|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|2|2.5|4|4|4|-37.5|2|2|2|2|0|4|4|4|4|0|Red||Child: Lost interest|55.1||1|1|1|1|M|Multi-race (Black & Hispanic)||15||Mother|28270|One Parent: Female|$25,000 to $29,999|Y|No||Therapist/Counselor|General Community||Match Support|M|White||51|28173|Bachelors Degree|Married|Consultant|28173|1|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020753|503007379|38|0|1|502935610|1|0|1|500623124|2||-2||4|3|||-2||-2|0|5|||7671|13|||1|476159|456253|4|3|45
503070961|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-21|2014-09-24|Baseline|2012-07-25|2012-08-21|Complete|Done|3|1|4|4|2|3|2.83|||||||||2|2|4|4|2|4|3|||||||||4|4|4|4||||||5|3|1|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|25.1||1|1|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|Amachi|Match Support|F|White||29|28209|||Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503072625|31|0|2|503034904|1|0|2|500628328|2||-2||4|3|500000294|500000294|-2||-2|0|4|||7464|9|||1|476341|-1|4|3|44
502183217|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-05|NaT|Followup|2013-08-05|2013-08-05|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|2|3||||||4|4|4|||||2|2||||4|4||||Green|Amachi||79.3||1|1|2|2|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|Black||50|28078|||Service: Restaurant|28082|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502183646|31|0|1|501733851|31|0|1|500462588|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|476381||4|3|45
502581001|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2014-01-30|Followup|2013-07-28|2013-08-21|Complete|Done|3|1|1|1|3|4|2.17|4|1|4|1|1|1|2|8.5|2|4|3|3|2|4|3|4|1|4|4|2|4|3.17|-5.36|4|4|4|4|4|4|3|3.67|8.99|4|2|3|5|3.5|5|4|4|5|4.5|-22.22|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|3|3.71|4.04|4|4|4|4|1|4|4|3|33.33|3|3|3|1|1|1|200|2|2|1|1|100|4|4||||Red||Volunteer: Feels incompatible with child/family|30.1||1|1|1|1|M|Black||15|No|Mother|28210|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013781|502581504|31|0|1|502650916|31|0|1|500547358|2||-2||4|3||500005291|-2|500000294|-2|34|2|||7496|10|||1|476512|321312|4|3|45
501618024|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-26|2016-01-08|Followup|2013-07-26|2013-07-24|Complete|Done|3|4|4|1|4|4|3.33|||||||||2|1|2|2|1|3|1.83|||||||||4|2|2|2.67||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|41.4||1|2|1|2|M|Hispanic||16||Mother|28031|Other/Unknown|Unknown||No||School|General Community||Match Support|M|White||65|28031|Some College|Married|Tech: Sales, Mktg|4241|5|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017777|501618344|3|0|1|501500078|1|0|1|500626248|2||-2||4|3|||-2||-2|0|4|||7462|13|||1|476703||4|3|45
502588461|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-22|2016-04-29|Followup|2013-07-22|2013-07-24|Complete|Done|4|3|3|2|4|4|3.33|3|3|2|2|2|3|2.5|33.2|3|4|3|4|3|3|3.33|3|4|4|3|2|4|3.33|0|4|3|4|3.67|4|3|4|3.67|0|4|4|4|4|4|4|5|4|5|4.5|-11.11|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|3|3|2|2.67|3|4|3|3.33|-19.82|2|3|2.5|4|4|4|-37.5|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Child: Graduated|57.3||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||46|28278|Bachelors Degree|Separated|Transport: Pilot|28208|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|502588977|31|0|1|502636478|31|0|1|500546741|2||-2||4|3|500005291|500005291|-2||-2|6854|8|||46|2|||1|476720|319772|4|3|45
501609876|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-13|2016-04-29|Followup|2013-07-13|2013-07-19|Comprehension|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Child: Graduated|81.5||1|2|1|2|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Black||38|28269|Masters Degree|Single|Medical: Nurse|28262|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501610196|31|0|2|501425392|31|0|2|500373716|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7464|9|||1|476780||4|2|45
503052850|BBBS of Greater Charlotte|Main Office|C|Active|2012-09-30|NaT|Baseline|2012-07-26|2012-09-29|Complete|Done|4|1|2|1|2|3|2.17|||||||||2|2|2|2|1|3|2|||||||||2|3|1|2||||||3|4|2|3|3|||||||4|4|4|4|4|3|4|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||53.5||1|1|1|1|F|Hispanic||13|No|Mother|28277|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||31|28210|Bachelors Degree|Single|Education: Teacher|29710|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020753|503027860|3|0|2|503028888|1|0|2|500626321|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|476823|-1|4|3|44
502980163|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-10|2013-08-30|Baseline|2012-07-26|2012-08-10|Complete|Done|3|2|2|1|2|2|2|||||||||1|1|3|2|2|3|2|||||||||3|3|3|3||||||2|3|5|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||2|3|1|2||||||2|2|2|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|12.6||1|1|1|1|M|Black||15|No|Mother|28105|One Parent: Female|$25,000 to $29,999|Y|No||Self|General Community||Match Support|M|Black||39|28110|Some College|Married|Business||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|502981615|31|0|1|502949611|31|0|1|500626324|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|476824|-1|4|3|44
501731841|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-05|2013-08-30|Followup|2013-06-05|2013-06-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|50.8||1|1|1|1|F|Black||18|Yes|Father|28210|One Parent: Male|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||49|28277|Bachelors Degree|Single|Business: Mgt, Admin||4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500008321|501732181|31|0|2|501182066|31|0|2|500367022|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||46|2|||1|477444||4|1|45
500478936|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-14|2013-11-11|Followup|2013-07-14|2013-08-28|Complete|Done|4|4|4|4|4|3|3.83|||||||||4|3|1|4|4|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|63.9||1|1|3|3|M|Black||21|No|Mother|28078|One Parent: Female|$25,000 to $29,999||No||Neighbor/Friend|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|500479187|31|0|1|501284751|31|0|1|500275964|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|8|||132|8|||1|477565||4|3|45
502252828|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2015-10-13|Followup|2013-08-03|2013-09-02|Declined|Done||||||||4|1|4|4|1|2|2.67|||||||||1|2|1|2|2|2|1.67||||||1|1|1|1|||||||4|3|2|1|2.5||||||||||4|4|4|4|4|4|4|4||||||2|2|3|2.33|||||4|3|3.5||||1|1||||4|4||Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|50.3||1|1|1|1|M|Black||15||GrandMother|28227|Grandparents|Unknown||No||Self|General Community|PERL 2014-2016|RTBM|M|White||27|28205|Associate Degree|Single|Law: Police Officer||0|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502253254|31|0|1|502602451|1|0|1|500547383|2||-2||4|1|500005291|500014681|-2|500005291|-2|0|10|||7496|10|||1|477589|320066|4|1|45
502802219|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-30|2014-02-27|Followup|2013-07-30|2013-08-28|Complete|Done|3|1|2|2|3|3|2.33|3|1|1|1|2|2|1.67|39.52|4|4|4|4|4|4|4|3|4|4|3|2|4|3.33|20.12|4|4|4|4|3|3|2|2.67|49.81|5|4|4|4|4.25|4|4|4|4|4|6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|4|4|3|3|3|3|33.33|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Time constraint|19||1|1|1|1|M|White||17|No|Mother|28209|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|M|White||35|28212|Some College|Single|Tech: Computer/Programmer|28212|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502803493|1|0|1|503060158|1|0|1|500623104|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|477748|470627|4|3|45
501994951|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2014-09-18|Followup|2013-06-15|2013-08-30|Expired|Late||||||||3|3|3|1|4|4|3|||||||||4|4|3|4|4|4|3.83||||||4|4|4|4|||||||4|5|5|4|4.5||||||||||4|4|4|3|3|3|3|3.43||||||3|3|3|3|||||3|1|2||||1|1|||||||Yellow||Volunteer: Lost contact with child/agency|51.1||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|Unknown||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||36|28078||Single|Customer Service||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501843047|31|0|2|502048623|31|0|2|500455478|2||-2||4|2|||-2||-2|7294|13|||7464|9|||1|477768|139614|4|0|45
500545328|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-02|2016-09-30|Followup|2013-07-02|2013-07-02|Complete|Done|3|4|4|2|3|2|3|||||||||3|4|4|2|2|3|3|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|3|2.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|99||3|3|1|1|F|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|F|Black||43|28208|Masters Degree|Single|Business: Sales|28078|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|2|501033808|31|0|2|500274449|2||-2||4|1|||-2||-2|0|10|||46|2|||1|477895||4|3|45
501240369|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-10-09|Followup|2013-07-10|2013-07-10|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|3|2|4|3|3.33|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|75||1|1|1|1|M|Black||20|Yes|Mother|28214|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||43|28269|Masters Degree|Single|Business: Mgt, Admin|28202|3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501240645|31|0|1|501240602|1|0|1|500272039|2||500003586||4|1|500000294|500000294|-2||-2|0|3|||131|1|||1|478020||4|3|45
502863776|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-31|NaT|Followup|2013-07-31|2013-09-13|Declined|Done||||||||2|2|3|4|3|4|3|||||||||2|3|3|3|3|3|2.83||||||4|4|4|4|||||||3|5|3|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||1|1|1||||1|1||||4|4||Green|||55.5||1|1|1|1|F|Black||14|No|Mother|28031|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Mgt, Admin|28078|1|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502865175|31|0|2|503029273|1|0|2|500622877|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|478193|434619|4|1|45
502863781|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-31|2015-01-30|Followup|2013-07-31|2013-09-13|Declined|Done||||||||3|4|3|2|3|4|3.17|||||||||2|4|3|2|1|2|2.33||||||4|4|4|4|||||||2|3|3|2|2.5||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||4|4|4||||1|1||||4|4||Red||Volunteer: Time constraint|30||1|1|1|1|M|Black||18|No|Mother|28031|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|M|White||26|28031|High School Graduate|Single|Personal Trainer/Coach|28117|0|4|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502865175|31|0|1|503002010|1|0|1|500621061|2||-2||4|3|||-2||-2|0|10|||17161|11|||1|478390|465050|4|1|45
501712048|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-22|NaT|Followup|2013-02-22|2013-03-07|Complete|Done|3|1|2|1|2|3|2|||||||||1|3|4|3|2|4|2.83|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green|Amachi||72.7||1|1|1|1|M|Black||13|Yes|Mother|28134|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||29|28273|Some College|Single|Govt: Mgmt/Admin|28208|2|0|Relative|Relative|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|501712386|31|0|1|502405439|1|0|1|500516322|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||17161|11|||1|478774||4|3|45
502859440|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-01|2014-04-21|Followup|2013-08-01|2013-08-28|Complete|Done|1|4|4|1|1|4|2.5|3|2|3|1|3|3|2.5|0|4|4|4|1|4|4|3.5|2|4|4|4|4|4|3.67|-4.63|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|4|4|5|4.5|11.11|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|4|3.5|14.29|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Time constraint|20.6||1|1|1|1|F|Hispanic|Mexican|15|No|Mother|28215|Two Parent|Unknown||Yes||School|General Community||Match Support|F|Multi-race (Hispanic & White)||30|28202|Bachelors Degree|Married|Finance: Banking|28255|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502860839|3|10|2|503046471|35|0|2|500623399|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|481257|401855|4|3|45
501938014|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-15|2013-04-10|Followup|2013-01-15|2013-04-01|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Feels incompatible with child/family|38.8||1|1|1|1|M|White||13|No|Mother|28083|One Parent: Female|Unknown|Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|RTBM|M|Hispanic||44|28081|Bachelors Degree|Single|Business: Mgt, Admin|28025|2|10|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|501938412|1|0|1|501874077|3|0|1|500426161|2||-2||4|1||500014681, 500016374|-2||-2|0|4|||7464|9|||1|481452||4|0|45
500186352|BBBS of Greater Charlotte|Main Office|C|Completed|2002-07-29|2014-01-02|Followup|2013-07-29|2013-08-29|Complete|Done|4|3|4|4|4|4|3.83|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|137.2||4|4|2|2|M|Black||21||Mother|28212|One Parent: Female|Unknown|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|White||45|28226|Masters Degree|Married|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500187945|31|0|1|500189280|1|0|1|500037290|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|481790||4|3|45
503044619|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-03|2016-09-15|Followup|2013-08-03|2013-09-02|Declined|Done||||||||3|1|4|1|2|2|2.17|||||||||4|4|4|4|4|4|4||||||3|2|4|3|||||||4|5|3|5|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||1|4|2.5||||2|2||||4|4||Green||Child/Family: Moved|49.4||1|1|1|1|M|Black||15|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance: Banking|28202|0|7|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020910|503046265|31|0|1|503021454|1|0|1|500624634|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|481833|474027|4|1|45
502353937|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-22|NaT|Followup|2012-11-22|2012-11-13|Complete|Done|4|4|4|1|4|4|3.5|||||||||3|4|4|1|3|4|3.17|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||75.8||1|1|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||31|29605|Bachelors Degree|Single|Business: Human Resources|29615|1|0|Local TV|Media|Big|General Community|Project Big AND Amachi|Match Support|277|60|598|500000170|500018851|502354375|31|0|2|501672025|1|0|2|500487322|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500004901|-2|0|4|||7438|1|||1|482089||4|3|45
502222545|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-03|2017-01-24|Followup|2013-08-03|2013-08-05|Complete|Done|1|3|1|4|1|2|2|||||||||1|1|3|1|2|3|1.83|||||||||4|4|4|4||||||2|2|5|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|77.7||1|1|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|F|White||37|28208|Masters Degree|Single|Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502222979|31|0|2|502196116|1|0|2|500462566|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|482120||4|3|45
502605331|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-13|NaT|Baseline|2012-08-06|2012-08-13|Complete|Done|3|4|4|1|3|3|3|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||1|1||||4|4||||Red|Cabarrus County||55.1||1|1|1|1|M|Hispanic||13|No|Mother|28027|One Parent: Female|$25,000 to $29,999||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||33|28036|Bachelors Degree|Married|Business||2|5|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502605848|3|0|1|503090281|1|0|1|500627504|2||500016307||2|3|500016374|500016374|-2|500016374|-2|34|2|||7464|9|||1|482204|-1|4|3|44
502839800|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-25|2014-08-12|Baseline|2012-08-06|2012-08-25|Complete|Done|4|3|3|3|3|3|3.17|||||||||2|4|4|3|3|4|3.33|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|23.6||1|1|1|1|M|Black||17|No|Mother|28213|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||29|28213|Bachelors Degree||Tech: Sales, Mktg|28213|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|503677894|31|0|1|502847446|1|0|1|500627524|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|482230|-1|4|3|44
501300101|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-14|2015-05-11|Followup|2013-08-14|2013-09-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|80.9||1|1|4|4|F|Black||19|Yes|GrandMother|28273|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501300379|31|0|2|500346193|31|0|2|500281421|2||500003586||4|2|500000294|500000294|-2||-2|7294|13|||46|2|||1|482413||4|1|45
501195410|BBBS of Greater Charlotte|Main Office|C|Active|2008-08-15|NaT|Followup|2013-08-15|2013-08-15|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|||103||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Asian||35|28210|Bachelors Degree|Married|Business: Sales|28217|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501195684|31|0|1|501277677|4|0|1|500278978|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|482414||4|3|45
502605248|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-07|2014-02-27|Followup|2013-08-07|2013-09-02|Declined|Done||||||||2|2|3|2|2|3|2.33|||||||||2|4|1|4|2|3|2.67||||||4|4|4|4|||||||4|2|5|4|3.75||||||||||4|4|4|4|4|4|4|4||||||3|3|2|2.67|||||4|4|4||||2|2||||4|4||Green||Volunteer: Time constraint|18.7||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|Unknown||Yes||Relative|General Community|Project Big|Enrollment|M|White||36|28205|Masters Degree|Single|Finance: Banking||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502137975|31|0|1|503049689|1|0|1|500623109|2||-2||4|1||500004640|-2||-2|0|3|||7496|10|||1|482516|470640|4|1|45
502142541|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-18|2015-07-23|Followup|2013-06-18|2013-07-31|Complete|Done|4|3|3|3|3|3|3.17|3|4|4|3|4|4|3.67|-13.62|4|4|4|3|3|4|3.67|3|3|3|3|3|3|3|22.33|4|4|4|4|4|4|4|4|0|5|5|5|5|5|4|4|5|3|4|25|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|3|4|4|3.67|4|4|4|4|-8.25|3|3|3|2|2|2|50|2|2|2|2|0|4|4||||Green||Child: Graduated|61.1||1|1|2|2|F|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502142970|31|0|2|501905673|31|0|2|500455759|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|482571|141478|4|3|45
501721760|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-22|2016-11-01|Followup|2013-06-22|2013-09-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Infraction of match rules/agency policies|88.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||59|28269|Masters Degree|Married|Clergy||0|0|Coca Cola|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|501722098|31|0|1|501755476|1|0|1|500368545|2||-2||4|1|||-2|500000294|-2|0|10|||9610|3|||1|482572||4|0|45
500910037|BBBS of Greater Charlotte|Main Office|C|Active|2009-06-22|NaT|Followup|2013-06-22|2013-09-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||92.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||46|28277||Married|Business: Mgt, Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|500910307|31|0|1|500856100|1|0|1|500368834|2||-2||2|1|||-2||-2|0|10|||46|2|||1|482573||4|0|45
501288021|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-27|2016-02-01|Followup|2013-08-27|2013-08-30|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|1|1.5|||||2|2||||4|4||||Green||Volunteer: Moved|89.2||1|1|1|1|F|Black||16|No|Mother|28211|Two Parent|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28027|PHD|Single|Education: College Professor|27411|1|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501288299|31|0|2|501249338|31|0|2|500281778|2||-2||4|1|||-2||-2|0|10|||46|2|||1|482701||4|3|45
501641325|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-24|2015-08-03|Followup|2013-06-24|2013-09-08|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|73.3||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Multi-race (Asian & White)||34|28205|Bachelors Degree|Single|Tech: Research/Design|28255|3|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|1|501715652|37|0|1|500366872|2||-2||4|1||500000294|-2|500000294|-2|6854|8|||7464|9|||1|482770||4|0|45
501488919|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-09|2015-08-25|Followup|2013-08-09|2013-08-08|Complete|Done|4|2|4|1|3|4|3|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|3|3|3.71||||||||||3|3|3|3||||||2|2|2|||||2|2||||4|4||||Yellow||Child: Lost interest|36.5||1|2|1|2|F|Black||17||Mother|28031|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||36|28205|Bachelors Degree|Single|Business: Mgt, Admin|28036|0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501489205|31|0|2|501392684|31|0|2|500626771|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|482974||4|3|45
501513669|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-09|2015-02-04|Followup|2013-08-09|2013-07-22|Complete|Early|3|3|2|3|1|2|2.33|||||||||3|3|3|2|3|3|2.83|||||||||4|4|4|4||||||3|3|4|4|3.5|||||||4|4|4|4|4|3|3|3.71||||||||||3|4|2|3||||||3|4|3.5|||||1|1||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|29.9||1|2|2|3|F|White||18|No|Mother|28031|Other/Unknown|Unknown||No||School|General Community||Match Support|F|White||68|28036||Divorced|Business: Sales||5|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011349|501513961|1|0|2|500824400|1|0|2|500626772|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|482975||4|3|45
502300563|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-09|NaT|Followup|2013-08-09|2013-08-20|Complete|Done|3|4|4|3|3|4|3.5|3|3|4|1|3|4|3|16.67|3|4|3|4|4|4|3.67|4|4|3|4|3|4|3.67|0|4|4|4|4|4|4|4|4|0|5|4|4|5|4.5|4|4|5|5|4.5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|2|3.71|4.04|4|4|4|4|4|4|3|3.67|8.99|4|2|3|2|3|2.5|20|2|2|1|1|100|4|4||||Green|||55.2||1|2|1|2|M|Black||15|No|Mother|28031|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Black||53|28078|PHD|Married|Medical|28078|2|0|AA Task Force|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020753|502300995|31|0|1|502101059|31|0|1|500626773|2||-2||2|1|||-2||-2|0|4|||11098|8|||1|482976|177594|4|3|45
501160242|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-09|2016-11-07|Followup|2013-08-09|2013-09-06|Complete|Done|3|2|2|3|1|2|2.17|||||||||2|2|2|2|2|3|2.17|||||||||3|3|3|3||||||3|2|4|3|3|||||||4|4|3|4|4|4|3|3.71||||||||||2|3|3|2.67||||||1|4|2.5|||||2|2||||4|4||||Red|Cabarrus County|Volunteer: Lost contact with child/agency|51||3|4|1|2|F|White||17|No|GrandFather|28147|Grandparents|Unknown||No||School|General Community|Cabarrus County|Match Support|F|White||29|28078||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501160516|1|0|2|502325100|1|0|2|500626774|2||500016307||4|3|500016374|500016374|-2|500016374|-2|0|4|||7496|10|||1|482977||4|3|45
501809541|BBBS of Greater Charlotte|Main Office|C|Active|2009-08-07|NaT|Followup|2013-08-07|2013-09-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||91.3||1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||49|28031|Bachelors Degree|Married|Transport: Pilot|40223|9|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501809896|36|0|1|501620528|1|0|1|500375025|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|482990||4|1|45
502529397|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-11|NaT|Followup|2013-08-11|2013-09-18|Complete|Done|2|1|4|1|4|4|2.67|||||||||1|3|3|2|2|4|2.5|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|Project Big||67.2||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||48|28216|Bachelors Degree|Married|Finance: Banking|28255|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502529850|31|0|1|500188946|31|0|1|500548763|2||500004641||2|1|500004640||-2||-2|6854|8|||7464|9|||1|483014||4|3|45
501092822|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-09|2014-04-23|Followup|2013-08-09|2013-09-22|Complete|Done|1|4|4|4|4|4|3.5|||||||||1|4|4|4|4|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Time constraint|20.4||3|4|2|3|F|Black||14|No|Mother|28217|Two Parent|$15,000 to $19,999|Y|No||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||34|28215|Bachelors Degree|Single|Tech: Computer/Programmer|28262|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501093096|31|0|2|500473347|31|0|2|500627441|2||-2||4|3||500014505, 500016394|-1||-2|0|4|||46|2|||1|483018||4|3|45
501631140|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-17|2016-03-03|Followup|2013-06-17|2013-07-22|Complete|Done|4|2|1|1|4|3|2.5|||||||||2|4|4|4|3|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|2|4|4|3.71||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Volunteer: Moved|80.5||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Service: Hotel|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501631463|31|0|1|501628976|1|0|1|500367187|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|483346||4|3|45
500185778|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-17|2016-06-23|Followup|2013-06-17|2013-06-19|Complete|Done|3|1|2|1|1|1|1.5|||||||||3|3|4|3|2|3|3|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||1|4|2.5|||||2|2||||4|4||||Green||Child: Graduated|144.2||1|1|1|1|M|Black||18||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||42|27514||Married|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187368|31|0|1|500188776|1|0|1|500036776|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|483347||4|3|45
500915359|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-10|2014-12-18|Followup|2013-08-10|2013-09-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|28.3||3|3|1|1|F|Black||19|No|Mother|28227|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28204|Bachelors Degree|Single|Medical: Nurse||0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500915629|31|0|2|503044413|1|0|2|500622861|2||-2||4|2|||-2||-2|34|2|||7496|10|||1|483354||4|1|45
502813454|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-13|NaT|Followup|2013-08-13|2013-08-12|Complete|Done|4|2|4|1|2|4|2.83|3|1|2|1|4|3|2.33|21.46|4|2|4|2|3|4|3.17|2|3|2|1|1|3|2|58.5|4|4|4|4|4|4|4|4|0|4|3|4|3|3.5|2|3|3|1|2.25|55.56|4|4|4|4|4|4|2|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|4|4|1|1|1|1|300|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|||55.1||1|2|1|2|F|White||14|No|Mother|28031|Two Parent|Unknown||Yes||School|General Community||Match Support|F|White||61|28031|Bachelors Degree|Divorced|Business: Mgt, Admin||5|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500020752|502814731|1|0|2|502855397|1|0|2|500627861|2||-2||2|1|||-2||-2|0|4|||129|1|||1|483723|390213|4|3|45
502605331|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-13|NaT|Followup|2013-08-13|2013-08-12|Complete|Done|3|4|4|2|4|4|3.5|3|4|4|1|3|3|3|16.67|2|3|3|2|3|3|2.67|2|4|3|4|4|3|3.33|-19.82|4|4|4|4|4|4|4|4|0|3|5|3|5|4|5|5|5|4|4.75|-15.79|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|3|4|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Red|Cabarrus County||55.1||1|1|1|1|M|Hispanic||13|No|Mother|28027|One Parent: Female|$25,000 to $29,999||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||33|28036|Bachelors Degree|Married|Business||2|5|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502605848|3|0|1|503090281|1|0|1|500627504|2||500016307||2|3|500016374|500016374|-2|500016374|-2|34|2|||7464|9|||1|483726|482204|4|3|45
502478700|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-09|2014-11-13|Followup|2013-08-09|2013-08-13|Complete|Done|4|3|4|4|3|4|3.67|4|4|4|2|2|4|3.33|10.21|2|2|4|1|4|4|2.83|2|4|4|3|4|4|3.5|-19.14|4|4|4|4|4|4|4|4|0|5|4|5|5|4.75|5|4|5|5|4.75|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|3|3|4|4|3|3.67|-18.26|3|3|3|2|2|2|50|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|39.2||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28027|Masters Degree|Single|Business: Engineer|28262|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|277|60|598|500000170|500013781|502881024|31|0|1|502578355|1|0|1|500544505|2||-2||4|3|500005291|500005291|-2|500015184|-1|0|5|||7462|13|||1|483769|315352|4|3|45
502869635|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-13|2014-08-21|Baseline|2012-08-13|2012-11-13|Complete|Done|4|4|4|4|3|4|3.83|||||||||3|3|4|3|3|3|3.17|||||||||4|4|4|4||||||4|4|5|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||4|3|3.5|||||2|2||||4|4||||Red||Volunteer: Moved|21.2||1|1|1|1|F|Black||17|No|Mother|28206|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community||Match Support|F|Black||34|28210|Bachelors Degree|Single|Business: Marketing||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502871029|31|0|2|503099564|31|0|2|500649374|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|483786|-1|4|3|44
501261979|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-22|2014-10-13|Followup|2013-07-22|2013-09-24|Complete|Late|3|4|4|2|4|3|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|74.7||1|1|3|3|F|Black||15|No|Mother|28134|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||55|28173||Married|Human Services: Non-Profit|28205|0|0|Coworker|Workplace Partner|Big|General Community|VOL - Maximizing Match Impact|Match Support|277|60|598|500000170|500011349|501262256|31|0|2|500418936|31|0|2|500278634|2||-2||4|1|||-2|500011314|-2|0|10|||7447|3|||1|483825||4|3|45
502249189|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-23|2016-09-22|Followup|2013-03-23|2013-04-29|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|66||1|1|1|1|M|Black||13|No|Mother|28277|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||34|28262||Married|Finance|29715|6|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Enrollment|277|60|598|500000170|500017732|502249620|31|0|1|502485458|31|0|1|500523907|2||-2||4|1|||-2||-2|34|2|||7462|13|||1|483965||4|1|45
501662021|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-14|2014-02-21|Followup|2013-08-14|2013-07-22|Complete|Early|3|1|4|1|2|3|2.33|3|1|4|1|1|3|2.17|7.37|2|4|4|3|2|3|3|2|4|4|4|4|3|3.5|-14.29|4|4|4|4|4|4|3|3.67|8.99|5|3|2|3|3.25|5|4|3|3|3.75|-13.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|2|4|1|2.33|3|4|3|3.33|-30.03|3|3|3|4|1|2.5|20|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|18.3||2|2|1|1|M|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|Black||50|28269|Some College|Divorced|Retired||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500011349|501090456|31|0|1|502902255|31|0|1|500627357|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|484022|468082|4|3|45
502236953|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-17|2015-01-30|Followup|2013-08-17|2013-10-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|53.5||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||50|28212|Some College|Married|Law: Police Officer||2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502237384|31|0|1|502232559|31|0|1|500464143|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|484159||4|1|45
501825910|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-24|2016-09-23|Followup|2013-08-24|2013-08-27|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|85||1|1|1|1|M|Black||16|Yes|Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|White||51|28214|Masters Degree|Married|Business: Sales|94108|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|501196986|1|0|1|500380446|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||7496|10|||1|484160||4|3|45
503023832|BBBS of Greater Charlotte|Main Office|C|Active|2013-05-31|NaT|Baseline|2012-08-14|2013-05-31|Complete|Done|4|2|2|2|2|2|2.33|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||45.5||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|White||33|28278|Bachelors Degree|Single|Arts, Entertainment, Sports|28269|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|503025372|31|0|1|503139766|1|0|1|500692957|2||-2||2|1|||-2||-2|0|10|||7671|13|||1|484219|-1|4|3|44
501721579|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-24|2016-06-17|Followup|2013-07-24|2013-09-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Moved|82.8||2|2|1|1|F|Multi-Race (None of the above)||14|No|Mother|28211|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||50|28227|Some College|Single|Human Services: Social Worker||2|5|St. Paul Baptist|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501721919|7|0|2|501687513|31|0|2|500375006|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||9609|7|||1|484529||4|1|45
502083465|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-06|2013-06-06|Followup|2012-10-06|2012-09-26|Complete|Done|3|1|1|1|3|3|2|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Moved|20||1|1|2|2|F|Black||13|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||69|28027||Married|Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500012459|502083880|31|0|2|502591360|31|0|2|500557052|2||-2||4|1|||-2|500016374|-2|0|10|||7464|9|||1|484562||4|3|45
501101149|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-01|NaT|Followup|2014-07-01|2014-08-15|Complete|Done|3|2|3|2|4|4|3|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||4|4|4|||||2|2||||4|4||||Yellow|||104.5||1|2|1|2|F|White||16||Mother|28270|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||55|28277|Masters Degree|Widowed|Consultant||5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|501101423|1|0|2|500834694|1|0|2|500276073|2||-2||2|2|||-2||-2|0|4|||7671|13|||1|484686||4|3|45
502785308|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-16|NaT|Followup|2013-08-16|2013-08-15|Complete|Done|4|4|4|1|4|4|3.5|3|2|2|2|1|3|2.17|61.29|4|4|4|4|1|3|3.33|2|4|3|1|2|4|2.67|24.72|4|4|4|4|2|2|2|2|100|2|4|5|5|4|2|5|2|5|3.5|14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Green|Cabarrus County||55||1|2|1|2|F|American Indian or Alaska Native||16|No|Aunt|28027|One Parent: Male|Unknown||Yes||School|General Community|Cabarrus County|Match Support|F|White||49|28027|Bachelors Degree|Married|Business: Marketing|28025|14|0|ACN|Workplace Partner|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|504347632|6|0|2|502736971|1|0|2|500628695|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|4|||13581|3|||1|484930|359572|4|3|45
502643010|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-30|2014-07-31|Baseline|2012-08-16|2013-03-30|Complete|Done|3|4|4|4|1|1|2.83|||||||||3|3|3|4|2|3|3|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Yellow||Volunteer: Lost contact with child/agency|16||1|1|1|1|M|Black||14|Yes|Mother|28262|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Enrollment|M|Black||30|28203|Bachelors Degree|Single|Finance|28255|3|5|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502643706|31|0|1|503262615|31|0|1|500686907|2||500003586||4|2||500000294|-2|500000294|-2|6854|8|||6247|12|||1|484989|-1|4|3|44
503043863|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-04|2014-02-27|Baseline|2012-08-16|2012-09-04|Complete|Done|3|3|4|4|4|4|3.67|||||||||1|3|3|2|2|3|2.33|||||||||4|4|3|3.67||||||3|5|3|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|2|3|||||1|1||||4|4||||Red||Volunteer: Feels incompatible with child/family|17.8||1|1|1|1|M|Hispanic||15|No|Mother|28211|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|Asian||32|28204|Bachelors Degree|Single|Medical: Admin|28203|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|503045507|3|0|1|502996721|4|0|1|500629081|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|484993|-1|4|3|44
503071479|BBBS of Greater Charlotte|Main Office|C|Active|2012-09-30|NaT|Baseline|2012-08-17|2012-09-30|Complete|Done|3|3|3|3|2|2|2.67|||||||||3|2|2|3|3|2|2.5|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3|||||||||||||2|2||||4|4||||Green|||53.5||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||28|28269|Some College|Single|Business: Clerical||0|3|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020910|503069483|31|0|1|503051382|1|0|1|500629193|2||-2||2|1|||-2||-2|0|10|||7671|13|||1|485271|-1|4|3|44
502619926|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-09|2015-05-05|Followup|2013-08-09|2013-08-14|Complete|Done|3|4|4|4|3|3|3.5|||||||||4|4|3|2|4|3|3.33|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Project Big|Volunteer: Lost contact with child/agency|44.8||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||38|28205|Bachelors Degree|Single|Law: Lawyer|28202|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502620542|31|0|2|502642260|1|0|2|500548116|2||500004641||4|1|500004640||-2||-2|0|10|||7464|9|||1|485286||4|3|45
502431187|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-17|2016-01-07|Followup|2013-08-17|2013-09-02|Declined|Done||||||||3|2|4|1|3|4|2.83|||||||||2|3|3|2|3|3|2.67||||||2|4|4|3.33|||||||4|3|5|3|3.75||||||||||4|4|4|4|4|4|3|3.86||||||3|2|3|2.67|||||2|3|2.5||||2|2||||4|4||Yellow||Volunteer: Time constraint|40.7||2|2|1|1|F|Black||17|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|RTBM|F|White||41|28105|Bachelors Degree|Divorced|Business|28112|1|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|502431630|31|0|2|503015009|1|0|2|500627361|2||-2||4|2||500005291|-2||-2|0|5|||46|2|||1|485331|272216|4|1|45
502631914|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2014-08-28|Followup|2013-07-28|2013-07-28|Complete|Done|4|4|4|4|4|4|4|4|4|4|1|4|4|3.5|14.29|2|3|4|3|1|4|2.83|1|1|3|3|1|4|2.17|30.41|4|4|4|4|4|4|4|4|0|4|5|5|5|4.75|4|5|5|4|4.5|5.56|4|4|4|4|3|4|4|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|3|2.5|1|3|2|25|2|2|1|1|100|4|4||||Red||Volunteer: Moved|37||1|1|1|1|F|Black||18|No|Mother|28215|One Parent: Female|$20,000 to $24,999||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||37|28205|Associate Degree|Single|Medical: Healthcare Worker|28205|7|10|Local Print|Media|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013781|502632569|31|0|2|502581901|1|0|2|500546271|2||-2||4|3||500005291|-2|500004640|-2|6854|8|||7439|1|||1|485397|318565|4|3|45
503070961|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-21|2014-09-24|Followup|2013-08-21|2013-11-05|Expired|Late||||||||3|1|4|4|2|3|2.83|||||||||2|2|4|4|2|4|3||||||4|4|4|4|||||||5|3|1|4|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Red|Amachi|Child/Family: Lost contact with volunteer/agency|25.1||1|1|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|Amachi|Match Support|F|White||29|28209|||Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503072625|31|0|2|503034904|1|0|2|500628328|2||-2||4|3|500000294|500000294|-2||-2|0|4|||7464|9|||1|486002|476341|4|0|45
502255223|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-11|NaT|Followup|2013-08-11|2013-08-28|Complete|Done|4|1|4|1|2|4|2.67|||||||||4|3|4|2|4|2|3.17|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||79.1||1|1|1|1|F|Hispanic||14|No|Mother|28212|One Parent: Female|Unknown|Y|No|Spanish Radio|Media|General Community||Match Support|F|White||33|28209||Single|Education: Teacher||0|0||High School Partner|Big|General Community||Match Support|277|60|598|500000170|500020753|502255655|3|0|2|501823103|1|0|2|500463922|2||-2||2|1|||-2||-2|7068|1|||0|4|||1|486331||4|3|45
501987736|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-29|2014-06-18|Followup|2013-06-29|2013-07-22|Complete|Done|3|2|2|3|1|2|2.17|4|4|4|2|4|4|3.67|-40.87|2|2|2|2|2|2|2|2|4|4|2|4|4|3.33|-39.94|4|4|3|3.67|4|2|2|2.67|37.45|2|3|4|4|3.25|4|3|3|3|3.25|0|4|3|4|3|4|4|4|3.71|4|4|4|4|4|4|4|4|-7.25|3|4|3|3.33|3|4|3|3.33|0|3|2|2.5|2|1|1.5|66.67|2|2|1|1|100|4|4||||Green||Child: Graduated|47.6||1|1|1|1|F|White||20|No|Father|28217|One Parent: Male|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||40|28203|Masters Degree|Single|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501988135|1|0|2|502109789|1|0|2|500456045|2||-2||4|1|||-2||-2|6855|8|||7464|9|||1|486806|142908|4|3|45
500881634|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-14|NaT|Followup|2013-07-14|2013-09-03|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||104||1|2|1|2|M|Black||18||Mother|28213|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||38|28213||Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500881903|31|0|1|500816190|31|0|2|500277615|2||-2||2|1|||-2||-2|0|4|||46|2|||1|486850||4|1|45
502097843|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-29|2016-08-11|Followup|2013-08-29|2013-10-14|Declined|Late||||||||3|2|2|1|4|3|2.5|||||||||2|3|3|2|3|3|2.67||||||4|4|4|4|||||||3|3|3|4|3.25||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||3||||||2|2||||4|4||Green|2010-2012 OJJDP JJI|Child: Lost interest|59.4||1|1|2|2|M|Black||17|No|Mother|28078|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500021785|502098263|31|0|1|502643791|3|0|1|500550390|2||-2||4|1|500005291||-2||-2|0|10|||7496|10|||1|486888|330290|4|1|45
502907527|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-23|2014-11-21|Followup|2013-08-23|2013-09-09|Complete|Done|4|4|4|1|4|4|3.5|4|1|4|1|4|4|3|16.67|4|4|4|1|4|4|3.5|4|4|4|4|1|4|3.5|0|4|4|4|4|4|4|4|4|0|4|5|4|3|4|3|5|3|3|3.5|14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Moved|26.9||1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community|Amachi|Match Support|M|White||55|28202|Associate Degree|Married|Business||30|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502908938|31|0|1|502996593|1|0|1|500624606|2||-2||4|2||500000294|-2||-2|0|10|||7464|9|||1|486927|473967|4|3|45
500280148|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-13|NaT|Followup|2013-07-13|2013-07-21|Complete|Done|3|3|4|4|4|4|3.67|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Yellow|Amachi||80.1||3|3|1|1|F|Black||16|Yes|Mother|28205|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|F|Black||30|28216|Bachelors Degree|Single|Human Services: Non-Profit|28216|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188151|31|0|2|502118494|31|0|2|500460767|2||500003586||2|2|500000294|500000294|-2||-2|0|3|||7464|9|||1|487274||4|3|45
502233625|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-24|2013-10-22|Followup|2013-08-24|2013-09-02|Declined|Done||||||||3|3|3|2|1|3|2.5|||||||||2|3|3|3|4|3|3||||||4|4|4|4|||||||3|5|4|4|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4||||2|2|||||||Red||Child/Family: Moved|13.9||3|3|1|1|F|Multi-race (Hispanic & White)||17|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||30|28209|Associate Degree|Single|Medical: Nurse|28210|2|6|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500011746|502234056|35|0|2|503081963|1|0|2|500628685|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|487374|168274|4|1|45
502272172|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-24|2014-09-04|Followup|2013-08-24|2013-09-02|Declined|Done||||||||3|4|4|1|4|4|3.33|||||||||2|4|2|1|3|3|2.5||||||4|4|4|4|||||||2|3|3|4|3||||||||||4|4|4|4|4|4|4|4||||||1|1|1|1|||||4|3|3.5||||1|1||||4|4||Yellow||Volunteer: Lost contact with child/agency|24.3||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||27|28036|Bachelors Degree|Single|Business|28078|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502272604|31|0|2|502965088|1|0|2|500626278|2||-2||4|2|||-2||-2|6854|8|||7464|9|||1|487378|243094|4|1|45
501641337|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-07|2015-03-13|Followup|2013-08-07|2013-10-03|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|67.2||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||31|28269|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|2|500835981|31|0|2|500373972|2||-2||4|1||500000294|-2|500000294|-2|0|10|||46|2|||1|487395||4|1|45
502839800|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-25|2014-08-12|Followup|2013-08-25|2013-09-02|Declined|Done||||||||4|3|3|3|3|3|3.17|||||||||2|4|4|3|3|4|3.33||||||4|4|4|4|||||||3|4|3|4|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Green||Volunteer: Moved|23.6||1|1|1|1|M|Black||17|No|Mother|28213|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||29|28213|Bachelors Degree||Tech: Sales, Mktg|28213|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|503677894|31|0|1|502847446|1|0|1|500627524|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|487525|482230|4|1|45
501726201|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2015-01-30|Followup|2013-07-08|2013-08-07|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Moved|66.8||1|1|1|1|F|Black||17|Yes|Mother|28212|One Parent: Female|Unknown||Yes|YeaGod|Faith Organization|General Community|Amachi|Match Support|F|Black||51|28262|PHD|Married|Real Estate: Realtor||0|0|Weeping Willow|Faith Organization|Big|General Community||Enrollment|277|60|598|500000170|500008321|501726541|31|0|2|501734664|31|0|2|500371036|2||-2||4|3|500000294|500000294|-2||-2|5634|9|||9218|7|||1|487887||4|1|45
502636177|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-29|2013-09-19|Followup|2013-08-29|2013-09-04|Complete|Done|4|1|3|1|4|4|2.83|4|1|4|1|4|3|2.83|0|4|4|4|4|3|4|3.83|4|4|4|4|3|4|3.83|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|4|4|4|4|4|25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|1|1|1|1|0|4|4|4|4|0|Green||Volunteer: Moved|24.7||1|1|1|1|F|Black||14|No|GrandMother|28216|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|Black||30|28212||Single|Medical||0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502636872|31|0|2|502643313|31|0|2|500551053|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|488268|330694|4|3|45
501749652|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-01|2013-11-07|Followup|2013-09-01|2013-10-29|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Moved|38.2||1|1|2|2|M|Black||18||Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|Black||52|28107|Some College|Divorced|Tech: Engineer|28262|3|0|Local Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500012459|501749994|31|0|1|501645507|31|0|1|500464305|2||-2||4|2|||-2||-2|0|10|||7437|1|||1|488859|38597|4|1|45
503158441|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-14|2014-07-03|Baseline|2012-08-29|2012-09-14|Complete|Done|4|3|4|1|4|4|3.33|||||||||2|3|4|2|1|4|2.67|||||||||4|4|4|4||||||5|3|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||4|2|3|||||2|2||||4|4||||Red||Volunteer: Moved|21.6||1|1|1|1|F|Black||19|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||27|28202|Bachelors Degree|Single|Business||1|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503160119|31|0|2|503130365|1|0|2|500631432|2||-2||4|3|||-2|500000294|-2|0|5|||7464|9|||1|488914|-1|4|3|44
500958307|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-19|NaT|Followup|2013-09-19|2013-09-16|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|2|2|3|2.83|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|Amachi, Cabarrus County||113.9|Y|1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$40,000 to $44,999|Y|No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|Black||62|28213||Married|Finance: Economist||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500958577|31|0|1|500876132|31|0|1|500193868|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|488936||4|3|45
503108699|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-14|2014-08-11|Baseline|2012-08-30|2012-09-14|Complete|Done|3|3|4|1|2|3|2.67|||||||||2|2|3|2|2|3|2.33|||||||||4|2|2|2.67||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|22.9||1|1|1|1|M|White||19|No|Mother|28031|One Parent: Female|$30,000 to $34,999|Y|No||Self|General Community||Match Support|M|White||37|28036|Bachelors Degree|Single|Business: Sales|28117|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503110361|1|0|1|503106216|1|0|1|500631547|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|489246|-1|4|3|44
503021417|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-11|2015-10-16|Baseline|2012-08-30|2012-09-11|Complete|Done|3|3|4|2|3|4|3.17|||||||||3|4|3|2|3|3|3|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Yellow||Child/Family: Moved|37.1||1|1|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|White||32|28204|Bachelors Degree|Single|Business: Marketing|29730|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|501428579|31|0|2|503115600|1|0|2|500631553|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|489252|-1|4|3|44
503017622|BBBS of Greater Charlotte|Main Office|C|Inactive|2012-09-19|NaT|Baseline|2012-08-31|2012-09-19|Complete|Done|3|2|2|2|2|||||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|||53.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|$30,000 to $34,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|F|White||33|28207|Bachelors Degree|Married|Business||0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|503019155|31|0|2|503095382|1|0|2|500631726|2||-2||3|1|||-2||-2|34|2|||7464|9|||1|489657|-1|4|3|44
500480596|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-13|2014-01-16|Followup|2013-09-13|2013-09-30|Complete|Done|4|3|4|4|4|4|3.83|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||5|5||5||||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|88.1||1|1|1|1|M|Black||21|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Married|Business: Sales|28203|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500480847|31|0|1|500491267|1|0|1|500120915|2||500003586||4|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|489671||4|3|45
503043863|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-04|2014-02-27|Followup|2013-09-04|2013-11-19|Expired|Late||||||||3|3|4|4|4|4|3.67|||||||||1|3|3|2|2|3|2.33||||||4|4|3|3.67|||||||3|5|3|5|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||4|2|3||||1|1||||4|4||Red||Volunteer: Feels incompatible with child/family|17.8||1|1|1|1|M|Hispanic||15|No|Mother|28211|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|Asian||32|28204|Bachelors Degree|Single|Medical: Admin|28203|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|503045507|3|0|1|502996721|4|0|1|500629081|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|490240|484993|4|0|45
501604443|BBBS of Greater Charlotte|Main Office|C|Active|2009-07-10|NaT|Followup|2013-07-10|2013-09-24|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||92.2||1|1|1|1|M|Black||18|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||35|28209|Bachelors Degree|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501729878|1|0|1|500371104|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|490282||4|0|45
502222992|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-16|2013-12-12|Followup|2013-07-16|2013-09-03|Declined|Late||||||||3|3|3|1|2|3|2.5|||||||||2|4|3|2|2|4|2.83||||||4|4|3|3.67|||||||3|4|4|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Child: Graduated|40.9||1|1|1|1|F|Black||21|No|Aunt|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||32|28213|Bachelors Degree|Single|Education|28223|7|0|BBBS National Site|Web Link|Big|General Site||Enrollment|277|60|598|500000170|500017732|502223423|31|0|2|502085103|31|0|2|500461244|2||-2||4|1|||-2||-1|6854|8|||46|2|||1|490284|157522|4|1|45
502034144|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-20|2014-12-04|Followup|2013-07-20|2013-07-12|Complete|Done|3|3|4|3|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|52.5||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||RTBM|M|Some Other Race||45|28210|Bachelors Degree|Married|Education: Teacher||0|0|CIS/Hidden Valley|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500018987|502034543|31|0|1|502212267|41|0|1|500460434|2||||4|1|||-2||-2|34|2|||11522|6|||1|490285||4|3|45
501831581|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-29|NaT|Followup|2013-09-29|2013-09-26|Complete|Done|3|4|1|2|4|3|2.83|||||||||2|4|3|2|1|3|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Amachi||89.5||1|1|2|3|F|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||38|28273||Single|Tech: Engineer||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501831944|31|0|2|500715453|31|0|2|500387624|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|490369||4|3|45
502296291|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-21|2013-08-15|Followup|2012-10-21|2012-10-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|33.8||1|1|1|1|M|White||13|No|Mother|28270|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||34|28278||Married|Self-Employed, Entrepreneur||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011746|502296723|1|0|1|502277214|1|0|1|500475457|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|490485||4|1|45
502179379|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-25|2015-07-31|Followup|2013-07-25|2013-09-13|Declined|Late||||||||4|4|4|4|2|4|3.67|||||||||1|4|4|1|2|4|2.67||||||4|4|4|4|||||||3|3|5|5|4||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||1|2|1.5||||2|2|||||||Red|Project Big|Volunteer: Lost contact with child/agency|60.2||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|Black||34|28269||Single|Student: College||0|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|502179808|31|0|2|502161458|31|0|2|500461681|2||-2||4|3|500004640|500004640|-2||-2|0|10|||9221|5|||1|490654|158340|4|1|45
500185723|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-05|2015-06-25|Followup|2013-09-05|2013-10-20|Complete|Done|4|2|3|2|4|4|3.17|||||||||2|3|3|4|4|4|3.33|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Child: Graduated|81.6||2|2|1|1|M|Black||19||Mother|28214|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|M|Black||36|28214|Bachelors Degree|Single|Tech: Computer/Programmer|28147|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187335|31|0|1|501310677|31|0|1|500284133|2||-2||4|3|||-2||-2|6855|8|||7464|9|||1|490655||4|3|45
502234504|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-28|NaT|Followup|2013-07-28|2013-09-13|Complete|Late|3|2|3|3|3|4|3|4|4|4|4|2|4|3.67|-18.26|4|4|4|4|4|4|4|1|4|4|1|2|4|2.67|49.81|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3|3|5|5|4|25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|1|4|2.5|1|3|2|25|2|2|2|2|0|4|4||||Yellow|Project Big||79.6||1|1|2|2|F|Black||16|No|GrandMother|28208|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|Project Big|Match Support|F|Black||37|28216|Bachelors Degree|Single|Customer Service||8|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500008321|502234935|31|0|2|502129464|31|0|2|500463451|2||500004641||2|2|500004640|500004640|-2||-1|0|4|||11247|3|1204|3|1|490660|155881|4|3|45
502221847|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-27|NaT|Followup|2013-09-27|2013-09-26|Complete|Done|2|1|2|1|3|2|1.83|3|1|2|1|4|2|2.17|-15.67|4|4|4|4|4|4|4|4|4|4|2|4|4|3.67|8.99|4|4|4|4|4|4|4|4|0|3|3|5|5|4|5|4|5|5|4.75|-15.79|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|1|2.33|3|4|4|3.67|-36.51|4|4|4|2|4|3|33.33|2|2|2|2|0|4|4||||Green|Amachi||65.6||2|2|1|1|F|Black||16|Yes|GrandMother|28213|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||24|28027|Some College|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502222278|31|0|2|502654877|31|0|2|500556560|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|490727|154081|4|3|45
502763586|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-06|2017-02-28|Followup|2013-09-06|2013-10-29|Complete|Late|4|1|1|1|4|2|2.17|3|2|3|2|4|3|2.83|-23.32|2|2|4|1|2|3|2.33|2|3|2|2|2|3|2.33|0|4|4|4|4|4|4|4|4|0|4|4|4|5|4.25|3|3|2|2|2.5|70|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|2|2|2|2|100|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|53.7||1|2|5|6|M|Black||16||Mother|28208|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Black|Other African|53|28277||Married|Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502764498|31|0|1|500189754|31|31|1|500632648|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|491029|358930|4|3|45
501604440|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-23|2014-11-19|Followup|2013-07-23|2013-09-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|63.9||1|1|1|1|M|Black||20|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||38|28269||Married|Govt||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501758365|3|0|1|500373108|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|491071||4|1|45
500186435|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-23|2015-08-20|Followup|2013-07-23|2013-09-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|144.9||1|1|1|1|M|Black||20||Mother|28216|One Parent: Female|Unknown||No|Brochure|Media|General Community||Match Support|M|White||45|28226|Bachelors Degree|Married|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187988|31|0|1|500189358|1|0|1|500037395|2||-2||4|1|||-2||-2|51|1|||7496|10|||1|491072||4|1|45
501524313|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-02|2014-04-21|Followup|2013-08-02|2013-09-02|Declined|Done||||||||2|2|3|2|3|3|2.5|||||||||3|3|3|3|3|3|3||||||3|3|3|3|||||||3|3|2|3|2.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||3|3|3||||2|2|||||||Green|2010-2012 OJJDP JJI|Volunteer: Moved|32.6||2|2|1|1|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28208|Bachelors Degree|Single|Finance: Economist|28202|5|6|Recruitment Event|BBBS Board/Staff|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|501524605|31|0|1|502615076|1|0|1|500547406|2||-2||4|1|500005291|500005291|-2|500005291|-2|0|10|||7462|13|||1|491106|4772|4|1|45
502934735|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-19|2013-06-18|Baseline|2012-09-06|2012-11-19|Complete|Done|3|2|3|2|4|4|3|||||||||2|4|3|3|2|4|3|||||||||4|4|3|3.67||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|1|2.5|||||1|1||||4|4||||Yellow||Volunteer: Lost contact with child/agency|6.9||1|1|1|1|F|Black||14|No|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|F|White||51|28031|Some College|Married|Finance: Banking||7|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502936158|31|0|2|502992001|1|0|2|500660486|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|491158|-1|4|3|44
500395038|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-01|2015-02-20|Followup|2013-08-01|2013-09-03|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|102.7||1|1|1|1|M|White||20||Mother|28226|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|M|White||39|28211|Masters Degree|Married|Law: Lawyer|28204|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500395288|1|0|1|500392006|1|0|1|500104016|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|491416||4|1|45
501000843|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-17|2015-09-24|Baseline|2012-09-07|2012-10-17|Complete|Done|4|3|4|2|4|4|3.5|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||2|5|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|1|1.5|||||1|1||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|35.2||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$25,000 to $29,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||26|28269|Bachelors Degree|Single|Business|28262|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|501001116|31|0|2|503106526|31|0|2|500632934|2||-2||4|3|||-2||-2|34|2|||7496|10|||1|491461|-1|4|3|44
502858216|BBBS of Greater Charlotte|Main Office|C|Active|2013-03-19|NaT|Baseline|2012-09-07|2013-03-19|Complete|Done|4|1|4|1|4|4|3|||||||||3|3|4|4|2|4|3.33|||||||||4|4|4|4||||||4|3|2|2|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||47.9||1|1|1|1|M|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||32|29708|Bachelors Degree|Married|Finance||0|9|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020752|502859613|31|0|1|503376842|1|0|1|500687641|2||-2||2|1|||-2||-2|0|10|||7438|1|||1|491466|-1|4|3|44
502108064|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-22|2014-02-06|Followup|2013-07-22|2013-07-23|Complete|Done|4|4|4|2|4|4|3.67|3|4|4|4|4|4|3.83|-4.18|1|4|3|1|2|4|2.5|1|4|3|1|1|3|2.17|15.21|4|4|4|4|4|4|4|4|0|3|4|5|3|3.75|5|5|5|5|5|-25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|3|2.5|1|1|1|150|1|1|1|1|0|4|4||||Yellow||Child: Graduated|42.5||1|1|1|1|F|White||21|No|Father|28277|One Parent: Male|Unknown||No||Relative|General Community||Match Support|F|White||48|28277|High School Graduate|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502108491|1|0|2|502146885|1|0|2|500460150|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|491490|155579|4|3|45
502576641|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-25|NaT|Followup|2013-05-25|2013-06-25|Complete|Done|3|2|3|2|3|3|2.67|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||3|4|3|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|||69.7||1|1|1|1|F|Black||13|No|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|White||41|28207|Masters Degree|Married|Business: Marketing|28202|2|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502577144|31|0|2|502537061|1|0|2|500535114|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|492140||4|3|45
502997224|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-21|2015-04-13|Followup|2013-05-21|2013-08-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|34.7||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||32|28210|Bachelors Degree|Married|Business: Human Resources|28269|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502998689|31|0|2|502939526|31|0|2|500613729|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|492142||4|0|45
502471024|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-09|2016-08-01|Followup|2012-09-09|2012-11-24|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Feels incompatible with child/family|58.7|Y|1|1|1|1|M|Black||13|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||51|28205|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502471471|31|0|1|502685747|1|0|1|500552890|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|492225||4|0|45
501842678|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2015-06-19|Followup|2013-06-27|2013-09-11|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Feels incompatible with child/family|47.7||2|2|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|White||53|28117|Bachelors Degree|Married|Real Estate: Realtor|28031|0|0|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|277|60|598|500000170|500015820|501843047|31|0|1|502335257|1|0|1|500542227|2||-2||4|2|||-2|500000294, 500004901|-2|0|10|||7464|9|||1|492696||4|0|45
503021417|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-11|2015-10-16|Followup|2013-09-11|2013-11-26|Expired|Late||||||||3|3|4|2|3|4|3.17|||||||||3|4|3|2|3|3|3||||||4|4|4|4|||||||4|5|3|4|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|3|2.5||||1|1||||4|4||Yellow||Child/Family: Moved|37.1||1|1|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|White||32|28204|Bachelors Degree|Single|Business: Marketing|29730|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|501428579|31|0|2|503115600|1|0|2|500631553|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|492829|489252|4|0|45
500186960|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-31|2013-08-15|Followup|2013-07-31|2013-08-15|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Time constraint|72.5||2|2|1|1|M|White||19|Yes|Mother|28227|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||40|28105|Some College|Married|Military|28112|11|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188147|1|0|1|500738970|1|0|1|500186719|2||500003586||4|3|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|493385||4|1|45
502247430|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-17|2014-01-23|Followup|2013-08-17|2013-09-27|Declined|Done||||||||3|1|1|1|2|3|1.83|||||||||2|2|3|1|2|2|2||||||4|3|3|3.33|||||||2|3|2|4|2.75||||||||||4|4|4|4|4|4|3|3.86||||||2|4|4|3.33|||||2|1|1.5||||1|1|||||||Yellow||Child: Lost interest|41.2||1|1|1|1|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||63|28078|Bachelors Degree|Married|Medical: Nurse||10|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502247861|31|0|2|502226106|1|0|2|500465539|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|493419|166252|4|1|45
503108699|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-14|2014-08-11|Followup|2013-09-14|2013-11-14|Complete|Late|4|4|3|2|3|4|3.33|3|3|4|1|2|3|2.67|24.72|2|3|3|2|2|3|2.5|2|2|3|2|2|3|2.33|7.3|4|4|3|3.67|4|2|2|2.67|37.45|4|3|4|3|3.5|3|4|3|4|3.5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|3|2.5|4|4|4|-37.5|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|22.9||1|1|1|1|M|White||19|No|Mother|28031|One Parent: Female|$30,000 to $34,999|Y|No||Self|General Community||Match Support|M|White||37|28036|Bachelors Degree|Single|Business: Sales|28117|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503110361|1|0|1|503106216|1|0|1|500631547|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|494022|489246|4|3|45
503158441|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-14|2014-07-03|Followup|2013-09-14|2013-10-09|Complete|Done|4|2|4|1|4|4|3.17|4|3|4|1|4|4|3.33|-4.8|2|4|4|4|2|4|3.33|2|3|4|2|1|4|2.67|24.72|4|4|4|4|4|4|4|4|0|5|4||5||5|3|4|3|3.75||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|1|2.67|3|3|2|2.67|0|3|1|2|4|2|3|-33.33|1|1|2|2|-50|4|4|4|4|0|Red||Volunteer: Moved|21.6||1|1|1|1|F|Black||19|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||27|28202|Bachelors Degree|Single|Business||1|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503160119|31|0|2|503130365|1|0|2|500631432|2||-2||4|3|||-2|500000294|-2|0|5|||7464|9|||1|494087|488914|4|3|45
501750647|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-31|2013-07-25|Followup|2013-08-31|2013-07-25|Declined|Early||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|46.8||2|2|1|1|F|Black||13|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Site||Match Support|F|White||31|28207||Single|Medical: Nurse|28054|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501750989|31|0|2|501584134|1|0|2|500374039|2||-2||4|3|||-1||-2|0|10|||7464|9|||1|494432||4|1|45
502217873|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2013-05-28|Followup|2012-10-27|2012-11-02|Complete|Done|3|1|3|4|2|3|2.67|||||||||2|3|3|2|2|3|2.5|||||||||3|4|3|3.33||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|31||1|1|1|1|F|Hispanic||13|No|Mother|28273|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||28|28273|Bachelors Degree|Single|Medical: Healthcare Worker|28211|0|9|Other|BBBS Board/Staff|Big|General Site|Amachi, mentor2.0 2014, Project Big|Enrollment|277|60|598|500000170|500011746|502218304|3|0|2|502223367|31|0|2|500478268|2||-2||4|3|||-2|500000294, 500004640, 500014506|-1|0|10|||7671|13|||1|494647||4|3|45
502627470|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-12|2014-05-19|Followup|2013-09-12|2013-11-27|Expired|Late||||||||4|4|4|3|2|4|3.5|||||||||2|2|4|1|4|4|2.83||||||3|4|4|3.67|||||||4|5|3|4|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||1|1||||4|4||Green||Volunteer: Lost contact with child/agency|32.2||1|1|1|1|M|Hispanic|Mexican|16|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|Asian||26|28105|Some College|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502628116|3|10|1|502672424|4|0|1|500552887|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|494671|335186|4|0|45
502455004|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-20|NaT|Followup|2013-09-20|2013-09-18|Complete|Done|4|4|4|4|4|4|4|4|2|4|1|1|4|2.67|49.81|2|4|1|2|4|4|2.83|4|4|4|2|4|4|3.67|-22.89|4|4|4|4|4|4|4|4|0|5|4|4|5|4.5|5|5|4|5|4.75|-5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||65.8||1|1|1|1|M|Black|Other African|15|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|29720|Bachelors Degree|Married|Business: Sales|28134|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|31|1|502680045|1|0|1|500553363|2||-2||2|1|500005291|500005291|-2||-2|0|4|||7464|9|||1|495182|336027|4|3|45
500185846|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-28|2014-10-23|Followup|2013-09-28|2013-09-23|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|3|4|5|4.25|||||||4|4|4|4|3|3|3|3.57||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|120.8||1|2|1|2|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||65|28256|Bachelors Degree||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187437|31|0|2|500188764|31|0|2|500038142|2||500003586||4|1|500000294|500000294|-2|500000294|-2|6854|8|||2238|7|||1|495189||4|3|45
503017622|BBBS of Greater Charlotte|Main Office|C|Inactive|2012-09-19|NaT|Followup|2013-09-19|2013-12-02|Declined|Late||||||||3|2|2|2|2|||||||||||3|4|4|3|3|4|3.5||||||4|4|4|4|||||||4|3|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||3|4|4|3.67|||||3|3|3||||2|2||||4|4||Green|||53.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|$30,000 to $34,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|F|White||33|28207|Bachelors Degree|Married|Business||0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|503019155|31|0|2|503095382|1|0|2|500631726|2||-2||3|1|||-2||-2|34|2|||7464|9|||1|495990|489657|4|1|45
503016111|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-30|2017-02-23|Baseline|2012-09-19|2012-09-29|Complete|Done|3|3|4|3|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|1|3.57||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Red||Volunteer: Time constraint|52.8||1|1|1|1|M|Black||14|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Black||32|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503013381|31|0|1|503135600|31|0|1|500636811|2||500003586||4|3||500000294|-2|500000294|-2|0|10|||7496|10|||1|496032|-1|4|3|44
501254255|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-23|2017-02-28|Followup|2013-09-23|2013-10-20|Complete|Done|4|4|4|3|2|2|3.17|||||||||4|4|4|2|3|4|3.5|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|101.2||1|1|1|1|F|Black||14|No|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28205|Masters Degree|Single|Finance: Banking|28217|0|4|Yahoo!|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501254531|31|0|2|501356688|1|0|2|500282157|2||-2||4|1|||-2|500000294|-2|0|10|||32|2|||1|496836||4|3|45
502939293|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-24|2013-11-21|Followup|2013-09-24|2013-10-07|Declined|Done||||||||4|1|4|1|4|4|3|||||||||4|4|4|4|4|4|4||||||4|4|4|4|||||||3|5|4|3|3.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|4|3.5||||2|2||||4|4||Red||Volunteer: Feels incompatible with child/family|13.9||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|F|White||48|28269|Bachelors Degree|Single|Finance: Banking||18|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502940718|31|0|2|502855925|1|0|2|500632744|2||-2||4|3|||-2||-2|0|4|||131|1|||1|497490|472079|4|1|45
502670071|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-26|2014-03-20|Followup|2013-10-26|2013-10-31|Complete|Done|2|4|4|4|4|2|3.33|4|4|4|1|4|4|3.5|-4.86|4|3|4|4|4|3|3.67|4|3|4|4|4|4|3.83|-4.18|4|4|4|4|4|4|4|4|0|5|3|5|5|4.5|5|5|5|5|5|-10|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|3|3|3|3|4|3|3.33|-9.91|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Yellow|Amachi, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|28.8||1|1|1|1|F|Black||16|Yes|Mother|28083|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|Black||36|28269|Masters Degree|Single|Human Services: Youth Worker|28027|2|2|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|502670906|31|0|2|502685522|31|0|2|500557057|2||500003586||4|2|500000294, 500005291|500005291|-2||-2|0|10|||9229|13|||1|498089|341113|4|3|45
501332658|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-01-19|Followup|2013-09-29|2013-10-01|Complete|Done|4|2|4|4|4|4|3.67|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||5|4|4|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Child: Severity of challenges|87.7||1|1|1|1|M|Black||15|Yes|GrandMother|28213|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||46|28227|High School Graduate|Single|Medical: Healthcare Worker|28269|4|0|Coworker|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500020752|501332937|31|0|1|501814288|1|0|1|500384166|2||-2||4|1|500000294|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||7447|3|||1|498110||4|3|45
503039131|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-26|2013-11-21|Baseline|2012-09-25|2013-07-25|Complete|Done|4|2|4|3|3|1|2.83|||||||||3|4|4|4|4|4|3.83|||||||||4|4||||||||4|5|4|5|4.5|||||||3|4|4|4|4|4|4|3.86||||||||||1|4|4|3||||||1|1|1|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|3.9||1|1|2|2|F|Black||18|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||45|28227|Bachelors Degree|Married|Customer Service|28262|18|0|Big For A Day|Special Event|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503040727|31|0|2|503483337|31|0|2|500703051|2||-2||4|3|||-2|500000294|-2|0|10|||16422|8|||1|498146|-1|4|3|44
503041998|BBBS of Greater Charlotte|Main Office|C|Active|2012-10-16|NaT|Baseline|2012-09-26|2012-10-16|Complete|Done|4|2|3|2|3|4|3|||||||||2|3|3|1|2|4|2.5|||||||||3|4|4|3.67||||||4|3|5|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Yellow|||53||1|1|1|1|M|Black||15|No|Mother|28214|One Parent: Female|$45,000 to $49,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28207|Masters Degree|Married|Finance|28273|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503043639|31|0|1|503110820|1|0|1|500638908|2||-2||2|2|||-2||-2|34|2|||7464|9|||1|498892|-1|4|3|44
502920861|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-29|2016-04-22|Baseline|2012-09-27|2012-10-29|Complete|Done|4|2|3|3|4|3|3.17|||||||||4|2|3|4|4|2|3.17|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|3|3.67||||||3|3|3|||||1|1||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|41.8||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||34|28203|Juris Doctorate (JD)|Single|Law: Lawyer||2|11|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502922278|31|0|1|503097126|1|0|1|500639233|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|499329|-1|4|3|44
503034234|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-29|2014-12-17|Baseline|2012-09-27|2012-10-29|Complete|Done|3|4|4|3|1|2|2.83|||||||||2|2|3|2|3|3|2.5|||||||||3|3|2|2.67||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Moved|25.6||1|1|1|1|M|Hispanic||13|No|Mother|28078|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Enrollment|M|White||30|28031|Bachelors Degree|Married|Finance|28036|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503035830|3|0|1|503070689|1|0|1|500639279|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|499356|-1|4|3|44
502264006|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-22|2017-02-26|Followup|2013-09-22|2013-11-21|Declined|Late||||||||2|1|3|1|2|3|2|||||||||1|3|2|2|1|3|2||||||4|4|4|4|||||||4|2|3|4|3.25||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||4|3|3.5||||1|1|||||||Red||Child: Lost interest|77.2||1|1|1|1|F|Hispanic||16|No|Mother|28211|One Parent: Female|Unknown||Yes|Spanish Print|Media|General Community||Match Support|F|Hispanic||38|28202|Bachelors Degree|Single|Tech: Engineer|28202|12|0|Big Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020753|502264438|3|0|2|502274748|3|0|2|500470897|2||-2||4|3|||-2||-2|7063|1|||7456|8|||1|499826|178842|4|1|45
500465511|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-21|2013-10-31|Followup|2013-08-21|2013-09-10|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child: Graduated|86.3||1|1|1|1|M|Black||21|Yes|Mother|28262|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|M|White||54|28210|Masters Degree|Married|Finance: Accountant||0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500527675|1|0|1|500118120|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|4|||2230|7|||1|500353||4|1|45
503016111|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-30|2017-02-23|Followup|2013-09-30|2013-09-30|Complete|Done|4|4|4|2|4|4|3.67|3|3|4|3|4|4|3.5|4.86|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|4|4.75|5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|1|3.57|12.04|4|4|4|4|4|4|3|3.67|8.99|3|3|3|2|2|2|50|1|1|2|2|-50|4|4|4|4|0|Red||Volunteer: Time constraint|52.8||1|1|1|1|M|Black||14|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Black||32|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503013381|31|0|1|503135600|31|0|1|500636811|2||500003586||4|3||500000294|-2|500000294|-2|0|10|||7496|10|||1|500501|496032|4|3|45
503052850|BBBS of Greater Charlotte|Main Office|C|Active|2012-09-30|NaT|Followup|2013-09-30|2013-10-02|Complete|Done|3|2|1|2|4|3|2.5|4|1|2|1|2|3|2.17|15.21|2|3|4|2|1|4|2.67|2|2|2|2|1|3|2|33.5|3|3|3|3|2|3|1|2|50|3|4|5|5|4.25|3|4|2|3|3|41.67|4|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Green|||53.5||1|1|1|1|F|Hispanic||13|No|Mother|28277|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||31|28210|Bachelors Degree|Single|Education: Teacher|29710|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020753|503027860|3|0|2|503028888|1|0|2|500626321|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|500581|476823|4|3|45
503071479|BBBS of Greater Charlotte|Main Office|C|Active|2012-09-30|NaT|Followup|2013-09-30|2013-11-21|Declined|Late||||||||3|3|3|3|2|2|2.67|||||||||3|2|2|3|3|2|2.5||||||4|4|4|4|||||||4|3|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||||||||2|2||||4|4||Green|||53.5||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||28|28269|Some College|Single|Business: Clerical||0|3|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020910|503069483|31|0|1|503051382|1|0|1|500629193|2||-2||2|1|||-2||-2|0|10|||7671|13|||1|500742|485271|4|1|45
500465506|BBBS of Greater Charlotte|Main Office|C|Active|2006-08-21|NaT|Followup|2013-08-21|2013-09-09|Complete|Done|3|1|4|4|3|3|3|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Yellow|Amachi||126.8||1|1|1|1|M|Black||16|Yes|Mother|28262|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||54|28226|Bachelors Degree|Married|Arts, Entertainment, Sports||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500496966|1|0|1|500118121|2||500003586||2|2|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|501159||4|3|45
502721278|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-12|NaT|Followup|2013-10-12|2013-10-10|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|1|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||4|4|4|||||1|1||||3|3||||Green|Amachi, Cabarrus County||65.1||1|1|1|1|M|White||13|Yes|Mother|28025|One Parent: Female|Unknown||Yes||School|General Community|Cabarrus County|Match Support|M|White||47|28025||Single|Tech: Support, Writing|28026|0|2|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501938680|1|0|1|502701096|1|0|1|500560499|2||500003586||2|1|500000294, 500016374|500016374|-2|500016374|-2|0|4|||7464|9|||1|501456||4|3|45
500961274|BBBS of Greater Charlotte|Main Office|C|Active|2007-08-27|NaT|Followup|2013-08-27|2013-09-24|Complete|Done|4|2|4|1|4|4|3.17|||||||||2|4|3|4|4|4|3.5|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||114.6||1|1|2|2|F|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28216|Bachelors Degree|Divorced|Business: Clerical|28204|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500934638|31|0|2|500403000|31|0|2|500186952|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|501812||4|3|45
500474486|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-23|2015-08-18|Followup|2013-08-23|2013-10-18|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|107.8||1|1|1|1|M|Black||20||Mother|28214|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||38|28209|Bachelors Degree|Single|Construction|28247|0|2|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500474735|31|0|1|500491064|31|0|1|500118168|2||-2||4|3|||-2||-2|34|2|||7447|3|||1|502317||4|1|45
500399844|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-20|2017-02-24|Followup|2013-08-20|2013-10-04|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Red||Child: Graduated|114.2||1|2|1|2|F|Black||16||Mother|28208|One Parent: Female|Unknown||No||School|General Site||Match Support|F|White||35|28210|Bachelors Degree|Single|Business: Mgt, Admin|29715|0|0|Radio|Media|Big|General Site||Match Support|277|60|598|500000170|500008321|500400094|31|0|2|500188569|1|0|2|500190707|2||-2||4|3|||-1||-1|0|4|||131|1|||1|502318||4|3|45
502445356|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-04|2016-06-20|Followup|2013-10-04|2013-10-06|Complete|Done|3|2|2|1|3|4|2.5|4|1|3|4|4|4|3.33|-24.92|1|4|4|2|2|4|2.83|4|4|4|4|4|4|4|-29.25|4|4|4|4|4|4|4|4|0|5|4|5|5|4.75|5|4|3|3|3.75|26.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|3|3.67|0|3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Green||Child: Lost interest|44.5||1|2|4|5|F|Black||16|Yes|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community|Amachi|Match Support|F|Black||52|28216|Some College|Divorced|Business: Clerical|28202|16|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|502445803|31|0|2|501026290|31|0|2|500641693|2||-2||4|1||500000294|-2||-2|0|4|||46|2|||1|502503|244170|4|3|45
502172536|BBBS of Greater Charlotte|Main Office|C|Active|2010-10-13|NaT|Followup|2013-10-13|2013-10-12|Complete|Done|3|3|3|3|4|4|3.33|3|2|4|3|1|1|2.33|42.92|3|4|4|3|3|4|3.5|2|4|4|2|2|4|3|16.67|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|4|4|4|4.25|17.65|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|2|3|0|2|2|2|2|0|4|4||||Green|||77.1||1|1|1|1|F|Black||17|No|Mother|28269|Two Parent|Unknown||Yes||Relative|General Community||Match Support|F|Multi-race (Asian & White)||33|28205|Masters Degree|Married|Finance: Economist|28223|7|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502172965|31|0|2|501279665|37|0|2|500475431|2||-2||2|1|||-2||-2|0|3|||129|1|||1|503027|184611|4|3|45
503225805|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-08|2016-05-24|Baseline|2012-10-08|2013-03-08|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|38.5||1|1|1|1|F|White||16|No|Mother|28082|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|F|White||33|28138|Associate Degree|Divorced|Insurance||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503227593|1|0|2|503317460|1|0|2|500680855|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|503767|-1|4|1|44
500867581|BBBS of Greater Charlotte|Main Office|C|Completed|2007-09-28|2014-02-06|Followup|2013-09-28|2013-09-26|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Child: Graduated|76.3||1|1|2|2|M|Black||21|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999||No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||40|28269|Masters Degree|Single|Finance: Accountant|28255|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|500867843|31|0|1|500708515|1|0|1|500195388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|5635|9|||2238|7|||1|504086||4|3|45
502206673|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-13|2015-06-23|Followup|2013-10-13|2013-11-11|Complete|Done|3|4|4|2|3|4|3.33|3|2|3|2|3|4|2.83|17.67|2|4|4|3|3|4|3.33|2|3|3|3|3|3|2.83|17.67|4|4|4|4|4|4|4|4|0|5|4|3|3|3.75|4|5|3|3|3.75|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Red|Amachi|Child: Lost interest|44.3||1|1|1|1|M|Black||17|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||47|28216|Bachelors Degree|Married|Business: Engineer|28255|18|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500013781|502207102|31|0|1|502668179|1|0|1|500557233|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|504104|341305|4|3|45
502593613|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2017-02-28|Followup|2013-08-19|2013-09-03|Declined|Done||||||||3|2||1|2|2||||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|3|3|3.33|||||3|3|3||||2|2||||4|4||Yellow||Volunteer: Lost contact with child/agency|66.4||1|1|1|1|F|Black||16|No|Mother|28208|Two Parent|$35,000 to $39,999|Y|Yes||Relative|General Community||Match Support|F|Hispanic||26|28217|Bachelors Degree|Single|Service: Restaurant||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502594130|31|0|2|502601730|3|0|2|500547881|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|504944|322561|4|1|45
501529924|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2017-02-28|Followup|2013-08-27|2013-10-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|78.1||2|2|1|1|F|Black||15|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||30|28209|Bachelors Degree|Single|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501530213|31|0|2|502199360|1|0|2|500465517|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|504946||4|1|45
500826596|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-28|2013-12-16|Followup|2013-07-28|2013-10-12|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|28.6||3|3|1|1|M|Black||17|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Black||29|28226|Some College|Single|Customer Service|28210|2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500826861|31|0|1|502549323|31|0|1|500544976|2||-2||4|2|500005291||-2|500000294|-2|0|5|||7464|9|||1|506270||4|0|45
502884974|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-09|2014-03-05|Followup|2013-07-09|2013-07-10|Complete|Done|4|1|4|1|3|4|2.83|||||||||2|3|4|1|2|4|2.67|||||||||4|4|4|4||||||5|5|3|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|1|3||||||2|4|3|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|19.8||1|1|1|1|M|Black||13|Yes|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community|Amachi|Match Support|M|White||34|28203|Some College|Single|Business: Marketing|28208|1|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011349|502875571|31|0|1|503036135|1|0|1|500621875|2||-2||4|2||500000294|-2||-2|0|10|||7496|10|||1|506716||4|3|45
501725168|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-31|2013-12-18|Followup|2013-08-31|2013-09-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|51.6||2|2|1|1|F|Multi-Race (None of the above)||15|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28269|Bachelors Degree|Married|Human Services: Non-Profit||2|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017777|501724831|7|0|2|501824761|1|0|2|500381463|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|506788||4|1|45
501347097|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-30|2014-10-16|Followup|2013-07-30|2013-07-22|Complete|Done|4|4|4|2|3|4|3.5|||||||||2|2|3|2|4|4|2.83|||||||||4|4|4|4||||||3|2|4|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|74.5||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||35|28078|Bachelors Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501347376|31|0|2|501099568|1|0|2|500278256|2||-2||4|2|||-2||-2|0|10|||46|2|||1|506852||4|3|45
501872144|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-30|NaT|Followup|2013-07-30|2013-08-01|Complete|Done|3|1|4|4|4|4|3.33|4|4|3|1|3|3|3|11|3|3|3|3|3|3|3|2|3|2|1|2|2|2|50|4|4|4|4|2|3|2|2.33|71.67|3|4|5|5|4.25|2|2|1|2|1.75|142.86|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|3|3|3|1|1|1|200|2|2|2|2|0|4|4||||Green|||79.5||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown|Y|Yes||Relative|General Community||Match Support|M|White||35|28205|Masters Degree|Married|Tech: Engineer|28115|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501872517|31|31|1|502063676|1|0|1|500460156|2||-2||2|1|||-2||-2|0|3|||46|2|||1|506862|155585|4|3|45
502171910|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2015-08-25|Followup|2013-07-30|2013-07-25|Complete|Done|3|4|3|1|2|3|2.67|3|1|2|2|2|3|2.17|23.04|2|4|3|3|1|3|2.67|2|3|3|4|2|4|3|-11|4|4|4|4|4|4|4|4|0|3|4|3|5|3.75|4|3|4|3|3.5|7.14|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|4|3.67|4|4|4|4|-8.25|4|3|3.5|4|4|4|-12.5|2|2|2|2|0|4|4||||Red|Amachi|Volunteer: Time constraint|60.8||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28214|Some College|Married|Medical||3|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502172339|31|0|1|502141964|31|0|1|500460627|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|5|||7464|9|||1|506864|156504|4|3|45
503061519|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-31|2014-08-13|Baseline|2012-10-16|2012-10-31|Complete|Done|3|1|2|1|2|4|2.17|||||||||1|2|4|1||4||||||||||4|4|4|4||||||2|5|5|||||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green||Child/Family: Moved|21.4||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||27|28031|Bachelors Degree|Married|Business: Mgt, Admin|28205|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|503063175|31|0|2|503115965|1|0|2|500646319|2||-2||4|1|||-2||-2|34|2|||7496|10|||1|507929|-1|4|3|44
503041998|BBBS of Greater Charlotte|Main Office|C|Active|2012-10-16|NaT|Followup|2013-10-16|2013-11-04|Complete|Done|3|1|4|1|1|4|2.33|4|2|3|2|3|4|3|-22.33|1|1|3|1|2|3|1.83|2|3|3|1|2|4|2.5|-26.8|3|4|3|3.33|3|4|4|3.67|-9.26|3|3|3|4|3.25|4|3|5|3|3.75|-13.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|1|2|2|4|3|-33.33|1|1|2|2|-50|4|4|4|4|0|Yellow|||53||1|1|1|1|M|Black||15|No|Mother|28214|One Parent: Female|$45,000 to $49,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28207|Masters Degree|Married|Finance|28273|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503043639|31|0|1|503110820|1|0|1|500638908|2||-2||2|2|||-2||-2|34|2|||7464|9|||1|507972|498892|4|3|45
501859854|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-29|2015-09-16|Followup|2013-09-29|2013-11-15|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|59.6||1|1|1|1|F|Black||13|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||28|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501860227|31|0|2|502044100|31|0|2|500469954|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|508458||4|1|45
501000843|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-17|2015-09-24|Followup|2013-10-17|2013-12-01|Complete|Done|3|3|3|3|3|4|3.17|4|3|4|2|4|4|3.5|-9.43|3|4|4|3|3|3|3.33|2|4|3|2|3|3|2.83|17.67|4|4|4|4|4|4|4|4|0|4|4|3|3|3.5|2|5|3|3|3.25|7.69|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|4|3|3.33|0|3|2|2.5|2|1|1.5|66.67|2|2|1|1|100|4|4|4|4|0|Red||Child/Family: Lost contact with volunteer/agency|35.2||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$25,000 to $29,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||26|28269|Bachelors Degree|Single|Business|28262|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|501001116|31|0|2|503106526|31|0|2|500632934|2||-2||4|3|||-2||-2|34|2|||7496|10|||1|508508|491461|4|3|45
502034298|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-19|2015-08-31|Followup|2013-10-19|2013-10-17|Complete|Done|4|4|4|4|4|4|4|3|4|4|2|4|4|3.5|14.29|4|4|4|3|4|4|3.83|2|4|3|4|3|4|3.33|15.02|4|4|4|4|4|4|4|4|0|4|5|5|4|4.5|5|5|5|4|4.75|-5.26|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|3|3.67|8.99|2|3|2.5|2|4|3|-16.67|2|2|1|1|100|4|4||||Red||Volunteer: Time constraint|34.4||2|3|4|6|M|White||16|Yes|Mother|28146|One Parent: Female|Unknown||Yes||School|General Community|Amachi|Match Support|M|White||41|28078|Bachelors Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502034697|1|0|1|500188638|1|0|1|500631278|2||-2||4|3||500000294|-2|500000294|-2|0|4|||7464|9|||1|510234|27853|4|3|45
501253195|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-24|NaT|Followup|2013-10-24|2013-10-20|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||100.7||1|1|2|2|M|Black||15|Yes|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28203|Masters Degree|Single|Medical: Doctor, Provider|28211|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501253471|31|0|1|500395148|1|0|1|500282924|2||500003586||2|1|500000294||-2||-2|0|10|||7464|9|||1|510241||4|3|45
500545326|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2016-09-02|Followup|2013-10-29|2013-11-13|Complete|Done|4|1|2|2|3|4|2.67|||||||||1|4|4|2|2|4|2.83|||||||||4|4|4|4||||||4|1|5|1|2.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|118.1|Y|1|1|1|1|M|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|Black||55|28214||Married|Clergy||12|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|1|500697845|31|0|1|500134545|2||-2||4|3|||-2||-2|0|10|||2238|7|||1|510384||4|3|45
500187075|BBBS of Greater Charlotte|Main Office|C|Completed|2004-09-21|2014-01-16|Followup|2013-09-21|2013-10-23|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|3|4|3.67||||||2|4|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|111.8||1|1|6|6|F|Black||21||Mother|28205|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|White||38|28209|Bachelors Degree|Single|Human Services: Non-Profit||0|0|Recruitment Event|Self|Big|General Site||Match Support|277|60|598|500000170|500012459|500188223|31|0|2|500189550|1|0|2|500037643|2||-2||4|1|||-2||-1|0|10|||7458|9|||1|511345||4|3|45
501989028|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-22|2016-08-30|Followup|2013-10-22|2013-11-18|Complete|Done|1|4|4|4|4|4|3.5|4|1|4|1|4|4|3|16.67|1|4|4|3|3|4|3.17|2|3|4|3|4|4|3.33|-4.8|4|4|4|4|4|3|4|3.67|8.99|4|3|5|5|4.25|5|4|4|4|4.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|2|3|2.5|60|2|2|2|2|0|4|4|4|4|0|Yellow||Child/Family: Moved|46.3||2|2|1|1|M|Black||15|No|Mother|28273|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28273|Juris Doctorate (JD)|Single|Law: Lawyer||0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502425720|31|0|1|503039778|31|0|1|500641725|2||-2||4|2||500005291|-2||-2|6855|8|||7496|10|635|1|1|511361|251884|4|3|45
503052841|BBBS of Greater Charlotte|Main Office|C|Active|2013-01-24|NaT|Baseline|2012-10-22|2013-01-24|Complete|Done|3|3|4|4|3|4|3.5|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|5|5|3|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||49.7||1|1|1|1|F|Hispanic||18|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||24|28104|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503027860|3|0|2|503122069|1|0|2|500660497|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|511402|-1|4|3|44
500931662|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-07|NaT|Followup|2013-09-07|2013-11-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||114.3||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$60,000 to $74,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||58|28270|Bachelors Degree|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500931932|31|0|1|500894084|1|0|1|500193824|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|511880||4|0|45
502510347|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-31|2016-08-30|Followup|2013-10-31|2013-12-02|Declined|Done||||||||4|1|2|1|4|4|2.67|||||||||1|4|2|2|2|2|2.17||||||4|4|4|4|||||||3|4|2|4|3.25||||||||||4|4|4|4|4|4|2|3.71||||||3|2|1|2|||||4|2|3||||1|1||||4|4||Green|2010-2012 OJJDP JJI|Child: Graduated|58||1|1|1|1|F|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28262|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502510796|31|0|2|502677833|31|0|2|500557844|2||-2||4|1|500005291|500005291|-2||-2|0|5|||7464|9|||1|512006|310349|4|1|45
502000252|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-22|NaT|Followup|2013-08-22|2013-09-02|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||78.8||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020910|502000651|31|0|1|502127058|1|0|1|500465318|2||-2||2|1|||-2||-2|0|10|||130|1|||1|512007||4|1|45
502602958|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-11|2017-02-23|Followup|2013-09-11|2013-11-26|Expired|Late||||||||4|1|1|2|3|4|2.5|||||||||4|3|4|4|4|4|3.83||||||4|4|4|4|||||||5|3|5|5|4.5||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||2|3|2.5||||2|2||||4|4||Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|65.4||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||52|28207|Masters Degree|Married|Business|28202|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501480402|31|0|1|502578040|1|0|1|500552390|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|512028|333955|4|0|45
500483980|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-01|2014-03-24|Followup|2013-09-01|2013-10-16|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|90.7||1|1|2|2|M|Black||21||Mother|28227|One Parent: Female|$10,000 to $14,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||71|28270||Single|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500484231|31|0|1|500423426|31|0|1|500120592|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|512562||4|1|45
502436202|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2015-07-13|Followup|2013-09-02|2013-10-17|Declined|Done||||||||3|2|2|1|3|3|2.33|||||||||3|3|3|4|2|4|3.17||||||4|4|4|4|||||||2|5|5|5|4.25||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||2|4|3||||1|1||||4|4||Green||Child: Graduated|46.3||1|1|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|Masters Degree|Single|Finance: Banking||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502436645|31|0|1|502642999|1|0|1|500549046|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|512564|327937|4|1|45
500970495|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-10|2017-03-09|Followup|2013-09-10|2013-11-25|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|101.9||3|3|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$35,000 to $39,999||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black|Other African|44|28212||Single|Consultant||1|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500970766|31|0|2|500965698|31|31|2|500285645|2||-2||4|2|||-2||-2|7294|13|||46|2|||1|512577||4|0|45
501309634|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-12|NaT|Followup|2013-09-12|2013-10-24|Complete|Done|2|4|4|4|4|4|3.67|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi||102.1||1|1|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||46|27704|Associate Degree|Divorced|Medical: Admin||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501309912|31|0|2|501046221|31|0|2|500281317|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7462|13|||1|512878||4|3|45
500382177|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-18|2015-08-25|Followup|2013-09-18|2013-11-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|107.2||1|1|2|2|M|Black||16||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||43|28215|Bachelors Degree|Single|Finance: Banking|28262|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|500382427|31|0|1|500188566|31|0|1|500122093|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|512879||4|1|45
501604446|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-19|NaT|Followup|2013-09-19|2013-12-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|2010-2012 OJJDP JJI||65.9||2|2|1|1|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28213|Bachelors Degree|Married|Tech: Support, Writing|28273|11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|502664359|31|0|1|500555050|2||-2||2|1|500005291|500005291|-2||-2|0|10|||7462|13|||1|512881||4|0|45
502064627|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-20|NaT|Followup|2013-08-20|2013-10-10|Complete|Late|3|2|4|2|3|4|3|2|2|4|2|3|4|2.83|6.01|2|3|3|2|3|3|2.67|3|3|4|3|2|4|3.17|-15.77|4|4|4|4|4|3|2|3|33.33|5|4|3|3|3.75|5|3|3|4|3.75|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|3|2|3|2.67|49.81|2|3|2.5|2|3|2.5|0|2|2|1|1|100|4|4||||Green|||78.9||1|1|2|2|M|Black||16|No|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|502065051|31|0|1|500773055|3|14|1|500462574|2||-2||2|1|||-2||-2|0|10|||46|2|||1|513771|159373|4|3|45
503026933|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-27|2013-07-31|Baseline|2012-10-25|2012-12-27|Complete|Done|2|2|3|2|3|3|2.5|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||2|2|3|3|2.5|||||||3|4|4|4|4|4|3|3.71||||||||||2|3|3|2.67||||||2|2|2|||||1|1||||4|4||||Red||Child/Family: Feels incompatible with volunteer|7.1||2|2|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28216|Two Parent|$35,000 to $39,999|Y|Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|Black||33|28216|Bachelors Degree|Single|Finance: Banking|28269|6|10|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503028507|38|0|2|503111607|31|0|2|500660471|2||-2||4|3||500011312|-2||-2|0|10|||7496|10|||1|513783|-1|4|3|44
500826594|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-21|2016-06-15|Followup|2013-08-21|2013-11-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|105.8||1|1|1|1|M|Black||18|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Some Other Race||36|28209|||Business: Sales||0|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|1|500920342|41|0|1|500185735|2||-2||4|1|||-2||-2|0|5|||6450|12|||1|514430||4|0|45
502129650|BBBS of Greater Charlotte|Main Office|C|Active|2012-10-26|NaT|Followup|2013-10-26|2013-10-24|Complete|Done|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|4|4|4|4|3.67|1|4|3|4|1|4|2.83|29.68|4|4|4|4|4|4|4|4|0|5|5|4|5|4.75|5|4|5|4|4.5|5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4||||Green|Cabarrus County||52.6||2|2|2|2|F|Black||17|No|GrandMother|28027|Grandparents|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|Black||42|28213|Bachelors Degree|Single|Finance: Banking|28202|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502130079|31|0|2|502598777|31|0|2|500646243|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|10|||7464|9|||1|514663|220242|4|3|45
502969236|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-14|2013-08-30|Followup|2013-05-14|2013-06-07|Complete|Done|3|2|3|2|3|4|2.83|||||||||4|4|4|4|4|3|3.83|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|15.5||2|2|1|1|F|Some Other Race||13||Mother|28277|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||34|28277|Bachelors Degree||Medical: Nurse||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|502970672|41|0|2|502938930|1|0|2|500612989|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|515403||4|3|45
501597228|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-04|NaT|Followup|2013-09-04|2013-10-03|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi||90.3||1|1|1|1|F|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||40|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28204|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501597548|31|0|2|501397328|31|0|2|500379964|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|515461||4|3|45
501725162|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2016-10-14|Followup|2013-10-29|2013-11-04|Complete|Done|3|3|2|1|4|4|2.83|4|1|2|1|4|4|2.67|5.99|2|2|2|3|4|2|2.5|3|4|2|3|3|3|3|-16.67|3|2|3|2.67|1|4|4|3|-11|2|3|3|3|2.75|5|1|5|5|4|-31.25|4|4|4|4|4|4|2|3.71|4|4|4|4|4|4|3|3.86|-3.89|2|4|2|2.67|4|4|2|3.33|-19.82|4|3|3.5|4|3|3.5|0|1|1|2|2|-50|4|4||||Green||Agency: Challenges with program/partnership|83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501724831|39|0|1|501833178|1|0|1|500394157|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|515608|16143|4|3|45
503034234|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-29|2014-12-17|Followup|2013-10-29|2013-10-09|Complete|Early|3|4|4|4|1|4|3.33|3|4|4|3|1|2|2.83|17.67|2|4|4|2|1|4|2.83|2|2|3|2|3|3|2.5|13.2|4|4|4|4|3|3|2|2.67|49.81|4|3|4|5|4|4|4|5|5|4.5|-11.11|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|3|3.67|8.99|2|3|2.5|2|2|2|25|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|25.6||1|1|1|1|M|Hispanic||13|No|Mother|28078|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Enrollment|M|White||30|28031|Bachelors Degree|Married|Finance|28036|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503035830|3|0|1|503070689|1|0|1|500639279|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|515837|499356|4|3|45
500185812|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-29|2016-05-26|Followup|2013-10-29|2013-12-13|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|42.9||2|3|2|3|F|Black||18|Yes|Mother|28210|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community|Amachi|Match Support|F|White||41|28214|Bachelors Degree|Single|Human Services: Non-Profit||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187400|31|0|2|500188912|1|0|2|500648551|2||-2||4|1||500000294|-2||-2|0|10|||7464|9|||1|515874||4|1|45
502920861|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-29|2016-04-22|Followup|2013-10-29|2013-12-13|Complete|Done|4|3|3|2|4|4|3.33|4|2|3|3|4|3|3.17|5.05|4|3|4|4|3|4|3.67|4|2|3|4|4|2|3.17|15.77|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|3|5|5|4.5|11.11|4|4|4|4|4|4|3|3.86|4|4|4|4|4|3|3|3.71|4.04|4|4|4|4|4|4|3|3.67|8.99|2|4|3|3|3|3|0|2|2|1|1|100|4|4|4|4|0|Yellow||Child/Family: Lost contact with volunteer/agency|41.8||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||34|28203|Juris Doctorate (JD)|Single|Law: Lawyer||2|11|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502922278|31|0|1|503097126|1|0|1|500639233|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|515903|499329|4|3|45
501224287|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-30|2014-01-23|Followup|2013-10-30|2014-01-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child: Lost interest|62.8||1|1|1|1|M|Black||19|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||43|28262|Bachelors Degree|Married|Customer Service|28211|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501224558|31|0|1|501343190|31|0|1|500298289|2||-2||4|3|500000294|500000294|-2|500000294|-2|5635|9|||2230|7|||1|516896||4|0|45
500970267|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-29|NaT|Followup|2013-09-29|2013-11-15|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||77.5||1|1|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||61|28204||Divorced|Self-Employed, Entrepreneur||0|0|Billboard|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|2|502084649|1|0|2|500468192|2||500003586||2|1|500000294|500000294|-2|500000294|-2|5635|9|||125|1|||1|516916|174196|4|1|45
501372080|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-31|2016-04-22|Followup|2013-10-31|2013-11-18|Complete|Done|4|2|2|2|3|4|2.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child/Family: Moved|41.7||2|2|2|2|M|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community||Match Support|M|White||31|28269|Masters Degree|Single|Insurance|28262|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|501372359|31|0|1|502500246|1|0|1|500640327|2||-2||4|2|||-2||-2|0|3|||7496|10|||1|517148||4|3|45
502926905|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-31|2014-09-18|Followup|2013-10-31|2013-10-28|Complete|Done|3|4|3|2|3|3|3|2|4|4|4|4|4|3.67|-18.26|4|4|4|3|3|4|3.67|2|3|3|2|2|3|2.5|46.8|4|4|4|4|4|3|3|3.33|20.12|3||4|5||2|3|3|2|2.5||4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|4|4|4|4|3|3.67|8.99|3|3|3|3|4|3.5|-14.29|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Feels incompatible with child/family|22.6||1|1|1|1|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||32|28216|Bachelors Degree|Single|Tech: Support, Writing|28117|1|9|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502928325|31|0|2|503096831|31|0|2|500635818|2||-2||4|2|||-2||-2|7294|13|||7438|1|||1|517308|415449|4|3|45
502698998|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2014-03-13|Followup|2013-11-11|2013-12-20|Declined|Done||||||||3|2|2|1|3|3|2.33|||||||||3|2|3|3|3|3|2.83||||||4|4|4|4|||||||3|4|4|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||4|3|3.5||||2|2||||4|4||Yellow||Child/Family: Lost contact with volunteer/agency|28||1|1|1|1|F|Black||18|No|GrandMother|28211|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28203|Masters Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500012459|502699843|31|0|2|502692148|1|0|2|500564380|2||-2||4|2||500005291|-2||-2|0|4|||7464|9|||1|517670|350301|4|1|45
503061519|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-31|2014-08-13|Followup|2013-10-31|2013-11-13|Complete|Done|4|4|4|1|1|4|3|3|1|2|1|2|4|2.17|38.25|1|1|4|1|4|1|2|1|2|4|1||4|||3|3|3|3|4|4|4|4|-25|3|4|2|3|3|2|5|5||||4|4|4|4|3|4|4|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|3|3.67|8.99|4|4|4|2|4|3|33.33|2|2|2|2|0|4|4|4|4|0|Green||Child/Family: Moved|21.4||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||27|28031|Bachelors Degree|Married|Business: Mgt, Admin|28205|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|503063175|31|0|2|503115965|1|0|2|500646319|2||-2||4|1|||-2||-2|34|2|||7496|10|||1|517783|507929|4|3|45
502728419|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-06|2013-08-22|Followup|2013-02-06|2013-02-26|Comprehension|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|18.5||2|2|1|1|M|Black||13|No|Mother|28214|One Parent: Female|$50,000 to $59,999||No|Big|Neighbor/Friend|General Community|PERL 2014-2016|Match Support|M|White||50|28105|Bachelors Degree|Married|Finance|28217|12|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502729316|31|0|1|502889543|1|0|1|500594026|2||-2||4|3||500014681|-2||-2|6854|8|||7496|10|||1|517966||4|2|45
502205848|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-18|NaT|Followup|2013-08-18|2013-11-02|Expired|Late||||||||3|4|3|2|4|4|3.33|||||||||3|2|3|4|3|3|3||||||4|4|4|4|||||||4|4|5|4|4.25||||||||||4|4|4|4|3|4|4|3.86||||||4|4|3|3.67|||||2|4|3||||1|1||||4|4||Green|2010-2012 OJJDP JJI||66.9||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Juris Doctorate (JD)|Single|Student: College|28208|0|0||Law Student Association|Big|General Community||Match Support|277|60|598|500000170|500020753|502206277|31|0|1|502624702|1|0|1|500549350|2||-2||2|1|500005291|500005291|-2||-2|0|10|||0|15|||1|518525|328511|4|0|45
503063881|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-30|2015-01-14|Baseline|2012-11-02|2012-11-30|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Yellow||Volunteer: Moved|25.5||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||34|28202|Associate Degree|Single|Medical: Healthcare Worker||6|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503065564|31|0|2|503125383|1|0|2|500656877|2||-2||4|2|||-2||-2|0|10|||46|2|||1|518880|-1|4|3|44
500868942|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-20|NaT|Followup|2013-09-20|2013-12-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||113.8|Y|1|1|1|1|M|Black||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|M|White||54|28207||Married|Business: Sales||0|0|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500869211|31|0|1|500947018|1|0|1|500195082|2||-2||2|1|||-2||-2|0|10|||7458|9|||1|519494||4|0|45
501771263|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-02-28|Followup|2013-09-29|2013-12-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|89||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||31|28262|Bachelors Degree|Single|Medical: Admin|28216|0|8|Recruitment Event|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501741899|31|0|2|501622704|31|0|2|500379993|2||-2||4|1|||-2||-2|0|10|||7443|2|||1|519500||4|0|45
502245129|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-22|NaT|Followup|2013-08-22|2013-09-25|Complete|Done|3|3|4|2|4|3|3.17|4|3|4|2|3|3|3.17|0|2|2|2|1|1|3|1.83|1|4|3|2|4|3|2.83|-35.34|4|3|3|3.33|4|3|2|3|11|3|4|5|5|4.25|5|4|3|2|3.5|21.43|4|4|4|4|4|3|4|3.86|4|3|4|3|2|4|3|3.29|17.33|2|4|2|2.67|4|4|3|3.67|-27.25|2|2|2|4|3|3.5|-42.86|2|2|1|1|100|4|4|4|4|0|Green|Amachi||66.8||1|1|1|1|M|Multi-race (Black & Hispanic)||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||28|28262|High School Graduate|Single|Laborer||0|8|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|502245570|38|0|1|502670839|31|0|1|500551050|2||-2||2|1|500000294||-2||-2|0|10|||7671|13|||1|519875|331272|4|3|45
501938282|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-17|NaT|Followup|2013-11-17|2013-11-16|Complete|Done|4|4|4|4|1|4|3.5|||||||||1|4|3|1|2|3|2.33|||||||||4|4|4|4||||||1|5|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green|Amachi, Cabarrus County||75.9||1|1|1|1|F|White||14|Yes|Mother|28025|Two Parent|Unknown|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||63|28027|High School Graduate|Married|Self-Employed, Entrepreneur|28027|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501938680|1|0|2|502356100|1|0|2|500493871|2||500016307||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|520829||4|3|45
502976039|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-16|2013-02-28|Baseline|2012-11-09|2012-11-16|Complete|Done|4|2|3|4|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Red||Child/Family: Infraction of match rules/agency policies|3.4||1|1|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|White||29|28205|Some College|Single|Medical||2|0|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500004169|502977487|31|0|1|503150561|1|0|1|500658198|2||-2||4|3|||-2||-2|0|10|||7438|1|||1|522750|-1|4|3|44
500185907|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2015-02-18|Followup|2013-10-29|2013-12-11|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|99.7||2|3|1|1|F|Black||19|Yes|Mother|28262|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||48|28212||Single|Medical: Healthcare Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187470|31|0|2|500697782|31|0|2|500134557|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|522867||4|3|45
500871683|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-01|2016-02-22|Followup|2013-10-01|2013-11-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|100.7||1|1|1|1|M|Black||19|Yes|Aunt|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|M|White||46|28209|Masters Degree|Single|Self-Employed, Entrepreneur|28209|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500871952|31|0|1|500933829|1|0|1|500199601|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|522869||4|1|45
501014187|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-07|NaT|Followup|2013-11-07|2013-11-22|Complete|Done|1|4|4|4|3|3|3.17|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||100.2||2|2|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||48|28205|Bachelors Degree|Living w/ Significant Other|Human Services: Non-Profit|28205|3|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501404007|1|0|2|500306699|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7671|13|||1|523375||4|3|45
500826592|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-08|2016-10-18|Followup|2013-10-08|2013-12-12|Complete|Late|3|4|4|4|3|4|3.67|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||2|2||||4|4||||Green||Child: Graduated|84.3||3|3|1|1|F|Black||20|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|F|White||33|28277|Bachelors Degree|Living w/ Significant Other|Unknown|28209|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|2|501314246|1|0|2|500382768|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|523408||4|3|45
500186133|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-14|2016-06-28|Followup|2013-10-14|2013-11-18|Complete|Done|3|2|3|2|3|3|2.67|||||||||2|3|3|3|4|4|3.17|||||||||4|4|4|4||||||4|3|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|140.5||1|1|1|1|M|White||18||Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||51|28262|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500187724|1|0|1|500188930|1|0|1|500036930|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|523889||4|3|45
502255225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-08|2016-08-26|Followup|2013-11-08|2014-01-10|Complete|Late|4|1|2|1|3|4|2.5|2|2|2|4|1|4|2.5|0|2|3|3|3|2|4|2.83|2|3|3|2|2|3|2.5|13.2|4|3|3|3.33|4|3|3|3.33|0|5|3|5|4|4.25|5|3|5|3|4|6.25|4|1|4|4|3|4|2|3.14|4|3|4|4|4|4|4|3.86|-18.65|4|4|4|4|4|4|4|4|0|3|4|3.5|1|1|1|250|2|2|1|1|100|4|4||||Red||Volunteer: Moved|69.6||1|1|1|1|M|Hispanic||15||Mother|28212|One Parent: Female|Unknown||No|Spanish Radio|Media|General Community||Match Support|M|White||33|28226|Bachelors Degree|Single|Education: Teacher||3|0|Spanish Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502255655|3|0|1|502312682|1|0|1|500487118|2||-2||4|3|||-2||-2|7068|1|||11662|1|||1|523901|199091|4|3|45
502353937|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-22|NaT|Followup|2013-11-22|2013-11-21|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|4|3|3|4|3.17|||||||||4|4|4|4||||||1|5|5|5|4|||||||4|4|4|4|4|4|2|3.71||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||75.8||1|1|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||31|29605|Bachelors Degree|Single|Business: Human Resources|29615|1|0|Local TV|Media|Big|General Community|Project Big AND Amachi|Match Support|277|60|598|500000170|500018851|502354375|31|0|2|501672025|1|0|2|500487322|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500004901|-2|0|4|||7438|1|||1|523903||4|3|45
502869635|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-13|2014-08-21|Followup|2013-11-13|2013-11-11|Complete|Done|3|4|4|4|4|4|3.83|4|4|4|4|3|4|3.83|0|3|4|3|4|1|4|3.17|3|3|4|3|3|3|3.17|0|4|4|4|4|4|4|4|4|0|3|3|4|4|3.5|4|4|5|3|4|-12.5|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|3|3|3|11|2|2|2|4|3|3.5|-42.86|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Moved|21.2||1|1|1|1|F|Black||17|No|Mother|28206|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community||Match Support|F|Black||34|28210|Bachelors Degree|Single|Business: Marketing||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502871029|31|0|2|503099564|31|0|2|500649374|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|524300|483786|4|3|45
502601023|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-31|2016-08-11|Followup|2013-08-31|2013-08-27|Complete|Done|2|2|4|2|2|2|2.33|3|2|3|1|3|4|2.67|-12.73|4|4|4|4|3|3|3.67|3|3|4|2|2|3|2.83|29.68|4|4|4|4|4|4|4|4|0|4|3|4|4|3.75|3|3|4|5|3.75|0|4|4|3|4|4|3|3|3.57|4|2|4|4|3|4|3|3.43|4.08|3|4|3|3.33|3|4|2|3|11|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child: Graduated|59.4||1|1|1|1|F|Black||19||Mother|28216|Two Parent|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||51|28277|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502601540|31|0|2|502546883|1|0|2|500550809|2||-2||4|1|500005291|500005291|-2||-2|6854|8|||7464|9|||1|525510|331012|4|3|45
502787401|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-30|2016-10-30|Baseline|2012-11-15|2013-04-29|Complete|Done|4|3|4|4|1|3|3.17|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|42||1|1|1|1|F|Black||16|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||41|28105|High School Graduate|Divorced|Business: Mgt, Admin|28207|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502788587|31|0|2|503122442|1|0|2|500692539|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|525811|-1|4|3|44
501237971|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-17|2016-03-03|Followup|2013-11-17|2013-11-16|Complete|Done|4|3|4|3|3|3|3.33|||||||||2|3|3|3|2|4|2.83|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Moved|39.5||2|2|3|3|F|Black||18|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||41|28269|||Business: Human Resources|28206|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503287812|31|0|2|501598429|31|0|2|500649363|2||-2||4|1||500000294|-2||-2|0|10|||7464|9|||1|526992||4|3|45
502273093|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-01|2015-03-31|Followup|2013-10-01|2013-11-15|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|53.9||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||37|28277|PHD|Single|Medical: Healthcare Worker||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502273525|31|0|2|502252422|31|0|2|500471568|2||-2||4|1|||-2|500000294|-2|0|4|||7496|10|||1|527621||4|1|45
502097794|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-20|NaT|Followup|2013-01-20|2013-01-31|Complete|Done|4|1|4|2|3|3|2.83|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||73.8||1|1|1|1|M|Black||13|No|Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28031|Bachelors Degree|Single|Business: Engineer|28036|0|8|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502098218|31|0|1|502425119|1|0|1|500510881|2||-2||2|1|||-2|500000294, 500004640|-2|34|2|||46|2|||1|528635||4|3|45
500252077|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-24|2016-01-20|Followup|2013-11-24|2013-11-21|Complete|Done|3|1|2|1|4|3|2.33|||||||||2|3|4|2|4|4|3.17|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|85.8||3|3|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Tech: Computer/Programmer||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501750989|31|0|1|501365749|1|0|1|500317108|2||500003586||4|3|500000294|500000294|-2||-2|7295|11|||46|2|||1|529037||4|3|45
502915950|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-02|2013-09-12|Followup|2013-04-02|2013-04-30|Complete|Done|1|4|2|4|3|3|2.83|||||||||2|3|4|2|4|4|3.17|||||||||3|4|3|3.33||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green||Volunteer: Moved|17.3||1|1|1|1|F|White||13|No|Mother|28031|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|F|White||34|28031|Masters Degree|Single|Education||3|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011349|502917364|1|0|2|502913149|1|0|2|500602723|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|529186||4|3|45
502471024|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-09|2016-08-01|Followup|2013-09-09|2013-10-10|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|3|3.67||||||4|5|4|3|4|||||||4|4|4|4|3|3|4|3.71||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green||Volunteer: Feels incompatible with child/family|58.7|Y|1|1|1|1|M|Black||13|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||51|28205|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502471471|31|0|1|502685747|1|0|1|500552890|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|529310||4|3|45
502859187|BBBS of Greater Charlotte|Main Office|C|Active|2012-11-24|NaT|Followup|2013-11-24|2014-01-08|Complete|Done|3|3|4|2|3|3|3|2|2|4|2|4|4|3|0|3|4|3|3|3|4|3.33|2|3|3|3|3|4|3|11|4|4|4|4|4|4|4|4|0|3|3|3|3|3|4|5|3|3|3.75|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|4|4|4|4|-16.75|3|2|2.5|4|4|4|-37.5|2|2|2|2|0|4|4|4|4|0|Green|VOL - PreMatch||51.7||2|2|1|1|F|Black||15|No|GrandMother|28205|Grandparents|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|White||31|28209|Associate Degree|Married|Retail: Mgt|28134|4|3|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500187987|31|0|2|503090888|1|0|2|500658723|2||-2||2|1|500007920||-2||-2|0|10|||9221|5|||1|529317|400467|4|3|45
501123191|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-20|2015-12-21|Followup|2013-10-20|2014-01-03|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|62||2|2|1|1|F|Black||15|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||48|28210|Some College|Single|Human Services||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500915629|31|0|2|502153920|1|0|2|500478644|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|530133||4|1|45
502499851|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2015-07-07|Followup|2013-11-11|2013-11-11|Complete|Done|3|3|4|3|3|2|3|3|1|1|1|2|2|1.67|79.64|3|3|4|3|4|4|3.5|4|4|4|2|2|4|3.33|5.11|4|4|4|4|4|4|4|4|0|3|5|4|5|4.25|5|5|5|4|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|3|3.33|20.12|4|4|4|2|4|3|33.33|2|2|2|2|0|4|4|4|4|0|Red||Agency: Concern with Volunteer re: child safety|43.8||1|1|1|1|M|White||18|No|Mother|28210|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||39|28210|Masters Degree|Single|Finance|28106|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|502500300|1|0|1|502690262|1|0|1|500562789|2||-2||4|3|||-2||-2|0|10|||46|2|||1|530351|348364|4|3|45
500186106|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-18|2015-08-13|Followup|2013-10-18|2013-11-01|Complete|Done|4|3|4|3|4|4|3.67|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Graduated|93.8||2|2|1|1|F|Black||20||Mother|28217|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||35|28211|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187698|31|0|2|500778380|1|0|2|500202993|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|530369||4|3|45
500936718|BBBS of Greater Charlotte|Main Office|C|Completed|2007-12-20|2016-06-16|Followup|2013-12-20|2014-03-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Agency: Challenges with program/partnership|101.9||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28210|Bachelors Degree|Married|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500017732|500915629|31|0|1|501027885|1|0|1|500224574|2||-2||4|1|||-2|500014505, 500015184|-1|34|2|||46|2|||1|530373||4|0|45
503163476|BBBS of Greater Charlotte|Main Office|C|Active|2012-11-30|NaT|Baseline|2012-11-27|2012-11-30|Complete|Done|3|1|1|1|1|3|1.67|||||||||2|3|4|2|3|3|2.83|||||||||3|4|4|3.67||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|||51.5||1|1|1|1|M|Black||13|No|Mother|28269|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|Black||32|28217|Masters Degree|Single|Consultant||0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503165154|31|0|1|503119713|31|0|1|500663695|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|530536|-1|4|3|44
503026286|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2017-02-26|Baseline|2012-11-28|2013-01-31|Complete|Done|3|3|4|4|3|3|3.33|||||||||3|3|3|3|3|2|2.83|||||||||4|4|4|4||||||5|2|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|48.9||1|1|1|1|M|Hispanic||17|No|Mother|28277|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Asian||30|28277|Bachelors Degree|Single|Finance||1|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503027860|3|0|1|503259120|4|0|1|500674960|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|530932|-1|4|3|44
502674024|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-07|2016-05-17|Followup|2013-12-07|2013-12-12|Complete|Done|3|4|4|4|4|4|3.83|4|4|4|3|4|4|3.83|0|2|4|4|4|4|3|3.5|2|4|4|4|4|3|3.5|0|4|4|4|4|4|4|4|4|0|2|5|5|4|4|4|4|4|3|3.75|6.67|2|3|4|4|4|3|3|3.29|4|4|4|4|4|4|3|3.86|-14.77|3|2|3|2.67|3|4|3|3.33|-19.82|2|4|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Green||Child: Lost interest|53.3||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Sales||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018851|502674852|31|0|2|502660051|1|0|2|500581910|2||-2||4|1||500005291|-2||-2|0|10|||7496|10|||1|530942|374331|4|3|45
502419933|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-07|2014-09-04|Followup|2013-12-07|2014-01-23|Complete|Late|3|4|3|3|4|4|3.5|3|2|3|3|3|3|2.83|23.67|2|4|4|2|2|4|3|3|3|3|2|3|4|3|0|4|4|4|4|4|4|4|4|0|3|3|4|4|3.5|4|4|4|4|4|-12.5|4|4|4|4|4|4|3|3.86||4|4|4|4|4|4|||4|4|4|4|4|4|4|4|0|3|2|2.5|4|4|4|-37.5|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Time constraint|32.9||2|2|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$40,000 to $44,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||58|28031|Bachelors Degree|Living w/ Significant Other|Business: Mgt, Admin||22|0|Big Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500011349|502371107|31|0|1|502669194|1|0|1|500571419|2||-2||4|2||500005291|-2||-2|0|10|||7456|8|||1|531566|254462|4|3|45
501273088|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-28|2017-02-28|Followup|2013-11-28|2013-12-20|Complete|Done|4|4|2|1|1|1|2.17|||||||||1|3|3|4|2|3|2.67|||||||||4|4|4|4||||||3|1|3|3|2.5|||||||4|4|4|4|3|3|3|3.57||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|51||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|F|Black||48|28213|Bachelors Degree|Single|Finance: Accountant||8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501273365|31|0|2|503079327|31|0|2|500659156|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|531597||4|3|45
502248033|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-06|2013-07-25|Followup|2013-02-06|2013-02-06|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|2|2|3|2.83|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Moved|17.6||1|1|1|1|M|Black||13|No|Mother|28273|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||28|28277|Bachelors Degree|Single|Business: Marketing||0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502248464|31|0|1|502841432|1|0|1|500591252|2||-2||4|3|||-2||-2|34|2|||7496|10|||1|531679||4|3|45
502604900|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-15|2015-05-14|Followup|2013-11-15|2013-12-23|Declined|Done||||||||3|1|1|1|1|1|1.33|||||||||1|1|2|1|1|3|1.5||||||4|4|4|4|||||||4|4|3|3|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|2|3||||1|1||||4|4||Green||Volunteer: Lost contact with child/agency|41.9||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||30|28211|Bachelors Degree|Single|Finance: Accountant|28204|0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502605417|1|0|1|502582742|1|0|1|500577855|2||-2||4|1|||-2|500000294|-2|6854|8|||7464|9|||1|532031|356462|4|1|45
502240205|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-22|2014-06-11|Followup|2013-09-22|2013-12-07|Expired|Late||||||||4|2|4|3|3|3|3.17|||||||||2|3|3|2|2|3|2.5||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||4|2|3||||2|2|||||||Green|Amachi|Child/Family: Lost contact with volunteer/agency|32.6||3|3|2|2|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||48|28203|Bachelors Degree|Married|Business: Mgt, Admin|28202|1|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002334|502240634|31|0|2|502657850|31|0|2|500553471|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|532548|156483|4|0|45
502507408|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-13|2016-08-22|Followup|2013-10-13|2013-12-28|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|58.3||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Less than $10,000||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||71|28277|Bachelors Degree|Married|Retired||0|0||Relative|Big|General Community||Match Support|277|60|598|500000170|500017732|502507857|31|0|1|502673562|31|0|1|500559678|2||-2||4|2|500005291||-2||-2|34|2|||0|11|||1|532549||4|0|45
500186192|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2014-10-13|Followup|2013-11-18|2013-11-16|Complete|Done|2|4|4|4|3|1|3|||||||||4|4|4|4|2|4|3.67|||||||||4|3|3|3.33||||||3|5|5|5|4.5|||||||4|3|3|4|4|4|4|3.71||||||||||3|4|1|2.67||||||2|1|1.5|||||1|1||||4|4||||Green||Child: Graduated|46.8||2|2|1|1|F|Black||20||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|Black||33|28208||Single|Service: Restaurant||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187762|31|0|2|502323059|31|0|2|500490136|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|532696||4|3|45
503163476|BBBS of Greater Charlotte|Main Office|C|Active|2012-11-30|NaT|Followup|2013-11-30|2014-01-14|Complete|Done|3|1|3|2|2|3|2.33|3|1|1|1|1|3|1.67|39.52|3|4|4|2|3|4|3.33|2|3|4|2|3|3|2.83|17.67|4|4|4|4|3|4|4|3.67|8.99|5|5|5|5|5|4|5|5|5|4.75|5.26|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|4|4|-8.25|2|2|2|1|2|1.5|33.33|2|2|2|2|0|4|4|4|4|0|Green|||51.5||1|1|1|1|M|Black||13|No|Mother|28269|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|Black||32|28217|Masters Degree|Single|Consultant||0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503165154|31|0|1|503119713|31|0|1|500663695|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|533054|530536|4|3|45
502359051|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-28|2017-02-28|Followup|2013-10-28|2013-11-18|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|3|4|3|4|4|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|76.1||1|1|1|1|F|Black||14|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||35|28213|Masters Degree|Married|Business: Clerical||3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502359489|31|0|2|502242295|31|0|2|500483954|2||500004772||4|3|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|10|||131|1|||1|533061||4|3|45
503063881|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-30|2015-01-14|Followup|2013-11-30|2014-01-14|Complete|Done|4|4|4|1|4|4|3.5|4|4|4|1|4|4|3.5|0|4|4|4|4|4|4|4|4|4|4|1|4|4|3.5|14.29|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|5|5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|4|4|4|-12.5|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Moved|25.5||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||34|28202|Associate Degree|Single|Medical: Healthcare Worker||6|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503065564|31|0|2|503125383|1|0|2|500656877|2||-2||4|2|||-2||-2|0|10|||46|2|||1|533107|518880|4|3|45
501234606|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-16|NaT|Followup|2013-09-16|2013-09-30|Complete|Done|3|3|4|3|4|4|3.5|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||2|2|2|2||||||4|4|4|||||2|2||||4|4||||Green|||101.9||1|1|1|1|F|Black||16|No|Mother|28216|Grandparents|Unknown||No|TV|Media|General Community||Match Support|F|Black||42|28212|Bachelors Degree|Single|Unknown|28202|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501234882|31|0|2|501233675|31|0|2|500287478|2||-2||2|1|||-2||-2|56|1|||7464|9|||1|533338||4|3|45
502261100|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-25|NaT|Followup|2013-01-25|2013-01-22|Complete|Done|4|4|4|1|2|4|3.17|||||||||2|2|4|3|3|4|3|||||||||2|4|4|3.33||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||73.7||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|F|White||35|28209|Bachelors Degree|Single|Retail: Sales||6|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502261532|31|0|2|502284382|1|0|2|500512216|2||-2||2|1|||-2||-2|0|3|||7464|9|||1|533437||4|3|45
503268271|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-27|2015-08-19|Baseline|2012-12-03|2012-12-21|Complete|Done|3|4|4|1|4|4|3.33|||||||||2|4|3|4|4|4|3.5|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|31.7||1|1|1|1|F|Black||13|No|Mother|28226|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||40|28273|Some College|Married|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503270085|31|0|2|502993922|1|0|2|500669147|2||-2||4|3|||-2||-2|6854|8|||7496|10|3|3|1|533978|-1|4|3|44
503029036|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-07|2014-02-10|Followup|2013-08-07|2013-08-28|Complete|Done|4|3|4|1|1|3|2.67|||||||||4|1|1|4|4|1|2.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Moved|18.1||1|1|1|1|M|Black||13|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Enrollment|M|Asian||33|30097|Bachelors Degree|Single|Business|28255|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002334|503030631|31|0|1|503070963|4|0|1|500626277|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|535519||4|3|45
501342393|BBBS of Greater Charlotte|Main Office|C|Completed|2008-10-22|2014-06-06|Followup|2013-10-22|2014-01-03|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Lost interest|67.4||1|1|1|1|F|White||19|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Business: Sales||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501342672|1|0|2|501210017|1|0|2|500293459|2||-2||4|1|||-2||-2|0|10|||46|2|||1|536486||4|1|45
500713817|BBBS of Greater Charlotte|Main Office|C|Active|2009-10-30|NaT|Followup|2013-10-30|2013-11-26|Complete|Done|4|3|4|3|3|4|3.5|||||||||3|2|4|3|3|4|3.17|||||||||4|4|4|4||||||5|5|3|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|||88.5||2|2|1|1|M|Black||16||Mother|28216|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28078|||Medical: Pharmacist|28210|10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|500714084|31|0|1|501834795|1|0|1|500396466|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|536487||4|3|45
502252822|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-11|2014-02-24|Followup|2013-10-11|2013-12-02|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|40.5||3|3|1|1|F|Black||13|No|GrandMother|28227|Grandparents|Unknown||No||Self|General Community||Match Support|F|White||34|28270||Single|Personal Trainer/Coach||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|502253254|31|0|2|502282155|1|0|2|500472826|2||-2||4|1|||-2||-2|0|10|||46|2|||1|536610||4|1|45
501853851|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-10-20|Followup|2013-04-30|2013-05-14|Complete|Done|3|2|3|2|4|4|3|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||3|4|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child/Family: Moved|41.7||2|2|1|1|M|Black||13|Yes|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||55|28105|Masters Degree|Married|Law: Lawyer||25|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|501854219|31|0|1|502922901|1|0|1|500608304|2||-2||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|537626||4|3|45
502083438|BBBS of Greater Charlotte|Main Office|C|Active|2012-02-02|NaT|Followup|2013-02-02|2013-01-02|Complete|Early|4|4|4|3|4|4|3.83|||||||||3|1|3|3|3|3|2.67|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|3|3|3.71||||||||||3|4|3|3.33||||||4|3|3.5|||||2|2||||4|4||||Green|Cabarrus County||61.4||1|1|1|1|F|Black||13|No|Mother|28083|One Parent: Female|Unknown||Yes||Self|General Community|Cabarrus County|Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502083853|31|0|2|502657267|31|0|2|500595491|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|10|||7496|10|||1|537634||4|3|45
502983808|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-15|2016-02-10|Baseline|2012-12-11|2012-12-15|Complete|Done|1|1|2|1|1|3|1.5|||||||||1|4|4|1|1|3|2.33|||||||||4|4|4|4||||||1|5|3|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|1|1|1.67||||||3|4|3.5|||||1|1||||4|4||||Yellow|Amachi|Volunteer: Time constraint|37.8||1|1|1|1|M|Black||15|Yes|Mother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||27|28203|Bachelors Degree|Single|Business||0|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502985262|31|0|1|503140432|1|0|1|500668771|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|538016|-1|4|3|44
502255210|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-27|NaT|Followup|2013-09-27|2013-10-03|Complete|Done|4|3|4|3|1|3|3|||||||||2|4|3|4|1|4|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||77.6||1|1|1|1|M|Black||14|No|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||29|28210|Bachelors Degree|Married|Business: Mgt, Admin|97224|6|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|500910307|31|0|1|502255794|1|0|1|500470233|2||-2||2|1|||-2|500000294|-2|0|10|||7496|10|||1|538393||4|3|45
500829028|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-30|NaT|Followup|2013-11-30|2013-12-02|Complete|Done|4|4|4|2|4|4|3.67|||||||||2|4|4|3|2|3|3|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|2|4|4|3|4|3|3.43||||||||||3|4|2|3||||||4|4|4|||||2|2||||4|4||||Green|||75.5||3|3|2|2|F|Black||17|No|Mother|28209|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||39|28210|Masters Degree|Single|Education|28212|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502254499|31|0|2|501978180|1|0|2|500498594|2||-2||2|1|||-2|500000294, 500004640|-2|0|10|||7464|9|||1|538585||4|3|45
502308197|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-03|2016-05-09|Followup|2013-12-03|2013-12-30|Complete|Done|4|4|4|4|4|4|4|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||5|3|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|65.2||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Enrollment|F|White||35|28210|Bachelors Degree|Living w/ Significant Other|Business: Sales|18034|2|7|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big AND Amachi|Match Support|277|60|598|500000170|500021785|502308629|31|0|2|502325667|1|0|2|500493122|2||500003586||4|1||500000294|-2|500000294, 500004901|-2|0|10|||7496|10|||1|538610||4|3|45
501060196|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-26|2015-08-03|Followup|2013-11-26|2014-02-10|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|92.2||1|1|1|1|M|Black||19|No|Mother|28205|One Parent: Female|$15,000 to $19,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28226|Masters Degree|Single|Finance: Accountant||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501060469|31|0|1|501036081|1|0|1|500223215|2||-2||4|1|||-2||-2|34|2|||46|2|||1|538697||4|0|45
502702145|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-21|2016-05-24|Followup|2013-12-21|2013-12-19|Complete|Done|4|3|4|3|4|4|3.67|3|3|4|3|4|4|3.5|4.86|4|4|4|1|4|4|3.5|3|4|4|4|4|4|3.83|-8.62|4|4|4|4|3|3|3|3|33.33|5|5|5|5|5|5|4|2|4|3.75|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|2|3|2.67|49.81|4|4|4|3|2|2.5|60|2|2|2|2|0|4|4|4|4|0|Red||Child: Graduated|53.1||1|1|2|2|F|Black||17|No|Mother|28083|One Parent: Female|$60,000 to $74,999||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020753|502702991|31|0|2|502204211|31|0|2|500582836|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|538711|375724|4|3|45
502753870|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2014-10-30|Followup|2013-11-30|2013-12-11|Complete|Done|4|4|4|3|3|4|3.67|3|3|3|2|3|3|2.83|29.68|4|4|4|4|4|4|4|4|1|2|3|3|3|2.67|49.81|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3||2|2|||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|2|3|2.67|49.81|3|4|3.5|3|4|3.5|0|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Time constraint|35||2|2|1|1|F|Hispanic||16|No|Mother|28262|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|F|White||31|28210|Masters Degree|Single|Medical: Doctor, Provider||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502751081|3|0|2|502785389|1|0|2|500574313|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|538724|363493|4|3|45
500186742|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-08|2016-06-30|Followup|2013-12-08|2013-12-13|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|Amachi|Child: Graduated|66.7||4|4|1|1|M|Black||19|Yes|Mother|28227|One Parent: Female|Unknown|Y|No||School|General Community|Amachi|Match Support|M|Black||52|28227|Masters Degree|Married|Education: Teacher|28227|2|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|502397541|31|0|1|500501282|2||500003586||4|1|500000294|500000294|-2|500000294, 500004640|-2|0|4|||12183|14|635|1|1|538738||4|3|45
502758832|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-17|2014-10-23|Followup|2013-12-17|2013-12-16|Complete|Done|4|2|4|2|4|4|3.33|4|4|4|4|3|3|3.67|-9.26|3|4|3|3|4|4|3.5|1|3|3|2|1|3|2.17|61.29|4|4|4|4|4|4|4|4|0|5|2|2|4|3.25|4|5|4|5|4.5|-27.78|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|3|3.67|3|4|3|3.33|10.21|4|4|4|3|4|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Green||Child: Family structure changed|34.2||1|1|1|1|F|White||14|No|Mother|28027|One Parent: Female|$50,000 to $59,999||No||Relative|General Community||Match Support|F|White||33|28027|Masters Degree|Single|Education: Teacher|28027|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502759744|1|0|2|502666962|1|0|2|500586238|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|538749|381135|4|3|45
502183420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-28|2015-01-15|Followup|2013-09-28|2013-12-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Time constraint|51.6||2|2|1|1|M|Multi-race (Black & White)||14|Yes|GrandMother|28215|Grandparents|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||58|28226|Masters Degree|Married|Tech: Sales, Mktg|28202|6|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502183840|36|0|1|502264770|1|0|1|500473793|2||500003586||4|2|500000294|500000294|-2||-2|7016|11|||7464|9|||1|539078||4|0|45
502866079|BBBS of Greater Charlotte|Main Office|C|Active|2013-03-26|NaT|Baseline|2012-12-13|2013-03-26|Complete|Done|4|1|1|1|1|1|1.5|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||5|5|4|3|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||1|3|1|1.67||||||4|1|2.5|||||2|2||||4|4||||Green|||47.7||1|1|1|1|M|White||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||32|28210|Bachelors Degree|Single|Business: Sales||4|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|502867478|1|0|1|503378886|1|0|1|500686789|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|539346|-1|4|3|44
502247579|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-02|2016-05-10|Followup|2013-12-02|2014-01-16|Declined|Done||||||||4|3|3|2|3|4|3.17|||||||||2|3|2|2|2|3|2.33||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|53.3||2|2|1|1|F|Black||15|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||47|28226|Bachelors Degree|Single|Education: Teacher||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500017732|502248010|31|0|2|502681447|31|0|2|500575685|2||500003586||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|10|||2238|7|||1|539835|194970|4|1|45
502760967|BBBS of Greater Charlotte|Main Office|C|Active|2011-12-08|NaT|Followup|2013-12-08|2014-02-12|Declined|Late||||||||1|2|4|1|3|3|2.33|||||||||4|4|4|4|3|4|3.83||||||4|2|2|2.67|||||||5|5|5|5|5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|3|3.5||||2|2||||4|4||Green|||63.2||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|$25,000 to $29,999|Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||29|28120|Bachelors Degree|Single|Govt: Clerical||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502761879|31|0|2|502666332|31|0|2|500579826|2||-2||2|1||500005291|-2||-2|2203|12|||7464|9|||1|539855|351583|4|1|45
502776341|BBBS of Greater Charlotte|Main Office|C|Active|2012-12-14|NaT|Followup|2013-12-14|2013-12-18|Complete|Done|4|4|4|4|3|3|3.67|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||51||1|2|1|2|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|White||31|28202|Bachelors Degree|Single|Retail: Mgt|28273|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502777520|31|0|2|502631040|1|0|2|500652764|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|539864||4|3|45
502180724|BBBS of Greater Charlotte|Main Office|C|Active|2010-12-30|NaT|Followup|2013-12-30|2013-12-23|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|3|2|2|4|2.83|||||||||4|4|4|4||||||2|2|2|2|2|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||74.5|Y|2|2|2|2|M|Black||15|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502181148|31|0|1|502391505|31|0|2|500505039|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7438|1|||1|539985||4|3|45
502983808|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-15|2016-02-10|Followup|2013-12-15|2014-03-01|Expired|Late||||||||1|1|2|1|1|3|1.5|||||||||1|4|4|1|1|3|2.33||||||4|4|4|4|||||||1|5|3|5|3.5||||||||||4|4|4|4|4|4|4|4||||||3|1|1|1.67|||||3|4|3.5||||1|1||||4|4||Yellow|Amachi|Volunteer: Time constraint|37.8||1|1|1|1|M|Black||15|Yes|Mother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||27|28203|Bachelors Degree|Single|Business||0|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502985262|31|0|1|503140432|1|0|1|500668771|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|540234|538016|4|0|45
502184849|BBBS of Greater Charlotte|Main Office|C|Active|2012-12-18|NaT|Followup|2013-12-18|2013-12-23|Complete|Done|3|4|4|3|3|4|3.5|||||||||3|4|4|3|4|3|3.5|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2|||||||||Green|||50.9||2|2|1|1|M|Multi-race (Hispanic & White)||13|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||28|28210|Bachelors Degree|Single|Business: Marketing|28224|1|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|502185278|35|0|1|503145815|1|0|1|500658541|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|541479||4|3|45
502551048|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-19|2015-01-15|Followup|2013-10-19|2013-10-29|Complete|Done|4|4|4|3|4|4|3.83|||||||||1|2|3|1|1|2|1.67|||||||||4|4|4|4||||||2|3|5|1|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Yellow||Volunteer: Moved|38.9||1|1|2|2|F|Hispanic||13|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Enrollment|F|Black||52|30080|Bachelors Degree|Single|Consultant|2451|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502551498|3|0|2|501472128|31|0|2|500554178|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|541738||4|3|45
501129781|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-15|2015-01-15|Followup|2013-11-15|2013-12-02|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|1|4|3.17|||||||||4|4|4|4||||||5|4|3|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Family structure changed|50||1|2|4|6|F|Black||17||Mother|28217|Two Parent|Unknown||No||School|General Community||Match Support|F|Black||48|28273|Bachelors Degree|Married|Business: Mgt, Admin|28273|4|0|Recruitment Event|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500018987|501130055|31|0|2|500189245|31|0|2|500494855|2||-2||4|1|||-2||-2|0|4|||7459|10|||1|541740||4|3|45
502589869|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2015-10-29|Followup|2013-11-30|2014-01-21|Declined|Late||||||||4|2|2|3|1|1|2.17|||||||||2|4|4|4|4|4|3.67||||||4|4|4|4|||||||4|5|4|5|4.5||||||||||4|3|4|4|4|4|3|3.71||||||4|3|4|3.67|||||2|3|2.5||||2|2||||4|4||Green|Project Big|Child/Family: Lost contact with volunteer/agency|46.9||2|2|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28205|Bachelors Degree|Married|Business|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502590381|31|0|2|502701252|1|0|2|500582617|2||500004641||4|1|500004640|500004640, 500005291|-2|500000294|-2|0|4|459|3|7496|10|||1|541741|290937|4|1|45
500186190|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-13|2014-08-20|Followup|2013-10-13|2013-10-18|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|4||3||||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|118.2||1|1|2|2|F|Black||20||Mother|28213|Other/Unknown|Unknown||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500187761|31|0|2|500189140|31|0|2|500037140|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|543014||4|3|45
500733695|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-26|2015-03-03|Followup|2013-12-26|2014-01-29|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|3|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.2||1|1|1|1|F|Black||19|Yes|GrandMother|28217|Grandparents|Less than $10,000|Y|No|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||34|28210|Bachelors Degree|Married|Finance: Accountant|28202|0|2|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500733962|31|0|2|500307108|1|0|2|500150172|2||500003586||4|3|500000294|500000294|-2||-2|7294|13|||2238|7|||1|543349||4|3|45
502173821|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-18|2014-08-29|Followup|2013-11-18|2014-01-02|Complete|Done|4|3|3|2|4|4|3.33|4|1|1|1|4|4|2.5|33.2|4|4|4|4|3|4|3.83|3|4|4|3|3|4|3.5|9.43|4|4|4|4|4|4|4|4|0|5|5|4|4|4.5|5|5|4|4|4.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|2|2|2|50|2|2|1|1|100|4|4||||Red|Amachi|Volunteer: Time constraint|45.3||2|2|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||32|28262|Masters Degree|Single|Finance: Banking|28262|3|11|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502174240|31|0|2|502264706|1|0|2|500491573|2||500003586||4|3|500000294|500000294|-2|500000294, 500004640|-2|7016|11|||7464|9|||1|543430|148526|4|3|45
501853848|BBBS of Greater Charlotte|Main Office|C|Completed|2009-11-30|2014-08-29|Followup|2013-11-30|2014-01-14|Complete|Done|4|3|4|2|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|56.9||1|1|1|1|M|Black||15|Yes|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|M|Black||33|28273|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501854219|31|0|1|501839466|31|0|1|500405366|2||-2||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|543431||4|3|45
502310004|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-26|2014-05-01|Followup|2013-10-26|2013-11-12|Complete|Done|4|2|4|3|3|3|3.17|4|4|4|4|3|3|3.67|-13.62|3|3|3|4|2|4|3.17|2|3|4|4|3|4|3.33|-4.8|4|4|4|4|4|4|4|4|0|4|3|4|2|3.25|3|3|3|3|3|8.33|4|4|4|3|1|3|3|3.14|4|4|4|4|4|4|3|3.86|-18.65|4|4|3|3.67|4|4|3|3.67|0|3|4|3.5|3|3|3|16.67|2|2|2|2|0|4|4||||Yellow|Amachi, Project Big, Project Big AND Amachi|Volunteer: Moved|42.2||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||No||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Enrollment|F|White||37|28078||Single|Business||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502310436|31|0|2|502331000|1|0|2|500483762|2||500003586||4|2|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7496|10|||1|543624|194875|4|3|45
502371558|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-31|NaT|Followup|2013-10-31|2013-11-25|Complete|Done|3|4|4|4|4|4|3.83|3|2|3|3|3|3|2.83|35.34|3|4|4|3|3|3|3.33|3|4|4|3|2|4|3.33|0|4|2|3|3|4|4|4|4|-25|5|4|3|3|3.75|4|4|4|5|4.25|-11.76|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|3|3.67|4|4|3|3.67|0|4|4|4|4|2|3|33.33|2|2|1|1|100|4|4|4|4|0|Green|||64.5||1|1|2|2|M|Black||17|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020752|502371997|31|0|1|502528355|1|0|1|500568298|2||-2||2|1||500000294, 500005291|-2||-2|0|10|||132|8|||1|543625|355033|4|3|45
502619306|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-22|2014-12-17|Followup|2013-10-22|2013-11-11|Complete|Done|3|4|4|1|4|4|3.33|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|37.8||1|1|2|2|F|Hispanic||13|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|White||35|28205|Masters Degree|Married|Education: Teacher|28205|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|277|60|598|500000170|500017777|502619917|3|0|2|502716664|1|0|2|500565374|2||-2||4|1|||-2|500015184|-1|0|10|||7462|13|||1|543725||4|3|45
503268271|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-27|2015-08-19|Followup|2013-12-27|2014-02-09|Complete|Done|3|2|4|2|3|3|2.83|3|4|4|1|4|4|3.33|-15.02|3|4|4|4|4|4|3.83|2|4|3|4|4|4|3.5|9.43|4|4|4|4|4|4|4|4|0|4|4|4|4|4|5|4|5|4|4.5|-11.11|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|2|3|33.33|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|31.7||1|1|1|1|F|Black||13|No|Mother|28226|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||40|28273|Some College|Married|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503270085|31|0|2|502993922|1|0|2|500669147|2||-2||4|3|||-2||-2|6854|8|||7496|10|3|3|1|543813|533978|4|3|45
502708670|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-23|2014-02-06|Followup|2013-12-23|2013-12-23|Complete|Done|3|1|2|1|2|2|1.83|||||||||2|1|3|2|1|2|1.83|||||||||4|4|4|4||||||2|4|3|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||1|3|1|1.67||||||4|2|3|||||1|1||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|25.5||1|1|1|1|F|Black||18|No|Mother|28209|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||28|28215|Bachelors Degree|Single|Customer Service|28078|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500015820|502709557|31|0|2|502756331|1|0|2|500584031|2||-2||4|3|||-2||-2|0|4|||7462|13|||1|544663|377810|4|3|45
501553422|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2014-07-17|Followup|2013-08-03|2013-08-03|Complete|Done|4|1|1|1|3|4|2.33|||||||||2|4|3|2|1|3|2.5|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|35.4||4|4|1|1|F|Black||13|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Enrollment|F|Black||31|28212|Masters Degree|Single|Human Services|28211|0|1|Sigma Gamma Rho|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500013781|501536657|31|0|2|502646582|31|0|2|500548206|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||8700|14|||1|544876||4|3|45
502083429|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-11|2016-08-19|Followup|2014-02-11|2014-03-05|Complete|Done|3|4|4|3|2|4|3.33|4|2|4|3|2|4|3.17|5.05|3|4|3|2|3|4|3.17|4|4|4|1|4|4|3.5|-9.43|4|4|4|4|4|3|3|3.33|20.12|2|5|4|5|4|3|5|4|4|4|0|4|4|4|4|4|4|3|3.86|4|2|4|4|4|4|3|3.57|8.12|3|4|4|3.67|4|4|4|4|-8.25|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Moved|54.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Cabarrus County|Match Support|F|Black||29|28027|Bachelors Degree|Single|Education: Teacher||1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|502083853|31|0|2|502653045|31|0|2|500590992|2||-2||4|3||500016374|-2|500016374|-2|7016|11|||7464|9|||1|544940|220254|4|3|45
502083438|BBBS of Greater Charlotte|Main Office|C|Active|2012-02-02|NaT|Followup|2014-02-02|2014-03-05|Complete|Done|2|1|4|4|1|2|2.33|||||||||1|2|3|1|4|4|2.5|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|Cabarrus County||61.4||1|1|1|1|F|Black||13|No|Mother|28083|One Parent: Female|Unknown||Yes||Self|General Community|Cabarrus County|Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502083853|31|0|2|502657267|31|0|2|500595491|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|10|||7496|10|||1|545066||4|3|45
502700500|BBBS of Greater Charlotte|Main Office|C|Active|2012-01-13|NaT|Followup|2014-01-13|2014-03-30|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||62.1||1|1|1|1|M|Black||13|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|White||30|28202|Bachelors Degree|Single|Business: Sales|28212|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502701345|31|0|1|502824634|1|0|1|500589524|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|545996||4|0|45
502435258|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-12|2014-10-30|Followup|2014-01-12|2014-03-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|33.6||2|2|1|1|F|Black||13|No|Relative: Other|28081|Other Relative|Unknown|Y|Yes||Self|General Community||Enrollment|F|Black||31|28025|Bachelors Degree|Single|Child/Day Care Worker|28027|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|502435701|31|0|2|502670193|31|0|2|500589905|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|546303||4|1|45
502882034|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-13|NaT|Followup|2013-06-13|2013-06-10|Complete|Done|4|2|1|4|1|4|2.67|||||||||1|4|4|2|1|4|2.67|||||||||4|4|4|4||||||5|3|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||57.1||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||27|28208|Bachelors Degree|Single|Business: Mgt, Admin|28213|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501390617|31|0|2|502983700|31|0|2|500615277|2||-2||2|1||500000294|-2||-2|0|10|||7464|9|||1|546619||4|3|45
500546821|BBBS of Greater Charlotte|Main Office|C|Completed|2007-02-21|2015-09-15|Followup|2014-02-21|2014-02-21|Complete|Done|4|4|4|4|3|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|102.8||1|1|3|3|M|Black||20|No|Mother|28083|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||52|28025||Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500012459|500547073|31|0|1|500790181|31|0|1|500159910|2||-2||4|1|||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|546699||4|3|45
501389722|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-06|2014-04-24|Followup|2014-02-06|2014-02-06|Complete|Done|2|3|3|2|4|4|3|||||||||3|3|3|3|3|4|3.17|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child: Graduated|62.5||1|1|1|1|F|White||21|No|Mother|28027|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||56|28027||Divorced|Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500012459|501390003|1|0|2|500787778|1|0|2|500337267|2||-2||4|1|||-2||-2|0|10|||46|2|||1|546701||4|3|45
501247269|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-21|NaT|Followup|2014-02-21|2014-02-21|Complete|Done|4|1|4|1|4|4|3|||||||||1|3|3|2|4|3|2.67|||||||||3|3|3|3||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|2010-2012 OJJDP JJI, Cabarrus County||72.8||2|2|1|1|F|White||15|No|Father|28025|One Parent: Male|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|White||43|28027|Associate Degree|Married|Student: College||4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500341682|1|0|2|501914025|1|0|2|500515263|2||500016307||2|1|500005291, 500016374|500016374|-2|500016374|-2|0|10|||7496|10|||1|546708||4|3|45
501023408|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-05|NaT|Followup|2013-11-05|2013-11-12|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Green|||100.3||1|1|1|1|M|Hispanic|Other South American|17|No|Mother|28273|One Parent: Female|Less than $10,000||Yes||Self|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501023677|3|15|1|501356600|1|0|1|500296545|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|546720||4|3|45
501092957|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-09|2014-05-15|Followup|2013-11-09|2013-12-16|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|42.2||2|2|1|1|M|Black||17|No|Mother|28027|One Parent: Female|$30,000 to $34,999||No|Radio|Media|General Community||Match Support|M|White||44|28269||Married|Finance: Banking||5|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|501093231|31|0|1|502294662|1|0|1|500484597|2||-2||4|1|||-2||-2|55|1|||7459|10|||1|546722||4|1|45
502728289|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-04|2017-03-09|Followup|2013-11-04|2014-01-03|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|64.1||1|1|1|1|F|Hispanic||13|No|Mother|28278|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community||Match Support|F|White||32|28211||Married|Finance||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|502729186|3|0|2|502339145|1|0|2|500565493|2||-2||4|1|||-2|500000294|-2|0|3|||7496|10|||1|546773||4|1|45
501252806|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-25|NaT|Followup|2013-11-25|2014-01-08|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|3|4|3|3|4|3.17|||||||||4|4|4|4||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||99.6||1|1|1|1|M|Black||13|No|Mother|28078|One Parent: Female|Unknown||No||Relative|General Community||Match Support|M|Black||45|28262|Bachelors Degree|Married|Business: Mgt, Admin||0|6|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|501253082|31|0|1|501320197|31|0|1|500310204|2||-2||2|1|||-2||-2|0|3|||6247|12|||1|547010||4|3|45
503170936|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-23|2013-01-31|Baseline|2013-01-10|2013-01-23|Complete|Done|3|1|3|2|3|2|2.33|||||||||2|3|4|1|4|4|3|||||||||3|4|4|3.67||||||5|5|5|5|5|||||||3|4|4|4|4|4|3|3.71||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green||Child: Severity of challenges|0.3||1|1|2|2|M|White||14|No|Mother|28277|Grandparents|Less than $10,000||Yes||Therapist/Counselor|General Community||Match Support|M|Asian|Indian|27|28277|Bachelors Degree|Single|Business|28277|0|2||Relative|Big|General Community||Enrollment|277|60|598|500000170|500004169|503172623|1|0|1|503258884|4|18|1|500674088|2||-2||4|1|||-2||-2|0|5|||0|11|||1|547194|-1|4|3|44
501353940|BBBS of Greater Charlotte|Main Office|C|Active|2011-11-30|NaT|Followup|2013-11-30|2014-01-02|Complete|Done|2|2|4|2|4|4|3|||||||||2|3|4|4|2|4|3.17|||||||||4|4|3|3.67||||||4|4|4|2|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|Amachi||63.5||3|3|1|1|M|Black||16|No|Relative: Other|28205|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||33|28226|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|10|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500020752|501354219|31|0|1|502710990|1|0|1|500574615|2||500003586||2|1|500000294|500000294, 500005291|-2||-2|34|2|||17161|11|||1|547265||4|3|45
502699353|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-31|2014-01-30|Followup|2013-10-31|2014-01-15|Expired|Late|3|2|2|1|2|||3|3|4|2|4|4|3.33||3|4|4|3|3|4|3.5|3|3|3|4|4|3|3.33|5.11|4|4|4|4|3|3|3|3|33.33|5|4|2|4|3.75|3|3|3|3|3|25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|3|3|3|3|22.33|2|2|2|3|3|3|-33.33|2|2|1|1|100|4|4|4|4|0|Yellow|Project Big|Volunteer: Moved|27||2|2|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown||No||School|General Community|PERL 2014-2016, Project Big|Match Support|F|White||29|28204|Bachelors Degree|Single|Business|28255|0|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502700198|31|0|2|502530062|1|0|2|500568290|2||-2||4|2|500004640|500004640, 500014681|-2|500000294|-2|0|4|||7464|9|||1|547937|355021|4|0|45
502469903|BBBS of Greater Charlotte|Main Office|C|Active|2012-02-22|NaT|Followup|2014-02-22|2014-02-24|Complete|Done|4|3|4|4|4|4|3.83|3|4|4|3|3|4|3.5|9.43|3|4|4|3|4|4|3.67|3|4|3|3|3|3|3.17|15.77|4|4|4|4|3|4|4|3.67|8.99|4|4|4|4|4|4|4|3|3|3.5|14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|2|1|1.5|100|2|2|1|1|100|4|4|4|4|0|Green|||60.7||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$15,000 to $19,999|Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||34|28269|Bachelors Degree|Single|Business: Human Resources|28025|2|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500020910|502470350|31|0|1|502868874|31|0|1|500594396|2||-2||2|1|||-2||-2|0|5|||4748|14|1360|3|1|548165|395896|4|3|45
501314104|BBBS of Greater Charlotte|Main Office|C|Active|2008-12-04|NaT|Followup|2013-12-04|2014-02-18|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|||99.4||1|1|1|1|M|Black||13|No|Mother|28217|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||39|28134|Bachelors Degree|Single|Business: Mgt, Admin||6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501314382|31|0|1|501170940|1|0|1|500315948|2||-2||2|2|||-2||-2|0|10|||7464|9|||1|548543||4|0|45
502255150|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-14|NaT|Followup|2014-02-14|2014-02-11|Complete|Done|4|1|1|1|4|4|2.5|1|2|1|1|1|4|1.67|49.7|1|3|4|1|1|4|2.33|1|4|3|1|1|3|2.17|7.37|4|4|4|4|4|4|4|4|0|1|3|1|1|1.5|2|3|3|2|2.5|-40|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|1|1|1|1|4|4|3|3.67|-72.75|1|1|1|1|1|1|0|2|2|2|2|0|4|4||||Green|Amachi||73||1|1|1|1|F|Black||17|Yes|Relative: Other|28227|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||34|28212|Masters Degree|Single|Education: Teacher|28216|6|3|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020752|502255582|31|0|2|502392989|1|0|2|500512287|2||500003586||2|1|500000294|500000294|-2|500000294, 500004640|-2|0|5|||7464|9|||1|548657|235505|4|3|45
501863951|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-18|2015-05-29|Followup|2013-12-18|2014-01-31|Complete|Done|3|4|3|2|4|4|3.33|||||||||3|4|4|4|3|4|3.67|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child: Lost interest|65.3||1|1|2|2|F|Black||14|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28078|Bachelors Degree|Single|Business: Human Resources|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501864324|31|0|2|501601161|31|0|2|500421259|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|549067||4|3|45
500938154|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-12|NaT|Followup|2014-01-12|2014-02-13|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||98.1||2|2|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||32|28208|Associate Degree|Single|Service: Restaurant|28211|4|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500938424|31|0|1|501446421|1|0|1|500323753|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|549612||4|3|45
501114434|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-23|2014-06-12|Followup|2013-12-23|2014-02-10|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|65.6||1|1|1|1|M|Black||20|No|Uncle|28206|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||33|28207|Masters Degree|Single|Finance: Accountant|28244|0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501114708|31|0|1|501315131|1|0|1|500324423|2||-2||4|3|500000294|500000294|-2||-2|0|10|||130|1|11|3|1|550779||4|1|45
502261100|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-25|NaT|Followup|2014-01-25|2014-01-24|Complete|Done|4|4|4|1|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||73.7||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|F|White||35|28209|Bachelors Degree|Single|Retail: Sales||6|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502261532|31|0|2|502284382|1|0|2|500512216|2||-2||2|1|||-2||-2|0|3|||7464|9|||1|550948||4|3|45
500796255|BBBS of Greater Charlotte|Main Office|C|Active|2010-01-20|NaT|Followup|2014-01-20|2014-02-21|Complete|Done|3|2|2|1|1|3|2|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4||3|3||||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||85.8||3|3|1|1|M|White||18|No|Mother|28031|One Parent: Male|$20,000 to $24,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||60|28269|||Medical: Admin|28207|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500796529|1|0|1|501846438|1|0|1|500424314|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|550962||4|3|45
502671406|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-14|2014-09-04|Followup|2014-02-14|2014-02-12|Complete|Done|1|4|4|4|4|4|3.5|3|4|4|3|3|3|3.33|5.11|2|3|3|2|2|3|2.5|3|3|2|3||3|||4|3|3|3.33|3|3|3|3|11|4|4|3|4|3.75|1|3|3|3|2.5|50|4|4|4|4|4|4|4|4|4|4|4|4|2|4|4|3.71|7.82|3|3|3|3|3|4|4|3.67|-18.26|2|1|1.5|3|1|2|-25|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Infraction of match rules/agency policies|30.7||1|1|1|1|F|Black||19|No|Mother|28210|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||34|28226|PHD|Single|Medical: Healthcare Worker|28207|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502672234|31|0|2|502885637|31|0|2|500597397|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|550978|400951|4|3|45
502634923|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-16|2015-02-20|Followup|2013-08-16|2013-09-26|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|42.2||1|1|1|1|F|Black||13|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community||Match Support|F|Black||42|28210|Masters Degree|Single|Business: Clerical|28036|3|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|502635617|31|0|2|501197016|31|0|2|500548227|2||-2||4|1|||-2||-2|0|3|||46|2|||1|551403||4|1|45
502934500|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-19|2013-10-31|Baseline|2013-01-24|2013-02-18|Complete|Done|2|2|4|2|2|3|2.5|||||||||4|4|3|4|4|4|3.83|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|3|4|2|3|4|3.43||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Red||Volunteer: Time constraint|8.3||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community||Match Support|M|Black||43|28216|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502935923|31|0|1|503123393|31|0|1|500676924|2||-2||4|3|||-2||-2|0|3|||7464|9|||1|552005|-1|4|3|44
503268324|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-26|2015-06-25|Baseline|2013-01-24|2013-01-26|Complete|Done|3|3|4|4|4|4|3.67|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|3|4|3|4|3|3.57||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Yellow||Child: Lost interest|28.9||1|1|1|1|M|Black||18|Yes|Mother|28226|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Asian||29|28277|Bachelors Degree|Single|Real Estate: Realtor|28277|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503270085|31|0|1|503253968|4|0|1|500676990|2||-2||4|2||500000294|-2||-2|6854|8|||7464|9|||1|552085|-1|4|3|44
502980965|BBBS of Greater Charlotte|Main Office|C|Active|2013-01-24|NaT|Followup|2014-01-24|2014-04-10|Expired|Late||||||||2|1|1||3|4||||||||||2|3|3|2|2|3|2.5||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|1|2||||2|2||||4|4||Green|||49.7||2|2|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||32|28210|High School Graduate|Single|Business: Sales|28277|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502982410|31|0|2|503091130|1|0|2|500676334|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|552155|447655|4|0|45
503052841|BBBS of Greater Charlotte|Main Office|C|Active|2013-01-24|NaT|Followup|2014-01-24|2014-01-21|Complete|Done|4|2|4|3|3|4|3.33|3|3|4|4|3|4|3.5|-4.86|3|3|4|3|4|4|3.5|4|4|4|3|4|4|3.83|-8.62|4|4|4|4|4|4|4|4|0|4|5|3|3|3.75|4|5|5|3|4.25|-11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green|||49.7||1|1|1|1|F|Hispanic||18|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||24|28104|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503027860|3|0|2|503122069|1|0|2|500660497|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|552190|511402|4|3|45
502839827|BBBS of Greater Charlotte|Main Office|C|Active|2013-01-31|NaT|Baseline|2013-01-24|2013-01-31|Complete|Done|3|4|4|3|3|4|3.5|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|4|4|2|3.71||||||||||4|3|4|3.67||||||2|2|2|||||1|1||||4|4||||Green|||49.4||1|1|1|1|M|Black||18|No|Mother|28215|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|Black||41|28105|Bachelors Degree|Single|Tech: Management|28202|0|6|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|502841119|31|0|1|503311280|31|0|1|500677083|2||-2||2|1|||-2||-2|0|10|||6247|12|||1|552197|-1|4|3|44
502839019|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-24|2016-01-28|Followup|2014-01-24|2014-03-04|Complete|Done|4|3|4|3|4|4|3.67|4|3|4|4|4|4|3.83|-4.18|3|3|4|4|3|3|3.33|3|4|3|2|4|4|3.33|0|4|4|4|4|4|4|4|4|0|4|5|4|4|4.25|5|4|4|5|4.5|-5.56|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|3|3.71|4.04|4|4|4|4|4|3|2|3|33.33|3|3|3|3|3|3|0|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Moved|36.1||1|1|1|1|M|Black||17|No|Mother|28210|One Parent: Female|$40,000 to $44,999|Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||32|28203|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502840311|31|0|1|502432390|31|0|1|500674451|2||-2||4|1|||-2||-2|6854|8|||7496|10|||1|552305|474477|4|3|45
502979759|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-12|2016-02-10|Baseline|2013-01-25|2013-03-12|Complete|Done|4|1|4|1|4|4|3|||||||||2|3|3|3|4|3|3|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||2|4|3|||||1|1||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|35||1|1|1|1|M|Black||16||Mother|28211|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||29|28211|Bachelors Degree||Construction|28208|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|502981210|31|0|1|503234517|1|0|1|500682418|2||-2||4|2|||-2||-2|0|10|||46|2|||1|552522|-1|4|3|44
503268324|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-26|2015-06-25|Followup|2014-01-26|2014-03-12|Complete|Done|3|3|3|2|4|3|3|3|3|4|4|4|4|3.67|-18.26|3|3|3|4|4|3|3.33|3|4|3|3|3|3|3.17|5.05|4|4|4|4|4|4|4|4|0|3|4|4|4|3.75|3|4|4|4|3.75|0|4|4|4|4|3|4|3|3.71|4|4|3|4|3|4|3|3.57|3.92|4|4|4|4|4|4|4|4|0|3|3|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Yellow||Child: Lost interest|28.9||1|1|1|1|M|Black||18|Yes|Mother|28226|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Asian||29|28277|Bachelors Degree|Single|Real Estate: Realtor|28277|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503270085|31|0|1|503253968|4|0|1|500676990|2||-2||4|2||500000294|-2||-2|6854|8|||7464|9|||1|552865|552085|4|3|45
501147999|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-26|2015-02-02|Followup|2014-01-26|2014-01-29|Complete|Done|4|1|4|4|4|4|3.5|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|24.2||2|2|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Unknown||No||School|General Community||Match Support|F|Black||35|28262|Bachelors Degree|Single|Insurance||6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|501148273|31|0|2|503112265|31|0|2|500665633|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|552868||4|3|45
502902269|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-26|2014-02-21|Followup|2014-01-26|2014-01-29|Complete|Done|1|2|4|2|3|3|2.5|4|3|4|1|3|4|3.17|-21.14|2|3|4|2|2|4|2.83|2|3|4|3|4|4|3.33|-15.02|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3|5|4|3|3.75|33.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|1|1|2|2|-50|4|4|4|4|0|Yellow||Child: Lost interest|12.8||1|1|3|3|M|Black||14|No|Mother|28215|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Enrollment|M|Black||31|28203|Juris Doctorate (JD)||Law: Lawyer|28203|1|0|Self|Self|Big|General Site|mentor2.0 2015|Match Support|277|60|598|500000170|500011349|502903679|31|0|1|501631588|31|0|1|500677452|2||-2||4|2|||-2|500015184|-1|0|10|||7464|9|||1|552870|417037|4|3|45
501529921|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2015-04-06|Followup|2014-01-23|2014-01-31|Complete|Done|3|2|2|2|3|2|2.33|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Time constraint|38.4||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||48|28031|Some College|Divorced|Medical|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501530213|31|0|2|502554719|1|0|2|500581908|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|553261||4|3|45
503010214|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-13|2013-06-19|Baseline|2013-01-28|2013-03-13|Complete|Done|4|2|4|4|3|4|3.5|||||||||2|3|3|2|3|3|2.67|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|1|2.5|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|3.2||1|1|1|1|M|Black||16|No|Mother|28226|One Parent: Female|$45,000 to $49,999||No||Self|General Community||Match Support|M|White||36|29708|Bachelors Degree|Married|Business: Sales|28216|10|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|503011744|31|0|1|503306996|1|0|1|500683223|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|553368|-1|4|3|44
503262762|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2014-01-06|Baseline|2013-01-29|2013-01-31|Complete|Done|4|4|4|4|4|4|4|||||||||3|3|3|3|4|3|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|2|3||||||2|4|3|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|11.2||1|1|1|1|F|Black||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||29|28203|Bachelors Degree|Single|Education: Teacher|28031|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503264570|31|0|2|503114924|1|0|2|500678106|2||-2||4|3|||-2||-2|34|2|||7464|9|||1|553946|-1|4|3|44
503238896|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2014-03-06|Baseline|2013-01-29|2013-01-31|Complete|Done|3|2|1|3|4|4|2.83|||||||||3|4|4|1|2|4|3|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|13.1||1|1|1|1|F|Black||16|No|Mother|28278|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|Black||27|28212|Bachelors Degree|Single|Finance: Banking||0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|503239061|31|0|2|503004093|31|0|2|500678152|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|553993|-1|4|3|44
503237270|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-08|2013-10-03|Baseline|2013-01-29|2013-02-08|Complete|Done|4|2|4|4|4|4|3.67|||||||||2|4|4|3|3|3|3.17|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|4|3.5|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|7.8||1|1|1|1|M|Black||17|No|Mother|28278|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||RTBM|M|Some Other Race||34|28212|Bachelors Degree|Single|Customer Service|28212|0|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|503239061|31|0|1|503022525|41|0|1|500678178|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|554016|-1|4|3|44
503015906|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-19|2013-05-23|Baseline|2013-01-30|2013-02-19|Complete|Done|4|1|2|2|3|3|2.5|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||5|2|3|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||2|4|3|||||1|1||||4|4||||Green||Child: Lost interest|3.1||1|1|2|2|M|White||17|No|Mother|28027|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|M|White||60|28027|Bachelors Degree|Separated|Insurance|28262|24|0|Local Radio|Media|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500015820|503017438|1|0|1|503041890|1|0|1|500678458|2||-2||4|1|||-2|500016374|-2|0|10|||7437|1|||1|554428|-1|4|3|44
500847570|BBBS of Greater Charlotte|Main Office|C|Active|2012-01-25|NaT|Followup|2014-01-25|2014-01-21|Complete|Done|3|2|3|2|3|4|2.83|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Yellow|Amachi||61.7||2|2|1|1|F|Black||16|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||52|28227|Bachelors Degree|Married|Insurance|28277|14|0|AA Task Force|Special Event|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188056|31|0|2|502542379|31|0|2|500592215|2||500003586||2|2|500000294|500000294|-2|500000294|-2|0|10|||11098|8|||1|554733||4|3|45
502555551|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-30|2016-08-18|Followup|2014-01-30|2014-01-31|Complete|Done|3|4|4|4|4|4|3.83|4|1|2|1|4|3|2.5|53.2|2|4|3|2|4|3|3|2|3|3|2|4|3|2.83|6.01|4|3|3|3.33|3|3|4|3.33|0|3|2|5|1|2.75|5|3|3|4|3.75|-26.67|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|3|3.67|3|4|3|3.33|10.21|4|4|4|4|4|4|0|2|2|2|2|0|4|4||||Green||Child/Family: Moved|42.6||2|2|1|1|M|Black||16|No|Aunt|28213|One Parent: Female|$40,000 to $44,999||Yes||School|General Community|Project Big|Match Support|M|White||33|28209|Associate Degree|Married|Business: Mgt, Admin||0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502556004|31|0|1|503207140|1|0|1|500674218|2||-2||4|1||500004640|-2||-2|0|4|||7464|9|||1|554735|318541|4|3|45
502097794|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-20|NaT|Followup|2014-01-20|2014-01-23|Complete|Done|3|3|3|2|3|3|2.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green|||73.8||1|1|1|1|M|Black||13|No|Mother|28269|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28031|Bachelors Degree|Single|Business: Engineer|28036|0|8|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502098218|31|0|1|502425119|1|0|1|500510881|2||-2||2|1|||-2|500000294, 500004640|-2|34|2|||46|2|||1|554834||4|3|45
502193174|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2015-07-30|Followup|2014-01-31|2014-01-29|Complete|Done|4|2|4|3|3|3|3.17|4|1|1|4|2|4|2.67|18.73|3|3|3|3|3|2|2.83|1|3|3|2|3|3|2.5|13.2|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|2|5|5|4|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|2|2|0|4|4||||Green||Volunteer: Moved|29.9||2|2|1|1|M|Black||16||Mother|28273|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|M|White||32|28273|Bachelors Degree|Single|Business: Mgt, Admin|28217|3|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|502193603|31|0|1|503100143|1|0|1|500677433|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|555022|168695|4|3|45
502254067|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2014-03-13|Followup|2014-01-31|2014-02-07|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|4|3.5|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|13.3||3|3|1|1|F|Black||14|No|Mother|28209|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|F|Black||39|28213|Bachelors Degree|Married|Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502254499|31|0|2|503047588|31|0|2|500677904|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|555196||4|3|45
503026286|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2017-02-26|Followup|2014-01-31|2014-01-29|Complete|Done|4|2|4|3|3|4|3.33|3|3|4|4|3|3|3.33|0|3|3|3|3|3|3|3|3|3|3|3|3|2|2.83|6.01|4|4|3|3.67|4|4|4|4|-8.25|4|3|2|3|3|5|2|3|4|3.5|-14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|48.9||1|1|1|1|M|Hispanic||17|No|Mother|28277|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Asian||30|28277|Bachelors Degree|Single|Finance||1|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503027860|3|0|1|503259120|4|0|1|500674960|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|555241|530932|4|3|45
502839827|BBBS of Greater Charlotte|Main Office|C|Active|2013-01-31|NaT|Followup|2014-01-31|2014-01-21|Complete|Done|3|2|3|2|3|4|2.83|3|4|4|3|3|4|3.5|-19.14|2|3|4|3|3|4|3.17|2|3|3|3|3|3|2.83|12.01|4|4|4|4|4|4|4|4|0|3|4|5|5|4.25|4|3|4|5|4|6.25|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|2|3.71|0|3|4|3|3.33|4|3|4|3.67|-9.26|2|3|2.5|2|2|2|25|2|2|1|1|100|4|4|4|4|0|Green|||49.4||1|1|1|1|M|Black||18|No|Mother|28215|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|Black||41|28105|Bachelors Degree|Single|Tech: Management|28202|0|6|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|502841119|31|0|1|503311280|31|0|1|500677083|2||-2||2|1|||-2||-2|0|10|||6247|12|||1|555427|552197|4|3|45
502980471|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-16|2013-07-16|Baseline|2013-01-31|2013-02-16|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|3|3|4|3|3|||||||||3|3|3|3||||||3|3|3|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|4.9||1|1|2|2|M|Black||18|No|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community|Project Big|Match Support|M|Asian|Indian|27|28277|Bachelors Degree|Single|Business|28277|0|2||Relative|Big|General Community||Enrollment|277|60|598|500000170|500008321|502981923|31|0|1|503258884|4|18|1|500678978|2||-2||4|3||500004640|-2||-2|34|2|||0|11|||1|555461|-1|4|3|44
503238896|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2014-03-06|Followup|2014-01-31|2014-02-13|Complete|Done|3|4|4|4|4|4|3.83|3|2|1|3|4|4|2.83|35.34|4|4|4|4|4|4|4|3|4|4|1|2|4|3|33.33|4|4|4|4|4|4|4|4|0|3|5|5|4|4.25|4|5|5|5|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|1|1|2|2|-50|4|4|4|4|0|Red||Volunteer: Time constraint|13.1||1|1|1|1|F|Black||16|No|Mother|28278|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|Black||27|28212|Bachelors Degree|Single|Finance: Banking||0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|503239061|31|0|2|503004093|31|0|2|500678152|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|555465|553993|4|3|45
501319029|BBBS of Greater Charlotte|Main Office|C|Completed|2013-01-31|2016-06-06|Followup|2014-01-31|2014-01-28|Complete|Done|1|1|2|1|1|1|1.17|||||||||4|3|4|4|1|4|3.33|||||||||4|4|4|4||||||3|5|5|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||1|2|1|1.33||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Moved|40.1||4|4|1|1|F|Black||13|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||28|28212|Bachelors Degree|Married|Child/Day Care Worker||0|3|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|503078205|1|0|2|500673752|2||-2||4|3||500014681|-2||-2|0|10|||7439|1|||1|555602||4|3|45
501536365|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-03|2014-07-17|Followup|2014-02-03|2014-03-12|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|1|4|4|3.57||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Time constraint|65.4||1|1|1|1|M|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Enrollment|M|Black||57|28105|Some College|Married|Retail: Sales|28105|10|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501536657|31|0|1|501443152|31|0|1|500336020|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|555785||4|3|45
501296349|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-01|2014-02-27|Followup|2013-12-01|2014-02-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|62.9||1|1|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||42|28214|Bachelors Degree|Single|Business: Mgt, Admin|28205|3|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501296627|31|0|2|501471640|31|0|2|500318555|2||||4|2|||-2|500000294|-2|0|4|||7464|9|||1|555887||4|0|45
501201377|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-31|2016-08-26|Followup|2014-01-31|2014-04-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|90.8||1|1|1|1|F|Hispanic||18|No|Mother|28212|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community||Match Support|F|Hispanic||65|28269|Masters Degree|Single|Medical: Admin|28262|8|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500017777|501201651|3|0|2|501497622|3|0|2|500331903|2||-2||4|3|||-2||-2|7016|11|||7446|3|||1|556272||4|0|45
501347056|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2015-10-12|Followup|2013-12-12|2014-02-26|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|82||1|1|1|1|M|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28226|Bachelors Degree|Married|Tech: Engineer|28202|2|8|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|501347335|31|0|1|501217000|1|0|1|500322327|2||-2||4|2|||-2||-2|34|2|||7446|3|||1|556345||4|0|45
502673798|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-30|2014-04-24|Followup|2014-01-30|2014-03-16|Declined|Done||||||||4|1|1|3|4|4|2.83|||||||||1|1|3|2|1|4|2||||||4|4|3|3.67|||||||5|5|3|3|4||||||||||4|4|4|4|1|4|4|3.57||||||4|3|4|3.67|||||2|1|1.5||||2|2||||4|4||Yellow||Volunteer: Time constraint|26.8||1|1|1|1|M|Black||17|No|Mother|28105|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|White||36|28173|Bachelors Degree|Separated|Business: Mgt, Admin|28110|15|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502674626|31|0|1|502860952|1|0|1|500590803|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|556488|389961|4|1|45
502236255|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-24|2014-11-30|Followup|2014-02-24|2014-04-03|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|4|3|2|2|4|2.83|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|45.2||1|1|1|1|M|Black||14|No|Father|28214|Two Parent|Unknown||Yes||Relative|General Community||Match Support|M|White||64|28207|Masters Degree|Married|Education: Teacher||0|0|Radio|Media|Big|General Site|mentor2.0 2015|Enrollment|277|60|598|500000170|500013781|502236686|31|0|1|502436546|1|0|1|500518376|2||-2||4|3|||-2|500015184|-1|0|3|||131|1|||1|556497||4|3|45
500843863|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-21|2016-06-17|Followup|2014-02-21|2014-03-23|Complete|Done|3|4|4|4|4|3|3.67|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||2|4|1|2.33||||||1|3|2|||||2|2||||4|4||||Green|Amachi|Volunteer: Changed workplace/school partnership|99.8||2|2|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|No|TV|Media|General Community|Amachi|Match Support|F|Black||32|28269|Bachelors Degree|Single|Business: Marketing|28273|0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500844129|31|0|2|501078655|31|0|2|500241388|2||500003586||4|1|500000294|500000294|-2|500000294|-2|56|1|||2238|7|||1|556789||4|3|45
502290605|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-09|2014-06-12|Followup|2013-05-09|2013-05-30|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red|Amachi|Volunteer: Moved|37.1||1|1|2|2|M|Black||13|Yes|Mother|28216|One Parent: Female|Unknown||Yes|Radio|Media|General Community|Amachi|Enrollment|M|Black||48|28269||Divorced|Tech: Engineer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502291037|31|0|1|500908500|31|0|1|500533937|2||-2||4|3|500000294|500000294|-2||-2|55|1|||7496|10|||1|557166||4|3|45
502244776|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-19|NaT|Followup|2014-01-19|2014-03-24|Declined|Late||||||||4|2|2|1|3|4|2.67|||||||||2|3|3|2|3|2|2.5||||||4|3|2|3|||||||2|3|3|4|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|4|3||||2|2||||4|4||Green|2010-2012 OJJDP JJI||73.9||1|1|2|2|F|Black||16|No|Mother|28216|Two Parent|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28209|Bachelors Degree|Single|Law|28273|5|0|Relative|Relative|Big|General Community|Amachi|Match Support|277|60|598|500000170|500021785|502245202|31|0|2|502143351|1|0|2|500511171|2||-2||2|1|500005291|500005291|-2|500000294|-2|0|4|||17161|11|||1|557615|233727|4|1|45
502308593|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-23|2015-05-28|Followup|2013-11-23|2014-02-07|Expired|Late||||||||4|2|3|1|3|4|2.83|||||||||3|3|4|4|3|3|3.33||||||3|2|3|2.67|||||||3|4|5|2|3.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|3|2.5||||1|1|||||||Red||Child/Family: Moved|54.1||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||40|28278|Bachelors Degree|Married|Tech: Computer/Programmer||3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502309025|31|0|1|502262702|31|0|1|500492994|2||-2||4|3|||-2||-2|0|10|||12183|14|1209|1|1|557682|206463|4|0|45
501390344|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-26|NaT|Followup|2014-02-26|2014-02-26|Complete|Done|4|3|3|3|4|4|3.5|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi||96.6||1|1|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Single|Tech: Computer/Programmer||0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|501390617|31|0|1|501380163|1|0|1|500342682|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|557877||4|3|45
502637766|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-12|2017-01-24|Followup|2013-07-12|2013-08-15|Complete|Done|3|3|3|2|2|2|2.5|||||||||2|3|2|1|2|3|2.17|||||||||4|4|4|4||||||2|3|4|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|54.4||1|1|1|1|M|Black||13|No|Mother|28262|One Parent: Female|$50,000 to $59,999||Yes||School|General Community||Match Support|M|Black||34|28269|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500021785|502638462|31|0|1|503016558|31|0|1|500619500|2||-2||4|1|||-2||-2|0|4|||7462|13|||1|558173||4|3|45
502335675|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-30|2016-10-31|Followup|2013-12-30|2014-02-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi, Project Big, Project Big AND Amachi|Child: Lost interest|70||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|Project Big AND Amachi|Match Support|M|White||27|28262||Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502336110|31|0|1|502305990|1|0|1|500495220|2||500004772||4|3|500000294, 500004640, 500004901|500004901|-2|500000294, 500004640|-2|0|4|||7496|10|||1|558644||4|1|45
502868923|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-27|2015-10-30|Followup|2014-01-27|2014-03-14|Complete|Late|4|4|4|2|4|4|3.67|||||||||2|4|4|3|4|3|3.33|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Volunteer: Moved|45.1||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Black||28|28262|Bachelors Degree|Single|Finance: Banking||0|0|AA Task Force|Special Event|Big|General Community||Match Support|277|60|598|500000170|500008321|502870324|31|0|2|502832013|31|0|2|500591320|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||11098|8|||1|558648||4|3|45
502580335|BBBS of Greater Charlotte|Main Office|C|Active|2011-11-30|NaT|Followup|2013-11-30|2013-12-17|Complete|Done|3|4|4|4|3|4|3.67|3|2|1|1|1|3|1.83|100.55|3|4|3|4|4|4|3.67|2|4|3|1|4|3|2.83|29.68|4|4|4|4|4|4|3|3.67|8.99|4|3|4|4|3.75|5|2|4|4|3.75|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|3|3.33|4|4|3|3.67|-9.26|2|3|2.5|3|2|2.5|0|2|2|2|2|0|4|4|4|4|0|Green|||63.5||1|1|1|1|F|Black||16||GrandMother|28269|Grandparents|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28269|Masters Degree|Single|Finance: Banking|28255|15|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502580838|31|0|2|502677590|31|0|2|500571804|2||-2||2|1||500005291|-2||-2|0|10|||7464|9|||1|558691|355336|4|3|45
502482642|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-11|2015-06-19|Followup|2014-02-11|2014-04-15|Declined|Late||||||||3|3|4|3|3|3|3.17|||||||||3|3|3|4|2|3|3||||||4|4|4|4|||||||3|4|4|4|3.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|2|2.5||||2|2||||4|4||Yellow||Child/Family: Moved|28.2||2|2|1|1|F|Black||16|No|Mother|28052|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||29|28277|Bachelors Degree|Single|Business|28217|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502391834|31|0|2|503118336|1|0|2|500679560|2||-2||4|2||500004640, 500005291|-2||-2|0|10|||7464|9|||1|558775|307140|4|1|45
501621811|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-16|2017-03-09|Followup|2014-03-16|2014-05-20|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Project Big|Child/Family: Lost contact with volunteer/agency|95.8||1|1|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||36|28269||Married|Self-Employed, Entrepreneur|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501622131|31|0|2|501621016|31|0|2|500344465|2||-2||4|2|500004640||-2||-2|0|10|||7464|9|||1|559357||4|1|45
502197486|BBBS of Greater Charlotte|Main Office|C|Active|2012-02-22|NaT|Followup|2014-02-22|2014-02-26|Complete|Done|4|1|3|2|4|4|3|||||||||4|4|3|3|2|4|3.33|||||||||4|4|4|4||||||4|3|2|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green|||60.7||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||30|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502197915|31|0|1|502870668|1|0|1|500597982|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|559362||4|3|45
501811395|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-10|NaT|Followup|2014-03-10|2014-03-10|Complete|Done|3|1|2|1|2|3|2|||||||||2|4|3|2|4|4|3.17|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||2|3|4|3||||||3|4|3.5|||||2|2||||4|4||||Green|Cabarrus County||84.2||1|1|1|1|F|Black||15|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||60|28213||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501811730|31|0|2|500876892|31|0|2|500436702|2||500016307||2|1|500016374|500016374|-2|500016374|-2|6854|8|||2238|7|||1|559515||4|3|45
502053779|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-13|2014-08-29|Followup|2014-02-13|2014-03-29|Complete|Done|4|3|3|3|4|4|3.5|3|3|3|2|3|4|3|16.67|3|3|3|3|4|4|3.33|2|3|3|1|2|3|2.33|42.92|4|4|4|4|4|4|4|4|0|4|4|2|4|3.5|3|3|2|4|3|16.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|3|3.67|8.99|3|2|2.5|3|3|3|-16.67|2|2|2|2|0|4|4||||Red||Volunteer: Feels incompatible with child/family|18.5||2|2|2|2|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community||Match Support|F|Black||49|28269|Bachelors Degree|Divorced|Finance|28282|0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500008321|502054203|31|0|2|500189241|31|0|2|500677878|2||-2||4|3|||-2||-2|7295|11|||7496|10|||1|559835|140517|4|3|45
502551047|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-21|2013-09-18|Baseline|2013-02-13|2013-02-21|Complete|Done|4|3|4|2|3|4|3.33|||||||||1|4|3|2|2|3|2.5|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|3|4|4|3|4|4|3.71||||||||||3|4|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|6.9||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Enrollment|M|White||28|28262|Some College|Single|Military|27260|6|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502551498|31|0|1|503347969|1|0|1|500681888|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|560049|-1|4|3|44
501227649|BBBS of Greater Charlotte|Main Office|C|Active|2013-02-14|NaT|Followup|2014-02-14|2014-02-13|Complete|Done|3|4|4|3|4|4|3.67|||||||||4|4|4|4|3|4|3.83|||||||||4|3|3|3.33||||||5|2|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|4|3|||||2|2||||4|4||||Green|Cabarrus County||49||2|2|1|1|M|White||16|Yes|GrandMother|28083|Grandparents|Unknown|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||51|28117|Masters Degree|Divorced|Consultant|28117|12|11|Local Print|Media|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501227925|1|0|1|503316978|1|0|1|500677437|2||500016307||2|1|500016374|500000294, 500016374|-2|500016374|-2|0|10|||7439|1|||1|560429||4|3|45
502663937|BBBS of Greater Charlotte|Main Office|C|Active|2013-02-27|NaT|Baseline|2013-02-15|2013-02-27|Complete|Done|2|4|4|4|3|4|3.5|||||||||3|2|4|2|3|4|3|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||48.6||1|1|1|1|M|Black||15|No|Mother|28212|Two Parent|$35,000 to $39,999||No||Relative|General Community||Match Support|M|White||30|28105|Bachelors Degree|Single|Business: Sales|17001|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502664764|31|0|1|503296990|1|0|1|500684232|2||-2||2|1|||-2||-2|0|3|||7496|10|||1|560917|-1|4|3|44
502551045|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-03-06|Followup|2014-02-22|2014-02-18|Complete|Done|2|1|1|1|2|3|1.67|4|1|1|2|1|4|2.17|-23.04|1|2|3|1|1|3|1.83|1|1|2|2|1|2|1.5|22|3|1|1|1.67|1|2|2|1.67|0|2|4|3|2|2.75|2|2|2|2|2|37.5|4|4|4|4|4|3|3|3.71|4|4|4|4|3|4|4|3.86|-3.89|2|4|3|3|3|4|2|3|0|2|2|2|2|2|2|0|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Health|24.4||2|2|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||54|28031|Bachelors Degree|Married|Business: Mgt, Admin|28262|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502551498|31|0|2|502864071|1|0|2|500597976|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|560956|401956|4|3|45
500186071|BBBS of Greater Charlotte|Main Office|C|Completed|2004-01-05|2014-04-30|Followup|2014-01-05|2014-02-12|Complete|Done|4|3|3|3|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|123.8||1|1|1|1|M|White||21|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||40|28277|Masters Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187670|1|0|1|500189012|1|0|1|500037012|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|561432||4|3|45
500892914|BBBS of Greater Charlotte|Main Office|C|Completed|2010-02-16|2014-09-11|Followup|2014-02-16|2014-02-15|Complete|Done|1|4|4|4|4|4|3.5|||||||||2|4|3|2|2|3|2.67|||||||||4|3|4|3.67||||||3|2|4|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||1|1||||4|4||||Red|Amachi|Child: Graduated|54.8||2|2|1|1|M|Black||20|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Sales|28269|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500893173|31|0|1|501964388|1|0|1|500429157|2||500003586||4|3|500000294|500000294|-2||-2|0|5|||7464|9|||1|561585||4|3|45
502747706|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-17|2015-10-09|Followup|2013-11-17|2013-12-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|46.7||1|1|1|1|F|Multi-Race (None of the above)||13|No|Mother|28229|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Enrollment|F|Black||34|28226|Bachelors Degree|Single|Business: Clerical|28208|0|6|Self|Self|Big|General Community|Project Big|Enrollment|277|60|598|500000170|500017777|502748616|7|0|2|502618438|31|0|2|500566066|2||-2||4|3|||-2|500004640|-2|0|10|||7464|9|||1|561609||4|1|45
502974629|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-25|2016-09-26|Baseline|2013-02-19|2013-02-25|Complete|Done|2|4|4|3|3|2|3|||||||||2|3|4|3|4|2|3|||||||||4|4|4|4||||||3|5|4|2|3.5|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|3|3.33||||||2|3|2.5|||||1|1||||4|4||||Red||Child/Family: Moved|43||1|1|1|1|M|Black||18|No|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||33|28209|Bachelors Degree|Married|Business: Mgt, Admin|28202|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502976067|31|0|1|503188801|1|0|1|500682863|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|561886|-1|4|3|44
502939347|BBBS of Greater Charlotte|Main Office|C|Completed|2014-02-25|2015-10-15|Baseline|2013-02-19|2014-02-25|Complete|Done|2|1|2|1|3|4|2.17|||||||||1|2|3|1|2|4|2.17|||||||||4|3|4|3.67||||||4|3|1|1|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green||Child/Family: Moved|19.6||1|1|1|1|F|Black||13|No|Mother|28052|Two Parent|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||32|28202|Masters Degree|Single|Medical: Doctor, Provider|28204|0|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|502940773|31|0|2|503598887|1|0|2|500748884|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|561889|-1|4|3|44
503166335|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-19|2014-09-24|Baseline|2013-02-20|2013-03-18|Complete|Done|4|3|4|4|4|4|3.83|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|18.2||2|2|1|1|F|White||14|No|Mother|28031|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|F|White||34|28031|Bachelors Degree|Single|Business: Marketing|28031|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503168022|1|0|2|503335465|1|0|2|500683005|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|562235|-1|4|3|44
501295538|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-30|NaT|Followup|2014-03-30|2014-04-03|Complete|Done|4|3|2|3|3|3|3|||||||||2|3|4|2|2|4|2.83|||||||||4|4|4|4||||||4|5|2|3|3.5|||||||4|4|4|4|4|3|2|3.57||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||59.5||2|2|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||31|28078|Bachelors Degree||Medical||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500740560|31|0|2|502897530|1|0|2|500603727|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|562354||4|3|45
503034769|BBBS of Greater Charlotte|Main Office|C|Active|2014-01-31|NaT|Baseline|2013-02-20|2014-01-31|Complete|Done|3|1|4|1|4|4|2.83|||||||||2|1|4|2|2|3|2.33|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|||37.5||1|1|1|1|M|Black||13|No|Mother|28226|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|M|Black||39|28210|Some College|Single|Arts, Entertainment, Sports|28202|7|2|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503036365|31|0|1|503650997|31|0|1|500744436|2||-2||2|1|||-2||-2|0|10|||7458|9|||1|562586|-1|4|3|44
502824908|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-21|2015-07-22|Followup|2014-02-21|2014-02-19|Complete|Done|3|1|2|3|2|3|2.33|3|2|3|2|3|3|2.67|-12.73|3|4|4|1|4|4|3.33|3|4|4|2|2|3|3|11|4|3|3|3.33|4|4|4|4|-16.75|4|5|3|3|3.75|5|5|4|4|4.5|-16.67|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|4|4|-7.25|4|3|4|3.67|4|4|4|4|-8.25|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green||Child: Graduated|41||1|1|1|1|F|Black||19|No|Mother|28226|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community||Match Support|F|White||34|28226|Bachelors Degree|Married|Unknown|29715|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502826191|31|0|2|502891382|1|0|2|500596373|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|562587|399457|4|3|45
501143676|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-28|2015-07-14|Baseline|2013-02-21|2013-02-28|Complete|Done|3|3|4|1|4|4|3.17|||||||||3|4|4|2|2|3|3|||||||||3|4|4|3.67||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|28.5||1|1|1|1|M|Black||14|No|Mother|28213|One Parent: Female|$10,000 to $14,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||50|28269|Associate Degree|Married|Self-Employed, Entrepreneur||12|0|Newspaper|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501143950|31|0|1|503315012|31|0|1|500683363|2||-2||4|3|||-2|500000294|-2|34|2|||129|1|||1|562841|-1|4|3|44
502714405|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-08|2015-08-06|Followup|2014-12-08|2015-01-22|Complete|Done|3|4|3|4|3|3|3.33|3|3|2|2|3|4|2.83|17.67|3|3|3|3|2|3|2.83|2|3|3|3|4|4|3.17|-10.73|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|5|3|3|3.5|-14.29|4|4|4|4|4|4|4|4|4|3|4|4|4|4|4|3.86|3.63|3|4|4|3.67|3|4|4|3.67|0|2|2|2|1|1|1|100|2|2|1|1|100|4|4|4|4|0|Green||Child: Graduated|43.9||1|1|1|1|M|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||33|28213|Associate Degree|Single|Transport: Driver|28205|5|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500017732|502715293|31|0|1|502764673|31|0|1|500577475|2||-2||4|1||500005291|-2||-2|56|1|||7446|3|||1|563250|367813|4|3|45
502974629|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-25|2016-09-26|Followup|2014-02-25|2014-04-11|Complete|Done|3|2|4|2|3|3|2.83|2|4|4|3|3|2|3|-5.67|2|4|3|3|3|4|3.17|2|3|4|3|4|2|3|5.67|4|4|4|4|4|4|4|4|0|2|3|3|3|2.75|3|5|4|2|3.5|-21.43|4|4|4|4|4|4|4|4|4|4|4|4|3|4|4|3.86|3.63|4|4|4|4|3|4|3|3.33|20.12|3|3|3|2|3|2.5|20|2|2|1|1|100|4|4|4|4|0|Red||Child/Family: Moved|43||1|1|1|1|M|Black||18|No|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||33|28209|Bachelors Degree|Married|Business: Mgt, Admin|28202|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502976067|31|0|1|503188801|1|0|1|500682863|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|564262|561886|4|3|45
502225378|BBBS of Greater Charlotte|Main Office|C|Active|2011-01-26|NaT|Followup|2014-01-26|2014-02-25|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||73.6||1|1|1|1|M|White||14|No|Mother|28277|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||67|28277|Bachelors Degree|Divorced|Tech: Sales, Mktg||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|502225809|1|0|1|502245842|1|0|1|500509780|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|564783||4|3|45
501735420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-26|2015-08-13|Followup|2014-01-26|2014-03-12|Complete|Done|4|4|4|2|3|3|3.33|||||||||2|2|3|2|2|3|2.33|||||||||4|4|4|4||||||5|1|3|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Child: Lost interest|66.5||2|2|2|2|F|Black||16||GrandMother|28215|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||41|28277|Bachelors Degree|Single|Business: Mgt, Admin||9|0|General|Other Big|Big|General Community||Enrollment|277|60|598|500000170|500017732|501735760|31|0|2|500956022|1|0|2|500428818|2||-2||4|1|||-2||-2|6854|8|||6450|12|||1|564838||4|3|45
502663937|BBBS of Greater Charlotte|Main Office|C|Active|2013-02-27|NaT|Followup|2014-02-27|2014-02-18|Complete|Done|4|4|4|4|4|4|4|2|4|4|4|3|4|3.5|14.29|3|3|3|3|3|3|3|3|2|4|2|3|4|3|0|4|4|4|4|4|4|4|4|0|3|5|5|4|4.25|3|4|5|5|4.25|0|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|3|3.71|4.04|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green|||48.6||1|1|1|1|M|Black||15|No|Mother|28212|Two Parent|$35,000 to $39,999||No||Relative|General Community||Match Support|M|White||30|28105|Bachelors Degree|Single|Business: Sales|17001|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502664764|31|0|1|503296990|1|0|1|500684232|2||-2||2|1|||-2||-2|0|3|||7496|10|||1|565627|560917|4|3|45
502304267|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-27|2016-09-01|Followup|2014-02-27|2014-05-14|Expired|Late||||||||3|1|2|1|1|2|1.67|||||||||2|2|3|4|2|3|2.67||||||3|4|2|3|||||||5|4|3|4|4||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||3|2|2.5||||1|1|||||||Yellow||Child/Family: Lost contact with volunteer/agency|42.1||2|2|1|1|M|White||16|No|Mother|28277|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||47|28277|Bachelors Degree|Married|Business|28217|20|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502304699|1|0|1|503343217|1|0|1|500682425|2||-2||4|2|||-2||-2|0|10|||7671|13|||1|565632|194371|4|0|45
502581328|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-28|2015-07-27|Followup|2014-02-28|2014-04-01|Complete|Done|2|2|3|4|3|2|2.67|3|2|3|2|1|3|2.33|14.59|4|4|4|3|4|4|3.83|4|4|4|4|4|4|4|-4.25|4|4|4|4|4|4|4|4|0|4|5|5|5|4.75|5|5|5|5|5|-5|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|4|3.86|0|3|3|3|3|4|4|3|3.67|-18.26|3|2|2.5|4|4|4|-37.5|2|2|2|2|0|4|4|4|4|0|Yellow||Child: Lost interest|28.9||1|1|1|1|F|Black||16|No|GrandMother|28212|One Parent: Female|$20,000 to $24,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||46|28262|PHD|Single|Education: College Professor|28223|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502581832|31|0|2|503144090|31|0|2|500681651|2||-2||4|2|||-2||-2|6854|8|||7464|9|||1|565906|306034|4|3|45
500185637|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-29|2014-12-11|Followup|2013-12-29|2014-01-02|Complete|Done|3|3|4|3|3|3|3.17|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|3|3.33||||||2|4|3|||||2|2||||4|4||||Green||Child: Graduated|107.4||1|1|2|2|M|Black||20||Mother|28206|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Black||55|28297|Masters Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500187271|31|0|1|500189284|31|0|1|500073080|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|565992||4|3|45
500261295|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-21|2017-03-09|Followup|2013-12-21|2014-02-12|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|134.6||1|1|1|1|M|White||20||Mother|28104|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||60|28270|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500261310|1|0|1|500188435|1|0|1|500073081|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|565993||4|1|45
501143676|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-28|2015-07-14|Followup|2014-02-28|2014-04-30|Declined|Late||||||||3|3|4|1|4|4|3.17|||||||||3|4|4|2|2|3|3||||||3|4|4|3.67|||||||4|5|5|4|4.5||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|1|1.5||||2|2||||4|4||Red||Child/Family: Lost contact with volunteer/agency|28.5||1|1|1|1|M|Black||14|No|Mother|28213|One Parent: Female|$10,000 to $14,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||50|28269|Associate Degree|Married|Self-Employed, Entrepreneur||12|0|Newspaper|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501143950|31|0|1|503315012|31|0|1|500683363|2||-2||4|3|||-2|500000294|-2|34|2|||129|1|||1|566520|562841|4|1|45
501936316|BBBS of Greater Charlotte|Main Office|C|Completed|2010-01-28|2016-08-29|Followup|2014-01-28|2014-03-24|Declined|Late||||||||3|3|3|2|2|2|2.5|||||||||3|3||3|3|3|||||||3|3|3|3|||||||4|5|4|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2|||||||Green||Child/Family: Lost contact with volunteer/agency|79||1|1|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||54|28203|||Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|501936714|31|0|1|501872326|1|0|1|500428557|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|566652|28181|4|1|45
500997880|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-19|2016-07-29|Followup|2014-02-19|2014-03-13|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|4|3|3|2|4|3.17|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||3|3|4|3|4|4|3|3.43||||||||||4|4|3|3.67||||||2|3|2.5|||||2|2||||4|4||||Green||Child: Graduated|101.3||1|1|1|1|M|Black||18|No|Mother|28204|Two Parent|$40,000 to $44,999||Yes||Self|General Community||Match Support|M|White||33|28202|Bachelors Degree|Married|Business: Marketing||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500998153|31|0|1|500990660|1|0|1|500237316|2||-2||4|1|||-2||-2|0|10|||46|2|||1|567670||4|3|45
502876870|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-05|2016-07-28|Followup|2014-03-05|2014-03-04|Complete|Done|4|4|4|4|4|4|4|3|3|4|1|4|4|3.17|26.18|4|4|4|4|4|4|4|3|4|4|4|1|4|3.33|20.12|4|3|4|3.67|4|4|4|4|-8.25|4|3|5|4|4|5|3|4|5|4.25|-5.88|4|4|4|4|4|4|3|3.86|4|4|4|4|2|3|2|3.29|17.33|4|4|4|4|4|4|3|3.67|8.99|2|3|2.5|1|2|1.5|66.67|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Changed workplace/school partnership|40.8||2|2|1|1|F|Black||16|No|GrandMother|28206|Grandparents|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Multi-race (Asian & White)||28|60654|Bachelors Degree|Single|Business: Mgt, Admin|60601|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502878273|31|0|2|503104166|37|0|2|500684838|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|567846|405521|4|3|45
501628854|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-05|2014-10-31|Followup|2014-03-05|2014-05-20|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Moved|19.9||3|3|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||42|28205|Associate Degree|Single|Transport: Flight Attendant||8|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|501629177|31|0|2|503374490|31|0|2|500682899|2||500003586||4|2||500000294|-2|500000294|-2|0|10|||7464|9|||1|568121||4|0|45
502873189|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-21|2016-09-01|Followup|2013-03-21|2013-05-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|53.4||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||40|28216|Masters Degree|Single|Finance||6|0|Charlotte Cares|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502874592|31|0|2|502882530|31|0|2|500600322|2||-2||4|2|||-2||-2|0|4|||11246|6|||1|568264||4|1|45
500577150|BBBS of Greater Charlotte|Main Office|C|Active|2011-03-22|NaT|Followup|2014-03-22|2014-03-31|Complete|Done|4|2|4|2|3|4|3.17|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||2|2|5|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||2|3|1|2||||||3|2|2.5|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI||71.8||4|5|1|2|F|Black||15||Aunt|28213|One Parent: Female|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||40|29715|||Customer Service||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500214349|31|0|2|501734288|1|0|2|500526894|2||500004641||2|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|568543||4|3|45
502787524|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-25|2014-08-29|Followup|2014-01-25|2014-03-10|Declined|Done||||||||3|4|4|4|4|4|3.83|||||||||2|4|3|4|4|4|3.5||||||4|3|3|3.33|||||||4|5|5|5|4.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4|||||||||4|4||Red||Child/Family: Lost contact with volunteer/agency|31.1||1|1|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28205|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Asian||29|28202||Single|Tech: Computer/Programmer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502788707|38|0|2|502272989|4|0|2|500587325|2||-2||4|3|||-2|500004640|-2|0|10|||7496|10|||1|568711|382987|4|1|45
502328599|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-22|2014-10-31|Followup|2014-02-22|2014-04-08|Declined|Done||||||||4|1|4|1|4|3|2.83|||||||||2|4|4|2|2|4|3||||||2|2|2|2|||||||4|3|4|5|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|4|3||||2|2||||4|4||Red||Volunteer: Time constraint|32.3||1|1|1|1|M|Black||15|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|M|White||73|28226|Bachelors Degree|Widowed|Construction||7|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502329034|31|0|1|502732347|1|0|1|500594124|2||-2||4|3|||-2||-2|0|10|||131|1|||1|568712|376848|4|1|45
501712048|BBBS of Greater Charlotte|Main Office|C|Active|2011-02-22|NaT|Followup|2014-02-22|2014-02-25|Complete|Done|1|2|4|4|4|4|3.17|||||||||2|4|3|4|4|4|3.5|||||||||4|2|2|2.67||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green|Amachi||72.7||1|1|1|1|M|Black||13|Yes|Mother|28134|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||29|28273|Some College|Single|Govt: Mgmt/Admin|28208|2|0|Relative|Relative|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|501712386|31|0|1|502405439|1|0|1|500516322|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||17161|11|||1|569030||4|3|45
502317500|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-08|2015-07-31|Followup|2014-02-08|2014-03-26|Declined|Late||||||||4|2|1|2|4|4|2.83|||||||||2|3|4|2|2|4|2.83||||||4|4|4|4|||||||4|3|2|3|3||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||3|2|2.5||||2|2||||4|4||Red|Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|41.7||1|1|2|2|M|Black||15|No|Mother|28214|One Parent: Female|Unknown||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|M|White||33|28214|Associate Degree|Single|Law: Security Officer|28208|2|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502317931|31|0|1|502658498|1|0|1|500587614|2||-2||4|3|500004640, 500004901|500004640, 500004901|-2||-2|0|4|||7464|9|||1|569099|383492|4|1|45
502051702|BBBS of Greater Charlotte|Main Office|C|Active|2013-04-16|NaT|Baseline|2013-03-08|2013-04-16|Complete|Done|3|3|4|3|1|3|2.83|||||||||1|4|3|2|1|4|2.5|||||||||4|4|4|4||||||5|4|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi||47||1|1|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||31|28262|Bachelors Degree|Single|Finance|28281|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501977740|31|0|2|503378835|31|0|2|500690864|2||-2||2|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|569232|-1|4|3|44
503296945|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-13|2015-04-06|Baseline|2013-03-08|2013-03-13|Complete|Done|3|3|4|3|3|3|3.17|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||2|3|4|4|3.25|||||||4|3|4|4|4|4|3|3.71||||||||||3|4|3|3.33||||||4|3|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|24.8||1|1|1|1|M|Black||16|Yes|Mother|28273|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||43|29707|Bachelors Degree|Separated|Govt||10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503298770|31|0|1|503381327|31|0|1|500687021|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|569268|-1|4|3|44
503225805|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-08|2016-05-24|Followup|2014-03-08|2014-03-06|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|3|3|2|3|3|2.83|||||||||4|4|4|4||||||3|4|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|4|2.5|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|38.5||1|1|1|1|F|White||16|No|Mother|28082|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|F|White||33|28138|Associate Degree|Divorced|Insurance||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503227593|1|0|2|503317460|1|0|2|500680855|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|569389|503767|4|3|45
501788776|BBBS of Greater Charlotte|Main Office|C|Active|2010-01-25|NaT|Followup|2014-01-25|2014-01-22|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi||85.7||1|1|1|1|M|Black||14|Yes|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||64|28117||Married|Business: Sales|28031|0|0|Alpha Kappa Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500020752|501789128|31|0|1|501698382|1|0|1|500418170|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||8697|14|||1|569580||4|3|45
500824037|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-15|NaT|Followup|2014-03-15|2014-03-17|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|||120||1|1|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community||Match Support|F|White||34|28210|Bachelors Degree|Single|Education: Teacher|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500824306|31|0|2|500789337|1|0|2|500165956|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|569719||4|3|45
500185601|BBBS of Greater Charlotte|Main Office|C|Completed|2008-01-28|2015-07-23|Followup|2014-01-28|2014-02-06|Complete|Done|4|3|4|2|4|4|3.5|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Graduated|89.8||2|2|1|1|M|Black||20||Mother|28210|Other/Unknown|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28078|High School Graduate|Single|Finance: Accountant|28202|0|4|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|500187235|31|0|1|501082220|1|0|1|500236473|2||-2||4|1|||-2||-2|6854|8|||7458|9|||1|569940||4|3|45
501516900|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-28|2015-08-27|Followup|2014-01-28|2014-01-16|Complete|Done|3|3|2|3|2|2|2.5|||||||||3|4|3|4|4|3|3.5|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|2|2.5|||||2|2||||4|4||||Green||Child: Graduated|78.9||1|1|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||39|28212|Bachelors Degree|Single|Medical: Healthcare Worker|28210|1|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500018987|501517192|31|0|2|501438601|31|0|2|500332399|2||-2||4|1|||-2||-2|6854|8|||7462|13|||1|569941||4|3|45
502979759|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-12|2016-02-10|Followup|2014-03-12|2014-04-30|Declined|Late||||||||4|1|4|1|4|4|3|||||||||2|3|3|3|4|3|3||||||4|4|4|4|||||||4|5|4|3|4||||||||||4|4|4|4|4|4|4|4||||||4|3|4|3.67|||||2|4|3||||1|1||||4|4||Yellow||Child/Family: Lost contact with volunteer/agency|35||1|1|1|1|M|Black||16||Mother|28211|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||29|28211|Bachelors Degree||Construction|28208|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|502981210|31|0|1|503234517|1|0|1|500682418|2||-2||4|2|||-2||-2|0|10|||46|2|||1|570163|552522|4|1|45
503110829|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-27|2016-05-24|Baseline|2013-03-12|2013-03-20|Complete|Done|2|4|3|3|3|4|3.17|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||1|1||||4|4||||Yellow||Volunteer: Moved|37.9||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|$45,000 to $49,999||No||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Mgt, Admin|28217|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503112489|31|0|1|503130981|1|0|1|500687926|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|570189|-1|4|3|44
501811385|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-23|2016-08-19|Followup|2014-03-23|2014-03-24|Complete|Done|4|3|1|1|4|3|2.67|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red|2010-2012 OJJDP JJI, Cabarrus County|Child: Graduated|64.9||2|2|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||43|28075|Bachelors Degree|Married|Business: Mgt, Admin||7|0|Recruitment Event|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501811730|31|0|2|502460013|31|0|2|500524684|2||-2||4|3|500005291, 500016374|500016374|-2|500016374|-2|6854|8|||7459|10|||1|570326||4|3|45
500186905|BBBS of Greater Charlotte|Main Office|C|Completed|2005-02-10|2015-11-04|Followup|2014-02-10|2014-02-10|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|1|1|||||2|2||||4|4||||Red|Amachi|Child: Graduated|128.8||1|1|1|1|F|Black||19|Yes|Mother|28205|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|F|Black||50|28215|Some College|Single|Finance: Banking||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188151|31|0|2|500189677|31|0|2|500037790|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||7453|7|||1|570506||4|3|45
501361902|BBBS of Greater Charlotte|Main Office|C|Active|2009-01-23|NaT|Followup|2014-01-23|2014-01-22|Complete|Done|4|4|3|3|3|4|3.5|||||||||3|4|3|3|3|4|3.33|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi||97.7||1|1|1|1|M|White||17|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28227|Bachelors Degree|Divorced|Business: Sales|28273|9|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501249611|1|0|1|501307192|1|0|1|500328424|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|570614||4|3|45
502275241|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-21|2015-10-15|Followup|2014-03-21|2014-03-24|Complete|Done|3|4|4|4|4|1|3.33|4|3|3|3|4|3|3.33|0|2|4|4|2|4|4|3.33|3|3|4|3|3|2|3|11|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|2|3|3|3|2.75|18.18|4|4|4|4|3|4|4|3.86|4|4|4|4|4|||||3|3|4|3.33|3|3|3|3|11|3|2|2.5|3|3|3|-16.67|2|2|2|2|0|4|4||||Green|Amachi|Child: Lost interest|54.8||1|1|1|1|F|Black||17|No|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||26|28031|Bachelors Degree|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|502275673|31|0|2|502394690|1|0|2|500521625|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7496|10|||1|570727|235273|4|3|45
503296945|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-13|2015-04-06|Followup|2014-03-13|2014-05-20|Declined|Late||||||||3|3|4|3|3|3|3.17|||||||||2|4|3|3|3|3|3||||||4|4|4|4|||||||2|3|4|4|3.25||||||||||4|3|4|4|4|4|3|3.71||||||3|4|3|3.33|||||4|3|3.5||||2|2||||4|4||Green||Volunteer: Lost contact with child/agency|24.8||1|1|1|1|M|Black||16|Yes|Mother|28273|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||43|29707|Bachelors Degree|Separated|Govt||10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503298770|31|0|1|503381327|31|0|1|500687021|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|570903|569268|4|1|45
502875279|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-19|2014-12-17|Followup|2014-03-19|2014-04-24|Complete|Done|3|2|1|1|3|1|1.83|3|2|2|2|3|3|2.5|-26.8|4|4|3|1|2|3|2.83|3|4|3|4|1|2|2.83|0|4|4|4|4|4|4|4|4|0|4|3|4|4|3.75|3|3|4|5|3.75|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|3|3.67|4|4||||3|2|2.5|3|2|2.5|0|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Time constraint|33||2|2|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||32|28210|Bachelors Degree|Single|Business: Sales||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502876679|31|0|2|502864263|31|0|2|500600651|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|571488|406736|4|3|45
503373647|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-21|2014-02-06|Baseline|2013-03-15|2013-03-21|Complete|Done|3|1|2|1|3|4|2.33|||||||||2|2|3|2|1|3|2.17|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||1|1||||4|4||||Yellow||Child/Family: Moved|10.6||1|1|2|2|F|Black||16|No|Mother|28213|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||30|28213|Some College|Single|Medical|28209|1|4|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500015820|503375503|31|0|2|503377601|31|0|2|500688140|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|571499|-1|4|3|44
500948129|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-18|2016-06-30|Followup|2014-03-18|2014-03-13|Complete|Done|3|3|4|3|3|3|3.17|||||||||2|3|4|3|2|4|3|||||||||4|4|4|4||||||4|4|5|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|75.4||2|2|1|1|F|Black||18|No|Mother|28217|One Parent: Female|$25,000 to $29,999|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||40|28203|Some College|Living w/ Significant Other|Finance: Banking|28281|1|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501891556|1|0|2|500438403|2||500003586||4|1|500000294|500000294|-2||-2|34|2|||7464|9|||1|571854||4|3|45
502106926|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-18|2014-09-24|Followup|2014-03-18|2014-06-02|Expired|Late||||||||4|4|4|1|2|4|3.17|||||||||1|2|4|3|3|3|2.67||||||4|4|4|4|||||||5|1|5|1|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Green||Child/Family: Moved|18.2||2|2|1|1|M|Black||17|No|Mother|28031|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||53|28036|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0||Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502107353|31|0|1|503230500|1|0|1|500686913|2||-2||4|1|||-2||-2|0|10|||0|11|||1|572232|40460|4|0|45
502278985|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-01|NaT|Followup|2014-03-01|2014-04-14|Complete|Done|3|4|4|2|3|3|3.17|||||||||4|3|2|3|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|3|2.5|||||2|2||||4|4||||Green|Project Big||60.5||1|1|2|2|M|Black||14|No|Mother|28213|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||40|28269||Married|Business: Marketing||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502279417|31|0|1|500220237|31|0|1|500599107|2||-2||2|1|500004640||-2|500000294|-2|6854|8|||2238|7|||1|572304||4|3|45
502211307|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-03|2014-04-24|Followup|2014-02-03|2014-03-23|Declined|Late||||||||4|4|4|3|4|3|3.67|||||||||4|3|3|4|3|3|3.33||||||4|4|4|4|||||||4|4|4||||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4||||||3|||||2|2|||||||Yellow|Amachi|Volunteer: Time constraint|38.6||1|1|1|1|M|Black||16|Yes|Mother|28278|One Parent: Female|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||51|28214|Bachelors Degree|Single|Business: Sales|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502211737|31|0|1|502371462|1|0|1|500512414|2||-2||4|2|500000294|500000294|-2|500000294|-2|7016|11|||7496|10|||1|572330|177660|4|1|45
500185630|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-19|2014-09-18|Followup|2014-03-19|2014-03-18|Complete|Done|3|4|3|2|3|3|3|||||||||2|3|3|3|2|3|2.67|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|18||3|3|2|2|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||39|28211|High School Graduate|Single|Finance: Banking|28208|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500015820|500187264|31|0|2|500542491|31|0|2|500688663|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|572493||4|3|45
503166335|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-19|2014-09-24|Followup|2014-03-19|2014-05-03|Complete|Done|4|3|4|3|4|4|3.67|4|3|4|4|4|4|3.83|-4.18|2|4|3|3|2|3|2.83|4|4|4|4|2|4|3.67|-22.89|4|3|3|3.33|4|4|4|4|-16.75|3|3|3|3|3|5|4|5|5|4.75|-36.84|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|2|2.5|4|4|4|-37.5|||2|2||4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|18.2||2|2|1|1|F|White||14|No|Mother|28031|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|F|White||34|28031|Bachelors Degree|Single|Business: Marketing|28031|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503168022|1|0|2|503335465|1|0|2|500683005|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|572539|562235|4|3|45
502866083|BBBS of Greater Charlotte|Main Office|C|Active|2013-03-26|NaT|Baseline|2013-03-19|2013-03-26|Complete|Done|3|3|2|3|2|3|2.67|||||||||3|3|4|1|4|3|3|||||||||3|4|4|3.67||||||5|4|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||2|2|2|||||1|1||||4|4||||Green|||47.7||1|1|1|1|M|White||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||32|28104|Bachelors Degree|Single|Business|20785|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502867478|1|0|1|503378884|1|0|1|500688846|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|572802|-1|4|3|44
502858216|BBBS of Greater Charlotte|Main Office|C|Active|2013-03-19|NaT|Followup|2014-03-19|2014-04-15|Complete|Done|4|2|2|1|2|2|2.17|4|1|4|1|4|4|3|-27.67|2|4|3|1|3|3|2.67|3|3|4|4|2|4|3.33|-19.82|4|4|4|4|4|4|4|4|0|4|3|3|3|3.25|4|3|2|2|2.75|18.18|2|4|4|4|4|4|4|3.71|4|4|4|4|4|4|3|3.86|-3.89|3|3|3|3|4|4|4|4|-25|1|3|2|2|2|2|0|2|2|1|1|100|4|4|4|4|0|Green|||47.9||1|1|1|1|M|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||32|29708|Bachelors Degree|Married|Finance||0|9|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020752|502859613|31|0|1|503376842|1|0|1|500687641|2||-2||2|1|||-2||-2|0|10|||7438|1|||1|572815|491466|4|3|45
501340097|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-23|2016-09-19|Followup|2014-03-23|2014-03-23|Complete|Done|3|4|4|2|4|4|3.5|||||||||4|4|4|2|4|3|3.5|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|77.9||2|2|1|1|M|Multi-race (Black & Hispanic)||17|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Hispanic||28|28277|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501340376|38|0|1|501934966|3|0|1|500440292|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|572977||4|3|45
500799303|BBBS of Greater Charlotte|Main Office|C|Completed|2007-03-27|2016-08-19|Followup|2014-03-27|2014-03-26|Complete|Done|3|3|3|2|3|4|3|||||||||3|4|3|3|3|3|3.17|||||||||4|3|4|3.67||||||3|4|4|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Red||Child: Graduated|112.8||1|1|1|1|M|White||19|No|Mother|28081|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||46|28202||Single|Business: Sales||0|4|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500799571|1|0|1|500798390|1|0|1|500167062|2||-2||4|3||500016374|-2|500016374|-2|34|2|||7464|9|||1|573470||4|3|45
501833031|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2015-11-04|Followup|2014-02-28|2014-03-20|Complete|Done|4|4|4|2|4|4|3.67|3|3|1|4|4|4|3.17|15.77|2|4|4|2|4|4|3.33|2|2|3|2|4|4|2.83|17.67|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Red|2010-2012 OJJDP JJI|Volunteer: Moved|56.2||1|1|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28205|Masters Degree|Single|Medical: Doctor, Provider|28277|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502427342|1|0|2|500518294|2||-2||4|3|500005291|500005291|-2||-2|0|10|||7464|9|||1|574188|157600|4|3|45
501833026|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-02|2016-09-30|Followup|2014-03-02|2014-03-04|Complete|Done|2|4|2|4|3|1|2.67|2|4|4|3|1|3|2.83|-5.65|2|4|4|2|3|4|3.17|2|1|3|2|3|2|2.17|46.08|4|4|4|4|4|4|4|4|0|2|5|4|4|3.75|3|4|3|3|3.25|15.38|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|2|3|33.33|3|3|3|2|4|3|0|2|2|1|1|100|4|4|4|4|0|Yellow|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|67||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28205|Masters Degree|Single|Education: Teacher|2122|1|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501833394|31|0|2|502451325|1|0|2|500518305|2||-2||4|2|500005291|500005291|-2|500000294|-2|0|10|||7464|9|||1|574189|157601|4|3|45
501132052|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-08|2015-10-15|Followup|2014-02-08|2014-04-15|Blank|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|44.2||2|3|1|2|F|Black||17||Mother|28213|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||35|85254|Bachelors Degree|Married|Medical: Admin|28217|2|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500018987|501076355|31|0|2|501356464|1|0|2|500597097|2||-2||4|1|||-2||-2|0|4|||7446|3|||1|574275||4|3|45
502610186|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-26|NaT|Followup|2014-03-26|2014-04-08|Complete|Done|4|1|4|1|4|4|3|4|1|4|1|4|4|3|0|2|4|3|2|4|4|3.17|3|3|3|2|2|3|2.67|18.73|4|4|4|4|4|4|4|4|0|2|3|3|3|2.75|2|4|2|4|3|-8.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|3|3|3|3|33.33|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Green|||59.7||1|1|1|1|F|Black||16|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Asian||35|28210|Masters Degree|Married|Arts, Entertainment, Sports|28202|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|502610737|31|0|2|502913393|4|0|2|500601697|2||-2||2|1|||-2||-2|6854|8|||7671|13|||1|574381|388768|4|3|45
501806165|BBBS of Greater Charlotte|Main Office|C|Active|2009-08-06|NaT|Followup|2013-08-06|2013-08-07|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||91.3||1|1|1|1|M|Black||12|Yes|GrandMother|28273|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|Black||40|28273|No High School|Single|Business: Human Resources||2|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500020752|501806520|31|0|1|501706064|31|0|1|500375643|2||-2||2|1|500000294|500000294|-2||-2|0|10|||7446|3|||1|574392||4|3|45
501074345|BBBS of Greater Charlotte|Main Office|C|Active|2008-03-31|NaT|Followup|2014-03-31|2014-03-31|Complete|Done|4|1|4|1|4|4|3|||||||||1|1|4|2|1|4|2.17|||||||||4|4|4|4||||||2|2|3|4|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi, Cabarrus County||107.5||1|1|1|1|M|White||16|Yes|GrandMother|28025|Grandparents|Unknown||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|White||46|28027|Bachelors Degree|Divorced|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501074618|1|0|1|501158523|1|0|1|500250038|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|5635|9|||46|2|||1|574566||4|3|45
502124485|BBBS of Greater Charlotte|Main Office|C|Active|2013-03-25|NaT|Followup|2014-03-25|2014-04-15|Complete|Done|3|3|2|3|3|3|2.83|4|1|2|1|2|4|2.33|21.46|2|3|3|3|2|3|2.67|3|4|4|4|4|4|3.83|-30.29|4|4|4|4|4|4|4|4|0|4|4|4|4|4|5|5|5|5|5|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|3|3|4|4|4|4|-25|3|3|3|2|4|3|0|2|2|2|2|0|4|4||||Green|||47.7||2|2|2|2|F|Black||17|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|502142970|31|0|2|501905673|31|0|2|500689671|2||-2||2|1|||-2||-2|0|4|||7496|10|||1|574570|132622|4|3|45
502725760|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2014-09-24|Followup|2014-01-23|2014-04-09|Expired|Late||||||||4|4|4|4|4|4|4|||||||||2|4|4|2|4|4|3.33||||||4|4|4|4|||||||5|4|4|5|4.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|2|3||||2|2||||4|4||Yellow|Amachi|Volunteer: Lost contact with child/agency|32||1|1|1|1|M|Black||16|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community|Amachi|Match Support|M|Black||28|28226|Bachelors Degree|Single|Business: Sales|28217|0|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502726656|31|0|1|502687867|31|0|1|500589763|2||-2||4|2|500000294|500000294|-2||-2|0|10|||4748|14|633|1|1|574785|388386|4|0|45
502825916|BBBS of Greater Charlotte|Main Office|C|Active|2012-01-23|NaT|Followup|2014-01-23|2014-04-09|Expired|Late||||||||4|2|1|2|2|4|2.5|||||||||2|3|4|3|4|3|3.17||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||4|4|4||||2|2||||4|4||Yellow|Amachi||61.7||1|1|2|2|F|Black||14|Yes|Mother|28273|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28208|Some College|Single|Education: Teacher|28226|1|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502827199|31|0|2|502367677|31|0|2|500589764|2||-2||2|2|500000294|500000294|-2|500000294, 500004640|-2|0|10|||7464|9|||1|574786|388387|4|0|45
502725777|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-23|2015-08-30|Followup|2014-01-23|2014-04-09|Expired|Late||||||||3|3|2|3|1|4|2.67|||||||||3|4|4|4|4|4|3.83||||||4|4|4|4|||||||3|5|3|3|3.5||||||||||4|4|4|4|4|4|2|3.71||||||4|4|3|3.67|||||4|4|4||||1|1||||4|4||Red|Amachi|Volunteer: Moved|43.2||1|1|1|1|F|Black||17|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||31|28217||Single|Customer Service||0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502726673|31|0|2|502710032|31|0|2|500590950|2||-2||4|3|500000294|500000294|-2||-2|34|2|||7464|9|||1|574787|390244|4|0|45
502866079|BBBS of Greater Charlotte|Main Office|C|Active|2013-03-26|NaT|Followup|2014-03-26|2014-03-31|Complete|Done|4|2|4|3|4|4|3.5|4|1|1|1|1|1|1.5|133.33|4|4|4|4|4|4|4|4|4|4|3|4|4|3.83|4.44|4|4|4|4|4|4|4|4|0|5|4|4|4|4.25|5|5|4|3|4.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|2|3|3|2.67|1|3|1|1.67|59.88|3|1|2|4|1|2.5|-20|2|2|2|2|0|4|4|4|4|0|Green|||47.7||1|1|1|1|M|White||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||32|28210|Bachelors Degree|Single|Business: Sales||4|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|502867478|1|0|1|503378886|1|0|1|500686789|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|574907|539346|4|3|45
502866083|BBBS of Greater Charlotte|Main Office|C|Active|2013-03-26|NaT|Followup|2014-03-26|2014-04-07|Complete|Done|3|2|3|3|2|3|2.67|3|3|2|3|2|3|2.67|0|3|3|4|4|4|4|3.67|3|3|4|1|4|3|3|22.33|4|4|3|3.67|3|4|4|3.67|0|4|5|4|5|4.5|5|4|3|4|4|12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|3|3.33|3|4|2|3|11|3|2|2.5|2|2|2|25|2|2|1|1|100|4|4|4|4|0|Green|||47.7||1|1|1|1|M|White||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||32|28104|Bachelors Degree|Single|Business|20785|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502867478|1|0|1|503378884|1|0|1|500688846|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|574912|572802|4|3|45
502945480|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-29|NaT|Followup|2014-03-29|2014-03-25|Complete|Done|1|4|4|4|3|4|3.33|1|4|3|1|4|4|2.83|17.67|3|4|3|4|2|3|3.17|1|4|3|3|2|2|2.5|26.8|4|4|4|4|4|4|4|4|0|2|4|4|3|3.25|5|5|3|4|4.25|-23.53|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|3|3.67|8.99|2|3|2.5|1|3|2|25|1|1|2|2|-50|4|4|4|4|0|Green|||59.6||1|1|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||54|28262|Bachelors Degree|Single|Business: Mgt, Admin||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502946906|31|0|2|502919780|31|0|2|500603409|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|574961|411819|4|3|45
503246887|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-10|2016-05-25|Baseline|2013-03-27|2013-04-10|Complete|Done|3|4|4|4|1|4|3.33|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|1|2.5|||||1|1||||4|4||||Green|Amachi|Volunteer: Moved|37.5||1|1|1|1|M|Black||15|No|Mother|28212|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||27|28209|Bachelors Degree|Single|Finance|28255|1|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|503248691|31|0|1|503253208|1|0|1|500690197|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||46|2|||1|575539|-1|4|3|44
503110829|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-27|2016-05-24|Followup|2014-03-27|2014-05-10|Complete|Done|3|2|3|2|3|3|2.67|2|4|3|3|3|4|3.17|-15.77|2|3|3|3|3|3|2.83|4|4|4|1|4|4|3.5|-19.14|3|3|3|3|4|4|4|4|-25|3|3||3||5|4|4|5|4.5||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|2|4|3|0|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Moved|37.9||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|$45,000 to $49,999||No||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Mgt, Admin|28217|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503112489|31|0|1|503130981|1|0|1|500687926|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|575634|570189|4|3|45
501631547|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2016-07-29|Followup|2014-03-31|2014-03-31|Complete|Done|4|3|3|3|3|3|3.17|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||5|3|4|3|3.75|||||||4|4|4|3|3|4|2|3.43||||||||||3|3|3|3||||||4|3|3.5|||||2|2||||4|4||||Green|Project Big, 2010-2012 OJJDP JJI|Child: Graduated|64||2|2|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||38|28277|Bachelors Degree|Single|Arts, Entertainment, Sports|28203|3|6|UnitedMethodistChrch|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|501631870|31|0|1|502170945|1|0|1|500528464|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||8529|7|||1|575650||4|3|45
501597169|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-06|2016-05-31|Followup|2014-04-06|2014-05-27|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Agency: Challenges with program/partnership|85.8||1|1|1|1|M|Black||13||Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||54|28262|High School Graduate|Married|Disabled||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501597489|31|0|1|501563612|31|0|1|500352827|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|575652||4|1|45
502700503|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-30|NaT|Followup|2014-03-30|2014-03-26|Complete|Done|3|4|4|4|4|4|3.83|4|1|1|1|3|1|1.83|109.29|2|4|4|4|4|4|3.67|2|3|3|2|2|2|2.33|57.51|4|4|4|4|4|4|4|4|0|4|4|3|3|3.5|3|2|2|3|2.5|40|4|4|4|4|4|4|4|4|4|4|4|4||4|3|||4|4|3|3.67|4|4|4|4|-8.25|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|||59.5||1|1|1|1|M|Black||14|No|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||36|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502701348|31|0|1|502931327|1|0|1|500605634|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|575659|415426|4|3|45
502571727|BBBS of Greater Charlotte|Main Office|C|Completed|2012-01-13|2017-03-09|Followup|2014-01-13|2014-03-30|Expired|Late||||||||3|4|4|3|1|4|3.17|||||||||2|4|2|3|4|3|3||||||4|4|4|4|||||||4|3|4|5|4||||||||||4|4|4|4|3|4|4|3.86||||||4|4|2|3.33|||||3|4|3.5||||2|2||||4|4||Green||Volunteer: Lost contact with child/agency|61.8||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|M|Black||45|28207|Masters Degree|Married|Tech: Management|28081|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|502572181|31|0|1|502769619|31|0|1|500586830|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|576878|382185|4|0|45
502643010|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-30|2014-07-31|Followup|2014-03-30|2014-06-14|Expired|Late||||||||3|4|4|4|1|1|2.83|||||||||3|3|3|4|2|3|3||||||4|4|4|4|||||||3|4|3|4|3.5||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|3|3||||1|1||||4|4||Yellow||Volunteer: Lost contact with child/agency|16||1|1|1|1|M|Black||14|Yes|Mother|28262|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Enrollment|M|Black||30|28203|Bachelors Degree|Single|Finance|28255|3|5|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502643706|31|0|1|503262615|31|0|1|500686907|2||500003586||4|2||500000294|-2|500000294|-2|6854|8|||6247|12|||1|576973|484989|4|0|45
502740493|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-12|2013-07-31|Followup|2013-04-12|2013-06-17|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|15.6||1|1|1|1|M|Black||12|No|Mother|28214|One Parent: Female|$60,000 to $74,999||Yes||Relative|General Community||Match Support|M|Black||45|28217|High School Graduate|Separated|Transport: Driver||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500008321|502741396|31|0|1|502875462|31|0|1|500605781|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|577028||4|1|45
501011735|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-11|2015-03-05|Followup|2014-04-11|2014-04-09|Complete|Done|3|4|4|3|3|4|3.5|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Yellow|2010-2012 OJJDP JJI|Child: Lost interest|46.8||3|3|1|1|F|Black||17||Mother|28215|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28215|High School Graduate|Married|Finance: Banking|28255|13|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|277|60|598|500000170|500012459|500417756|31|0|2|502473442|31|0|2|500528270|2||-2||4|2|500005291|500005291|-2||-2|0|10|||7446|3|||1|577350||4|3|45
502893765|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-08|2015-05-11|Followup|2014-03-08|2014-03-16|Complete|Done|1|4|4|4|3|4|3.33|4|4|4|2|3|3|3.33|0|3|4|3|4|2|3|3.17|3|3|3|3|3|3|3|5.67|4|4|4|4|4|4|4|4|0|2|4|4|3|3.25|2|2|3|3|2.5|30|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|2|4|3|3|33.33|2|3|2.5|2|2|2|25|1|1|1|1|0|4|4|4|4|0|Green||Child: Graduated|38.1||1|1|1|1|F|Black||19|No|Mother|28213|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||32|28262|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502895172|31|0|2|502874079|31|0|2|500599963|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|577448|405542|4|3|45
502912141|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-05|2016-06-17|Followup|2014-04-05|2014-04-05|Complete|Done|3|4|4|3|4|4|3.67|2|4|4|3|4|4|3.5|4.86|2|4|3|2|2|4|2.83|2|4|3|2|2|4|2.83|0|4|4|4|4|4|4|4|4|0|4|5|4|5|4.5|3|4|5|5|4.25|5.88|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|4|4|-7.25|4|4|4|4|4||3|||3|2|2.5|4||||2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Moved|50.4||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Business: Marketing|28203|0|8|Other Church Partner|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|502913549|31|0|2|502932948|1|0|2|500605880|2||-2||4|3|||-2||-2|34|2|||7453|7|||1|577451|415863|4|3|45
503230648|BBBS of Greater Charlotte|Main Office|C|Active|2013-07-17|NaT|Baseline|2013-04-02|2013-07-17|Complete|Done|3|2|4|4|3|4|3.33|||||||||2|3|4|4|4|3|3.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|||44||1|1|1|1|F|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|Black||39|28214|Bachelors Degree|Single|Govt||1|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502841119|31|0|2|503169561|31|0|2|500700323|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|577620|-1|4|3|44
503110827|BBBS of Greater Charlotte|Main Office|C|Active|2013-04-22|NaT|Baseline|2013-04-02|2013-04-22|Complete|Done|4|4|1|4|4|4|3.5|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|||46.8||1|1|1|1|M|Black||18|Yes|Mother|28262|One Parent: Female|$45,000 to $49,999|Y|No||Self|General Community||Match Support|M|White||31|28203|Masters Degree|Single|Consultant||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503112489|31|0|1|503278385|1|0|1|500691045|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|577768|-1|4|3|44
503318449|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-06|2014-02-10|Baseline|2013-04-02|2013-05-02|Complete|Done|1|2|4|4|4|4|3.17|||||||||2|4|3|3|3|4|3.17|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|9.2||2|2|2|2|F|Black||15|No|Mother|28215|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||28|28213|Masters Degree|Single|Student: College||0|0||Law Student Association|Big|General Community||Match Support|277|60|598|500000170|500017777|503320281|31|0|2|500716763|31|0|2|500694861|2||-2||4|1|||-2||-2|0|10|||0|15|||1|577769|-1|4|3|44
500961015|BBBS of Greater Charlotte|Main Office|C|Completed|2008-04-11|2014-10-02|Followup|2014-04-11|2014-05-08|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|77.7||1|1|1|1|M|Black||20|Yes|Mother|28227|Two Parent|Unknown||No||Self|General Community|Amachi|Match Support|M|Black||43|28104||Married|Tech: Computer/Programmer|29607|10|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500013781|500934638|31|0|1|501210561|31|0|1|500257073|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||17161|11|||1|578005||4|3|45
501376745|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-01|2016-01-11|Followup|2014-04-01|2014-04-17|Complete|Done|3|4|4|3|3|3|3.33|||||||||3|3|3|2|3|3|2.83|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|4|3.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|81.3||1|1|3|4|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28269|||Business: Marketing||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|501377024|31|0|2|500725077|31|0|2|500350905|2||-2||4|1|||-2||-2|6854|8|||46|2|||1|578426||4|3|45
502681380|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-21|2014-12-18|Followup|2014-03-21|2014-04-16|Complete|Done|3|3|3|2|3|3|2.83|3|4|4|4|3|4|3.67|-22.89|3|4|3|2|3|3|3|4|4|3|4|1|4|3.33|-9.91|4|3|3|3.33|3|3|3|3|11|4|3|3|3|3.25|4|4|5|5|4.5|-27.78|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|2|3|33.33|3|2|2.5|2|3|2.5|0|1|1|2|2|-50|4|4|4|4|0|Green||Volunteer: Lost contact with child/agency|32.9||1|1|1|1|M|White||14|No|Mother|28075|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|M|White||29|28277|Bachelors Degree|Single|Insurance|28262|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502682208|1|0|1|502847991|1|0|1|500603939|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|578434|412646|4|3|45
502813442|BBBS of Greater Charlotte|Main Office|C|Active|2013-04-04|NaT|Followup|2014-04-04|2014-04-03|Complete|Done|4|4|4|2|3|4|3.5|4|4|4|2|3|4|3.5|0|3|3|4|2|3|4|3.17|4|4|4|2|4|4|3.67|-13.62|4|4|4|4|4|4|4|4|0|3||4|||5|5|5|4|4.75||4|4|4|4|3|4|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Green|||47.4||1|2|1|2|M|Hispanic|Mexican|15|No|Mother|28031|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28036|Some College|Married|Self-Employed, Entrepreneur|28036|20|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|502814719|3|10|1|502656402|1|0|1|500690220|2||-2||2|1||500005291|-2||-2|0|4|||7671|13|||1|578438|362674|4|3|45
501428903|BBBS of Greater Charlotte|Main Office|C|Completed|2009-01-21|2015-02-25|Followup|2014-01-21|2014-04-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|73.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|White||53|15001|Masters Degree|Single|Consultant|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501429188|31|0|1|501441245|1|0|1|500331206|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|579204||4|0|45
500887862|BBBS of Greater Charlotte|Main Office|C|Active|2011-04-13|NaT|Followup|2014-04-13|2014-04-14|Complete|Done|3|3|3|2|4|3|3|||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|3|2|||||2|2||||4|4||||Green|Cabarrus County||71.1||2|2|2|2|F|Black||18|Yes|Mother|28025|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|F|Black||43|28027||Divorced|Finance: Banking||0|7|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500888132|31|0|2|500923430|31|0|2|500530980|2||500016307||2|1|500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|579309||4|3|45
503246887|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-10|2016-05-25|Followup|2014-04-10|2014-05-24|Complete|Done|3|2|4|3|3|4|3.17|3|4|4|4|1|4|3.33|-4.8|2|4|4|4|4|4|3.67|4|3|4|4|4|4|3.83|-4.18|3|3|3|3|4|4|4|4|-25|4|4||3||5|4|4|4|4.25||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|2|4|3|4|1|2.5|20|2|2|1|1|100|4|4|4|4|0|Green|Amachi|Volunteer: Moved|37.5||1|1|1|1|M|Black||15|No|Mother|28212|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||27|28209|Bachelors Degree|Single|Finance|28255|1|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|503248691|31|0|1|503253208|1|0|1|500690197|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||46|2|||1|580262|575539|4|3|45
502431164|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-30|2015-10-12|Followup|2014-03-30|2014-04-07|Complete|Done|4|4|4|4|4|4|4|4|4|4|3|4|4|3.83|4.44|4|4|4|4|4|1|3.5|4|4|4|4|4|4|4|-12.5|4|4|4|4|4|4|4|4|0|3|5|5|5|4.5|3|4|4|2|3.25|38.46|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|3|4|3.5|-14.29|2|2|2|2|0|4|4|4|4|0|Green||Child: Graduated|42.4||1|1|1|1|M|Black||19|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community||Match Support|M|White||59|28277|Masters Degree|Single|Tech: Computer/Programmer|28203|3|4|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502431607|31|0|1|502850528|1|0|1|500606503|2||-2||4|1|||-2||-2|0|5|||7439|1|||1|580357|417125|4|3|45
500874765|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-11|2015-07-23|Followup|2014-04-11|2014-04-15|Complete|Done|2|3|4|2|3|2|2.67|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|4|3|||||2|2||||4|4||||Green||Child: Graduated|27.4||4|4|2|2|F|Black||20|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|501755813|31|0|2|502038804|31|0|2|500692473|2||-2||4|1|||-2||-2|34|2|||7496|10|||1|580684||4|3|45
502307585|BBBS of Greater Charlotte|Main Office|C|Active|2011-03-21|NaT|Followup|2014-03-21|2014-03-21|Complete|Done|4|4|4|1|4|4|3.5|4|1|2|1|1|1|1.67|109.58|4|4|4|4|4|4|4|2|2|4|1|2|3|2.33|71.67|4|4|4|4|4|4|4|4|0|5|3|3|4|3.75|4|5|5|5|4.75|-21.05|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|3|3|3|16.67|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi||71.9||1|1|1|1|F|Black||17|Yes|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||53|28031||Divorced|Medical: Admin|28207|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500020910|502308017|31|0|2|501519450|1|0|2|500521250|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|4|||7446|3|||1|581063|251051|4|3|45
501378357|BBBS of Greater Charlotte|Main Office|C|Active|2009-02-13|NaT|Followup|2014-02-13|2014-02-26|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|2|3|4|3.5|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||97||1|1|2|2|M|Multi-race (Black & White)||18|No|Mother|28213|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Mgt, Admin|28215|10|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501378636|36|0|1|501174997|31|0|1|500339619|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|581064||4|3|45
502859604|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-26|2014-12-18|Followup|2014-03-26|2014-04-16|Complete|Done|2|4|4|4|3|4|3.5|3|4|4|3|3|4|3.5|0|2|2|2|3|3|3|2.5|4|2|4|4|4|3|3.5|-28.57|4|4|4|4|4|4|4|4|0|1|1|1|1|1|5|3|5|1|3.5|-71.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|3|3.67|0|1|1|1|3|3|3|-66.67|1|1|1|1|0|4|4|4|4|0|Green||Volunteer: Time constraint|32.8||1|1|1|1|F|Hispanic|Other Central American|19|No|Mother|28205|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Hispanic||40|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502860998|3|14|2|502863229|3|0|2|500604130|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|581068|407511|4|3|45
502030263|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2014-03-31|2014-05-22|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||83.5||1|1|1|1|M|White||15|No|Mother|29710|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community||Match Support|M|White||38|28210|||Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502030662|1|0|1|501923553|1|0|1|500438867|2||-2||2|1|||-2||-2|6855|8|||7464|9|||1|581074||4|1|45
501434147|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-31|NaT|Followup|2014-03-31|2014-05-22|Declined|Late||||||||3|1|4|3|1|3|2.5|||||||||2|4|4|4|4|4|3.67||||||4|4|4|4|||||||4|5|2|5|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||2|2|||||||Green|||83.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||26|28215|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501434432|31|0|1|501926474|31|0|1|500441566|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|581077|29966|4|1|45
502472483|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-28|2014-08-28|Followup|2014-02-28|2014-03-05|Complete|Done|4|4|4|1|4|3|3.33|3|1|4|4|1|1|2.33|42.92|2|3|3|1|2|3|2.33|2|2|3|3|4|3|2.83|-17.67|4|4|4|4|4|4|4|4|0|2|3|3|4|3|3|3|3|3|3|0|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|3|3.71|4.04|2|2|2|2|4|4|4|4|-50|3|2|2.5|2|3|2.5|0|2|2|1|1|100|4|4||||Red|Amachi|Volunteer: Time constraint|42||1|1|1|1|F|Black||18|Yes|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi|Match Support|F|White||33|28202|Bachelors Degree|Single|Education|28208|4|10|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500013781|502472930|31|0|2|502453698|1|0|2|500518061|2||500003586||4|3|500000294|500000294|-2|500004640|-2|0|10|||7464|9|||1|581287|245268|4|3|45
502051702|BBBS of Greater Charlotte|Main Office|C|Active|2013-04-16|NaT|Followup|2014-04-16|2014-06-03|Declined|Late||||||||3|3|4|3|1|3|2.83|||||||||1|4|3|2|1|4|2.5||||||4|4|4|4|||||||5|4|4|3|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Yellow|Amachi||47||1|1|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||31|28262|Bachelors Degree|Single|Finance|28281|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501977740|31|0|2|503378835|31|0|2|500690864|2||-2||2|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|582107|569232|4|1|45
501185594|BBBS of Greater Charlotte|Main Office|C|Completed|2008-02-29|2016-06-15|Followup|2014-03-01|2014-03-06|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|99.5||1|1|1|1|M|Multi-race (Black & White)||19|No|Mother|28227|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Consultant|28226|0|8|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501153366|1|0|1|500248756|2||-2||4|1|||-2||-2|0|4|||7452|6|||1|583129||4|3|45
501868921|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-31|2016-07-29|Followup|2014-03-31|2014-03-31|Complete|Done|4|4|4|4|4|4|4|3|1|1|1|1|2|1.5|166.67|4|4|3|4|2|4|3.5|3|2|4|4|4|4|3.5|0|3|2|2|2.33|4|3|3|3.33|-30.03|1|3|4|2|2.5|4|5|5|4|4.5|-44.44|4|4|4|4|4|3|3|3.71|4|4|4|4|3|3|3|3.57|3.92|2|2|1|1.67|2|4|3|3|-44.33|2|2|2|2|1|1.5|33.33|2|2|1|1|100|4|4||||Green|2010-2012 OJJDP JJI|Child/Family: Moved|64||2|2|2|2|F|Black||19|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28211||Married|Finance: Banking|28255|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501869291|31|0|2|501382633|1|0|2|500524206|2||-2||4|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|583135|4527|4|3|45
501626218|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-24|2014-12-18|Followup|2014-03-24|2014-03-31|Complete|Done|3|4|4|3|3|3|3.33|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|68.8||1|1|1|1|F|Black||20|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||30|11215|Bachelors Degree|Single|Consultant|11215|0|5|other|College Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501622822|31|0|2|501587214|31|0|2|500350222|2||-2||4|1|||-2|500000294|-2|0|10|||7670|5|||1|583137||4|3|45
503346838|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-29|2013-11-08|Baseline|2013-04-19|2013-05-21|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|4|5|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Yellow||Child/Family: Unrealistic expectations|5.4||1|1|1|1|M|Black||15|Yes|Mother|28213|One Parent: Female|$50,000 to $59,999|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||49|28078|Masters Degree|Divorced|Finance||0|3|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500004169|503348683|31|0|1|503369070|1|0|1|500693781|2||-2||4|2||500000294|-2||-2|34|2|||7464|9|||1|583755|-1|4|3|44
503110827|BBBS of Greater Charlotte|Main Office|C|Active|2013-04-22|NaT|Followup|2014-04-22|2014-06-06|Complete|Done|4|3|4|2|3|3|3.17|4|4|1|4|4|4|3.5|-9.43|2|4|4|3|3|3|3.17|3|4|4|4|4|4|3.83|-17.23|4|4|4|4|4|4|4|4|0|4|4|4|||4|5|5|5|4.75||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Green|||46.8||1|1|1|1|M|Black||18|Yes|Mother|28262|One Parent: Female|$45,000 to $49,999|Y|No||Self|General Community||Match Support|M|White||31|28203|Masters Degree|Single|Consultant||0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503112489|31|0|1|503278385|1|0|1|500691045|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|584225|577768|4|3|45
500765381|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-26|2015-10-20|Followup|2014-02-26|2014-03-27|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|4|3|4|4|3.83|||||||||4|4|3|3.67||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green||Volunteer: Moved|79.7||1|1|1|1|M|Black||16|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||33|10019|Bachelors Degree|Single|Business: Marketing|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500739190|31|0|1|501579025|1|0|1|500342803|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|584239||4|3|45
502753873|BBBS of Greater Charlotte|Main Office|C|Active|2013-04-22|NaT|Followup|2014-04-22|2014-04-30|Complete|Done|4|4|4|2|4|4|3.67|3|3|3|3|4|4|3.33|10.21|2|4|4|2|2|4|3|3|2|3|3|2|3|2.67|12.36|4|4|4|4|4|4|4|4|0|5|4|5|5|4.75|3|3|3|3|3|58.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|3|3|3|3|22.33|2|3|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Green|||46.8||2|2|1|1|F|Hispanic||14|No|Mother|28262|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||43|28216|Masters Degree|Single|Finance: Accountant|28685|1|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502751081|3|0|2|503146044|31|0|2|500691867|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|584348|399995|4|3|45
500814240|BBBS of Greater Charlotte|Main Office|C|Active|2008-04-24|NaT|Followup|2014-04-24|2014-04-23|Complete|Done|4|4|4|4|4|4|4|||||||||1|4|4|4|1|4|3|||||||||4|4|4|4||||||1|4|3|4|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||106.7||1|1|1|1|M|Black||18|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||46|28215|Bachelors Degree|Single|Business: Mgt, Admin|28226|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500814509|31|0|1|500981509|31|0|1|500248568|2||500003586||2|1|500000294|500000294|-2|500000294|-2|34|2|||2238|7|||1|584617||4|3|45
503012569|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-24|2015-03-26|Followup|2014-04-24|2014-04-24|Complete|Done|3|4|4|1|3|4|3.17|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|23||2|3|1|2|F|American Indian or Alaska Native||13|No|Aunt|28027|Other Relative|Unknown||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||38|28027|Some College|Single|Arts, Entertainment, Sports|28025|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|504347632|6|0|2|502966672|1|0|2|500693960|2||-2||4|2||500014681, 500016374|-2||-2|0|4|||7496|10|1360|3|1|585216||4|3|45
500186702|BBBS of Greater Charlotte|Main Office|C|Completed|2004-04-28|2014-11-25|Followup|2014-04-28|2014-04-30|Complete|Done|3|4|4|3|4|3|3.5|||||||||4|4|4|3|3|4|3.67|||||||||4|4|4|4||||||3|5|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|1|2.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|126.9||1|2|1|2|F|Black||20|Yes|GrandMother|28208|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||57|28212|Some College|Married|Unknown||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|RTBM|277|60|598|500000170|500017732|500188150|31|0|2|500189528|31|0|2|500038225|2||500003586||4|1|500000294|500000294|-2|500015184|-1|0|10|||7462|13|||1|585342||4|3|45
502478428|BBBS of Greater Charlotte|Main Office|C|Active|2011-04-28|NaT|Followup|2014-04-28|2014-05-08|Complete|Done|4|4|4|3|4|4|3.83|4|4|1|4|4|4|3.5|9.43|4|4|3|4|4|4|3.83|4|2|4|2|4|4|3.33|15.02|4|4|4|4|4|4|4|4|0|3|4|5|5|4.25|4|5|5|5|4.75|-10.53|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|4|3.5|2|4|3|16.67|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||70.6||1|1|1|1|M|White||16|No|Mother|28277|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||54|28205|Some College|Separated|Self-Employed, Entrepreneur|28214|29|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502478875|1|0|1|502555822|1|0|1|500533009|2||-2||2|1|500005291|500005291|-2||-2|0|10|||7464|9|||1|585453|270021|4|3|45
501222138|BBBS of Greater Charlotte|Main Office|C|Completed|2010-04-30|2015-05-07|Followup|2014-04-30|2014-05-01|Complete|Done|2|1|2|2|3|4|2.33|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|60.2||2|2|2|3|F|Black||14|Yes|GrandMother|28227|Grandparents|Unknown||No||Self|General Community|Amachi|Enrollment|F|Black||53|28269|Some College|Married|Business: Sales|28227|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500012459|501222414|31|0|2|500189173|31|0|2|500447311|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|585472||4|3|45
503292494|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-24|2015-08-25|Followup|2014-04-24|2014-04-24|Complete|Done|4|2|4|1|4|4|3.17|||||||||1|4|4|1|4|4|3|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green||Child/Family: Moved|28||1|2|1|2|F|White||14|No|Mother|28083|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Some Other Race||44|28107|Bachelors Degree|Married|Finance|28025|0|0|ACN|Workplace Partner|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|277|60|598|500000170|500012459|503294318|1|0|2|503216525|41|0|2|500693959|2||-2||4|1|||-2|500007920, 500011315, 500011316|-1|0|4|||13581|3|||1|585512|523398|4|3|45
502197477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-02-10|2016-10-03|Followup|2014-02-10|2014-04-11|Declined|Late||||||||4|3|4|4|4|4|3.83|||||||||2|3|3|4|3|3|3||||||3|3|3|3|||||||5|3|3|5|4||||||||||4|4|4|3|3|4|4|3.71||||||4|4|3|3.67|||||4|4|4||||1|1||||4|4||Green|2010-2012 OJJDP JJI|Volunteer: Moved|67.7||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28202|Bachelors Degree|Single|Business: Sales|27560|1|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017732|502197915|31|0|1|502422929|1|0|1|500515536|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|0|4|||7464|9|||1|586507|241218|4|1|45
503452081|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-09|2014-10-20|Baseline|2013-04-29|2013-05-09|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|2|4|4|4|4|3.67|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green||Volunteer: Moved|17.4||1|1|1|1|M|White||15|No|Mother|28227|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||26|28269|Bachelors Degree|Single|Business: Engineer||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503453947|1|0|1|503371848|1|0|1|500694854|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|586808|-1|4|3|44
501525308|BBBS of Greater Charlotte|Main Office|C|Completed|2009-02-16|2015-06-18|Followup|2014-02-16|2014-02-27|Complete|Done|4|4|4|2|3|4|3.5|||||||||2|4|3|2|2|3|2.67|||||||||3|3|3|3||||||2|1|4|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|76||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28205|Some College|Married|Retail: Sales|28206|1|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|501525600|31|0|1|501536144|1|0|1|500335230|2||-2||4|1|||-2||-2|6854|8|||7464|9|||1|586891||4|3|45
501506214|BBBS of Greater Charlotte|Main Office|C|Completed|2009-03-28|2016-06-23|Followup|2014-03-28|2014-05-20|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|86.9||1|1|1|1|M|Black||19|No|Mother|28105|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||55|28173|||Unknown|28203|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501506506|31|0|1|501588885|31|0|1|500351462|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|586893||4|1|45
502249189|BBBS of Greater Charlotte|Main Office|C|Completed|2011-03-23|2016-09-22|Followup|2014-03-23|2014-04-10|Complete|Done|4|2|2|1|3|2|2.33|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|3|4|4|3.86||||||||||4|3|4|3.67||||||2|2|2|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|66||1|1|1|1|M|Black||13|No|Mother|28277|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||34|28262||Married|Finance|29715|6|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Enrollment|277|60|598|500000170|500017732|502249620|31|0|1|502485458|31|0|1|500523907|2||-2||4|1|||-2||-2|34|2|||7462|13|||1|586895||4|3|45
500186798|BBBS of Greater Charlotte|Main Office|C|Completed|2005-03-30|2015-10-20|Followup|2014-03-30|2014-03-31|Complete|Done|4|3|4|4|4|4|3.83|||||||||4|4|4|1|4|4|3.5|||||||||4|4|4|4||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||4|2|3|||||2|2||||4|4||||Green||Child/Family: Time constraints|126.7||1|2|1|2|F|Multi-Race (None of the above)||19|No|Father|28208|Two Parent|Unknown||No||Self|General Community||Match Support|F|White||45|28226|Bachelors Degree||Business: Human Resources||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|500187961|7|0|2|500189825|1|0|2|500038158|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|586897||4|3|45
500378354|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-01|NaT|Followup|2014-05-01|2014-05-07|Complete|Done|3|4|4|3|4|4|3.67|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||5|3|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||106.5||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$40,000 to $44,999||No|Big|Neighbor/Friend|General Community||Match Support|M|White||36|28270|Juris Doctorate (JD)|Married|Law: Lawyer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500378596|31|0|1|501181060|1|0|1|500264206|2||-2||2|1|||-2||-2|6854|8|||46|2|||1|586913||4|3|45
500361200|BBBS of Greater Charlotte|Main Office|C|Active|2006-03-21|NaT|Followup|2014-03-21|2014-03-21|Complete|Done|3|3|3|3|3|3|3|||||||||2|4|4|1|2|3|2.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Cabarrus County||131.8||2|2|1|1|F|White||17|No|Mother|28027|Two Parent|Unknown||No||Relative|General Community|Cabarrus County|Match Support|F|White||32|28115|Bachelors Degree|Single|Human Services: Social Worker||0|0|other|College Partner|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500361450|1|0|2|500368628|1|0|2|500085591|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|3|||7670|5|||1|587266||4|3|45
502885468|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-30|NaT|Followup|2014-04-30|2014-05-13|Complete|Done|3|4|4|2|4|4|3.5|4|4|4|4|1|4|3.5|0|4|4|4|2|2|4|3.33|4|4|4|1||3|||4|3|4|3.67|1|4|1|2|83.5|5|5|4|3|4.25|3|3|2|1|2.25|88.89|4|4|4|4|4|4|3|3.86|2|1|3|4|4|4|4|3.14|22.93|4|4|4|4|1|1|1|1|300|2|3|2.5|1|2|1.5|66.67|1|1|1|1|0|4|4|4|4|0|Green|||58.5||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Black||47|28227|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502886874|31|0|1|502954219|31|0|1|500610806|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|587355|425685|4|3|45
500740296|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-04|NaT|Followup|2014-05-04|2014-05-05|Complete|Done|3|4|3|4|3|4|3.5|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Yellow|||58.4||2|2|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Therapist/Counselor|General Community||Match Support|F|Asian||32|28216|Bachelors Degree|Single|Business: Mgt, Admin|28208|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500740560|31|0|2|502893901|4|0|2|500611525|2||-2||2|2|||-2||-2|0|5|||7464|9|||1|587499||4|3|45
502787401|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-30|2016-10-30|Followup|2014-04-30|2014-06-14|Complete|Done|3|2|3|2|3|3|2.67|4|3|4|4|1|3|3.17|-15.77|2|4|3|3|3|3|3|2|4|4|2|2|4|3|0|4|4|3|3.67|4|4|4|4|-8.25|2|3|3|3|2.75|4|4|4|4|4|-31.25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|3|3|3|3|3|4|4|3.67|-18.26|2|2|2|3|2|2.5|-20|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Lost contact with child/agency|42||1|1|1|1|F|Black||16|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||41|28105|High School Graduate|Divorced|Business: Mgt, Admin|28207|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502788587|31|0|2|503122442|1|0|2|500692539|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|587515|525811|4|3|45
502137546|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-29|2015-10-20|Followup|2014-04-29|2014-06-13|Declined|Done||||||||4|4|2|2|4|4|3.33|||||||||2|4|3|2|2|3|2.67||||||4|4|4|4|||||||4|3|5|4|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|4|3.5||||2|2|||||||Red|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|53.7||1|2|1|2|F|Black||16||Mother|28213|Other/Unknown|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28262|||Business: Mgt, Admin|75234|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502137975|31|0|2|501641708|31|0|2|500520728|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|587870|36419|4|1|45
502570188|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Followup|2014-04-30|2014-04-29|Complete|Done|4|3|3|3|4|4|3.5|4|3|3|2|4|4|3.33|5.11|3|4|4|4|2|4|3.5|2|4|4|2|3|4|3.17|10.41|4|4|4|4|4|4|4|4|0|4|3|3|4|3.5|5|5|5|4|4.75|-26.32|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|2|4|3|2|2|2|50|2|2|2|2|0|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|69.8||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||56|28226|Masters Degree|Married|Medical: Nurse|28217|34|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570642|31|0|2|502366830|1|0|2|500533448|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2|500004640|-2|0|4|||10326|3|||1|587871|271777|4|3|45
502570183|BBBS of Greater Charlotte|Main Office|C|Completed|2011-04-30|2017-02-23|Followup|2014-04-30|2014-04-29|Complete|Done|4|3|4|2|3|4|3.33|3|3|4|3|4|3|3.33|0|2|3|3|3|3|3|2.83|4|4|4|4|4|3|3.83|-26.11|4|4|3|3.67|4|4|3|3.67|0|4|4|3|3|3.5|3|3|4|3|3.25|7.69|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Agency: Challenges with program/partnership|69.8||1|1|1|1|F|Black||17|Yes|Mother|28206|Other/Unknown|Unknown||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||61|28134|Bachelors Degree|Married|Medical: Admin||33|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502570637|31|0|2|502570153|31|0|2|500534090|2||500004772||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|587878|273709|4|3|45
500783100|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-08-29|Followup|2014-04-30|2014-06-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|112||1|1|1|1|M|Black||16||Mother|28206|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||36|28203|||Retail: Sales|28226|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|500783368|31|0|1|500777047|1|0|1|500174449|2||-2||4|2|||-2||-2|0|10|||46|2|||1|587880||4|1|45
500271303|BBBS of Greater Charlotte|Main Office|C|Completed|2009-04-30|2015-08-03|Followup|2014-04-30|2014-05-21|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|1|2|4|2.83|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|75.1||2|2|1|1|F|Black||17|Yes|Mother|28227|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|White||31|28204|Bachelors Degree|Single|Business: Engineer|28269|0|2|TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|500271368|31|0|2|501291358|1|0|2|500354049|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||130|1|||1|588080||4|3|45
501390345|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-08|NaT|Followup|2014-05-08|2014-05-08|Complete|Done|3|4|4|2|3|3|3.17|||||||||2|4|3|1|2|3|2.5|||||||||4|3|3|3.33||||||3|3|3|3|3|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green|Amachi||58.3||2|2|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||35|28206|Bachelors Degree|Single|Business: Sales|28117|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501390617|31|0|1|502966998|1|0|1|500609269|2||-2||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|588756||4|3|45
502873189|BBBS of Greater Charlotte|Main Office|C|Completed|2012-03-21|2016-09-01|Followup|2014-03-21|2014-05-03|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|3|4|4|3|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|53.4||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||40|28216|Masters Degree|Single|Finance||6|0|Charlotte Cares|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502874592|31|0|2|502882530|31|0|2|500600322|2||-2||4|2|||-2||-2|0|4|||11246|6|||1|590511||4|3|45
502982301|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-22|2015-08-06|Baseline|2013-05-07|2013-05-21|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|3|4|4|4|3.33|||||||||4|4|4|4||||||2|4|4|4|3.5|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|2|3||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|26.5||1|1|2|2|M|Black||18|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||54|28262|Bachelors Degree|Married|Business||7|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|502983753|31|0|1|503442370|31|0|1|500695892|2||-2||4|1|||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|590573|-1|4|3|44
503452081|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-09|2014-10-20|Followup|2014-05-09|2014-05-16|Complete|Done|4|3|4|2|4|4|3.5|3|4|4|4|4|4|3.83|-8.62|4|1|4|3|4|4|3.33|4|2|4|4|4|4|3.67|-9.26|4|4|4|4|4|4|4|4|0|3|5|5|4|4.25|5|4|5|4|4.5|-5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|2|4|3|16.67|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|17.4||1|1|1|1|M|White||15|No|Mother|28227|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||26|28269|Bachelors Degree|Single|Business: Engineer||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503453947|1|0|1|503371848|1|0|1|500694854|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|591905|586808|4|3|45
500727291|BBBS of Greater Charlotte|Main Office|C|Completed|2007-05-17|2016-07-29|Followup|2014-05-17|2014-07-23|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|110.4||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|Black||46|28269|||Human Services: Non-Profit||0|0|BBBS National Site|Web Link|Big|General Community|VOL - Adjudicated, VOL - Cultural Comp, VOL - PreMatch|Match Support|277|60|598|500000170|500008321|500727558|31|0|1|500857838|31|0|1|500176403|2||-2||4|1|||-2|500007913, 500007920, 500011311|-2|0|10|||46|2|||1|592046||4|1|45
503216769|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-21|2017-02-28|Baseline|2013-05-10|2013-06-21|Complete|Done|4|4|4|4|4|3|3.83|||||||||2|3|3|3|2|3|2.67|||||||||4|3|3|3.33||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||3|4|3.5|||||2|2||||4|4||||Red||Child/Family: Moved|44.3||1|1|2|2|F|Black||18|No|Mother|28262|Two Parent|$75,000 to $99,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||25|28269|Bachelors Degree|Single|Education: Teacher|28210|0|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503218550|31|0|2|503344849|31|0|2|500698465|2||-2||4|3|||-2||-2|34|2|||46|2|||1|592542|-1|4|3|44
503469094|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-10|2016-04-29|Baseline|2013-05-10|2013-05-10|Complete|Done|3|3|2|1|2|3|2.33|||||||||2|3|3|3|2|4|2.83|||||||||4|2|2|2.67||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Green||Volunteer: Moved|35.6||1|1|1|1|F|Black||18|No|Mother|28216|Two Parent|Unknown|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||33|28269|Bachelors Degree|Single|Human Services: Non-Profit|28202|0|8|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|503470960|31|0|2|501717376|1|0|2|500696470|2||-2||4|1|||-2|500000294|-2|6854|8|||7464|9|||1|592583|-1|4|3|44
503469094|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-10|2016-04-29|Followup|2014-05-10|2014-07-03|Declined|Late||||||||3|3|2|1|2|3|2.33|||||||||2|3|3|3|2|4|2.83||||||4|2|2|2.67|||||||3|4|5|5|4.25||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||1|2|1.5||||2|2||||4|4||Green||Volunteer: Moved|35.6||1|1|1|1|F|Black||18|No|Mother|28216|Two Parent|Unknown|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||33|28269|Bachelors Degree|Single|Human Services: Non-Profit|28202|0|8|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|503470960|31|0|2|501717376|1|0|2|500696470|2||-2||4|1|||-2|500000294|-2|6854|8|||7464|9|||1|592599|592583|4|1|45
502904444|BBBS of Greater Charlotte|Main Office|C|Completed|2013-03-06|2014-10-22|Followup|2014-03-06|2014-04-03|Complete|Done|2|4|2|2|1|4|2.5|||||||||1|4|2|3|2|1|2.17|||||||||4|4|4|4||||||3|5|2|1|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child: Family structure changed|19.5||1|1|1|1|M|Black||12|Yes|Mother|28278|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|M|White||36|29715|Bachelors Degree|Single|Tech: Research/Design|28226|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502905855|31|0|1|502883475|1|0|1|500683493|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|593099||4|3|45
501247286|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-14|2016-11-08|Followup|2014-05-14|2014-05-14|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|101.8||1|1|1|1|M|White||15|No|Father|28025|One Parent: Male|Unknown||No||Self|General Community|Cabarrus County|Enrollment|M|White||49|27103|Masters Degree|Single|Education: Teacher|27282|0|0|Other|Service Organization|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|500341682|1|0|1|501247141|1|0|1|500264655|2||-2||4|1||500016374|-2|500016374|-2|0|10|||7452|6|||1|593183||4|3|45
503149009|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-13|2015-07-28|Baseline|2013-05-13|2013-06-13|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|2|3|2|3|2.67|||||||||4|4|4|4||||||2|4|4|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|25.5||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|$15,000 to $19,999|Y|Yes|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||37|28269|Masters Degree|Single|Business: Human Resources|28262|1|3|Recruitment Event|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|503150686|31|0|2|503199095|31|0|2|500696674|2||-2||4|3|||-2||-2|6855|8|||7460|12|||1|593541|-1|4|3|44
503209438|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-31|2014-04-30|Baseline|2013-05-13|2013-08-31|Complete|Done|3|4|4|3|3|4|3.5|||||||||4|3|3|4|3|4|3.5|||||||||4|4|3|3.67||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||1|1||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|8||1|1|1|1|F|Black||17||Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|F|White||29|28205|Masters Degree|Single|Finance: Accountant|28277|1|10|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503211213|31|0|2|503464333|1|0|2|500707202|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|593576|-1|4|3|44
502787404|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-26|NaT|Baseline|2013-05-14|2013-06-22|Complete|Done|3|2|1|1|4|4|2.5|||||||||1|4|4|2|2|4|2.83|||||||||3|4|2|3||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||2|4|4|3.33||||||1|1|1|||||1|1||||4|4||||Yellow|||44.6||1|1|1|1|M|Black||12|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Black||32|28262|Some College|Single|Business||0|5|United Way|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502788587|31|0|1|503485414|31|0|1|500701279|2||-2||2|2|||-2||-2|0|10|||16263|6|||1|593927|-1|4|3|44
501092911|BBBS of Greater Charlotte|Main Office|C|Completed|2008-05-01|2015-08-18|Followup|2014-05-01|2014-06-13|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|3|4|4|4|3.83|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5||||||||||4|4||||Red||Child: Graduated|87.6||1|1|1|1|M|Black||19||Mother|28226|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|M|White||37|28210|Some College|Single|Business: Mgt, Admin||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|501064244|31|0|1|501176101|1|0|1|500261235|2||-2||4|3|||-2||-2|0|4|||46|2|||1|594455||4|3|45
500185571|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-02|2015-07-14|Followup|2014-05-02|2014-06-16|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|110.4||1|1|1|1|M|Black||19||Mother|28215|Other/Unknown|Unknown||No|Other|Faith Organization|General Community||Match Support|M|Black||49|28213|Bachelors Degree|Married|Finance: Banking|28288|4|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187198|31|0|1|500188438|31|0|1|500089543|2||-2||4|3|||-2||-2|5635|9|||7464|9|||1|594456||4|1|45
502526965|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-03|NaT|Followup|2014-04-03|2014-05-15|Complete|Done|4|4|4|2|4|4|3.67|4|3|3|4|4|4|3.67|0|2|4|3|4|3|4|3.33|2|4|2|3|2|3|2.67|24.72|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|4|3|5|3.75|-20|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green|||59.4||1|1|1|1|M|Black||17|No|Mother|28278|Two Mothers|$50,000 to $59,999||No||Self|General Community||Match Support|M|White||32|28278|Bachelors Degree|Single|Medical|28208|3|5|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502527418|31|0|1|502881104|1|0|1|500606886|2||-2||2|1|||-2||-2|0|10|||17161|11|||1|594460|417778|4|3|45
502809446|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-12|2016-06-20|Followup|2014-04-12|2014-05-26|Complete|Done|2|2|3|1|4|3|2.5|4|4|4|4|3|4|3.83|-34.73|1|3|3|3|3|3|2.67|2|4|4|3|4|4|3.5|-23.71|3|3|3|3|3|4|4|3.67|-18.26|2|3|3|||4|3|5|4|4||4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|4|4|4|4|4|4|2|3.33|20.12|2|2|2|4|4|4|-50|2|2|1|1|100|4|4|4|4|0|Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|50.3||1|1|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Multi-race (Black & White)||33|28269|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502810724|31|0|2|502909383|36|0|2|500608444|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7462|13|||1|594462|421044|4|3|45
502710796|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-13|NaT|Followup|2014-04-13|2014-05-28|Complete|Done|4|4|4|2|4|4|3.67|4|1|2|1|4|4|2.67|37.45|2|4|4|4|4|4|3.67|1|1|3|1|1|4|1.83|100.55|4|4|4|4|3|4|3|3.33|20.12|4|4|4|4|4|3|4|4|2|3.25|23.08|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|4|3|3.5|1|4|2.5|40|2|2|2|2|0|4|4|4|4|0|Green|Project Big||59.1||1|1|1|1|M|Black||17|No|GrandMother|28208|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|Project Big|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502711683|31|0|1|502926804|1|0|1|500608316|2||500004641||2|1|500004640|500004640|-2||-2|6854|8|||7464|9|||1|594467|420876|4|3|45
502765606|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-03|2014-09-24|Followup|2014-04-03|2014-05-15|Complete|Done|2|2|4|2|4|4|3|4|1|2|2|2|4|2.5|20|2|3|3|2|2|3|2.5|3|2|3|2|2|2|2.33|7.3|3|3|3|3|4|4|4|4|-25|2|2|3|3|2.5|3|3|4|3|3.25|-23.08|4|4|4|4|4|4|4|4|3|4|3|4|2|4|4|3.43|16.62|4|4|4|4|3|4|4|3.67|8.99|2|2|2|3|2|2.5|-20|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Moved|29.7||1|1|1|1|F|Black||19|No|Mother|28105|One Parent: Female|$15,000 to $19,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28209|Some College|Single|Finance: Accountant|28232|0|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502766519|31|0|2|502842142|31|0|2|500607132|2||-2||4|3|||-2||-2|6854|8|||7462|13|||1|594470|418328|4|3|45
501212047|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-07|NaT|Followup|2014-05-07|2014-07-03|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||106.3||1|1|1|1|F|White||18|No|Father|28207|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||33|28226||Single|Human Services: Non-Profit|28205|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501212321|1|0|2|501242250|1|0|2|500264889|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|594471||4|1|45
501853851|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-10-20|Followup|2014-04-30|2014-06-14|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|Amachi|Child/Family: Moved|41.7||2|2|1|1|M|Black||13|Yes|Mother|28210|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||55|28105|Masters Degree|Married|Law: Lawyer||25|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|501854219|31|0|1|502922901|1|0|1|500608304|2||-2||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|594472||4|3|45
503292427|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-16|2015-09-15|Followup|2014-05-16|2014-05-19|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|4|3|4|3.5|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child/Family: Moved|28||1|2|1|2|M|White||13|No|GrandMother|28083|Grandparents|Unknown||No||School|General Community||Match Support|M|White||57|28027||Married|Business: Sales|28025|3|0|ACN|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500012459|503248831|1|0|1|503282196|1|0|1|500695385|2||-2||4|1|||-2||-2|0|4|||13581|3|||1|595612||4|3|45
502552445|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-12|NaT|Followup|2013-06-12|2013-06-24|Complete|Done|4|3|3|1|4|4|3.17|||||||||3|4|4|4|4|3|3.67|||||||||4|3|3|3.33||||||3|3|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||3|3||||Green|Project Big||69.1||1|1|1|1|F|Black||12|No|GrandMother|28208|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Project Big|Match Support|F|White||28|28209|Bachelors Degree|Single|Business: Sales|28277|0|9|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502552891|31|0|2|502545537|1|0|2|500539524|2||500004641||2|1|500004640|500004640|-2|500000294, 500004640|-2|0|4|||7464|9|||1|595996||4|3|45
501716720|BBBS of Greater Charlotte|Main Office|C|Completed|2010-03-02|2017-02-06|Followup|2014-03-02|2014-05-17|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Cabarrus County|Child/Family: Lost contact with volunteer/agency|83.2||1|1|1|1|M|Black||15|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||52|28075||Married|Medical: Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501716992|31|0|1|501878786|31|0|1|500435676|2||500016307||4|3|500016374|500016374|-2|500016374|-2|6854|8|||7464|9|||1|596020||4|0|45
502627468|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-17|2014-05-19|Followup|2014-05-17|2014-05-19|Declined|Done||||||||2|4|4|4|3|3|3.33|||||||||4|2|2|3|4|4|3.17||||||4|4|4|4|||||||4|4|5|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|4|3.5||||2|2||||4|4||Green||Child: Lost interest|12.1||1|1|1|1|M|Hispanic|Mexican|18|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||30|28036|Some College|Single|Business|28078|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500017777|502628116|3|10|1|503419352|1|0|1|500696276|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|596076|393156|4|1|45
502874566|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-24|2015-10-16|Followup|2014-05-24|2014-06-24|Complete|Done|3|3|1|2|3|3|2.5|3|1|3|1|3|4|2.5|0|2|3|4|2|2|3|2.67|2|3|4|2|3|4|3|-11|4|4|4|4|4|4|4|4|0|4|4|5|4|4.25|4|4|5|5|4.5|-5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|4|4|0|2|2|2|2|0|4|4||||Green||Volunteer: Moved|40.7||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|White||28|27235|Bachelors Degree||Business: Engineer||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502875969|3|10|2|502894480|1|0|2|500607372|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|596289|411252|4|3|45
503379566|BBBS of Greater Charlotte|Main Office|C|Active|2013-05-23|NaT|Baseline|2013-05-17|2013-05-23|Complete|Done|4|3|4|2|4|4|3.5|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Cabarrus County||45.8||1|1|1|1|M|Black||16||Mother|28027|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||51|28269|Bachelors Degree|Married|Business: Sales||6|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|503381423|31|0|1|503407492|1|0|1|500697331|2||500016307||2|1|500016374|500016374|-2|500016374|-2|34|2|||46|2|||1|596320|-1|4|3|44
502973981|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-02|2014-01-24|Baseline|2013-05-17|2013-07-02|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Feels incompatible with child/family|6.8||1|1|1|1|F|Black||18|No|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||55|28217|Masters Degree|Widowed|Education: Teacher|28208|0|6|BBBS National Site|Web Link|Big|General Community||RTBM|277|60|598|500000170|500011349|502875571|31|0|2|503484061|31|0|2|500701296|2||-2||4|1|||-2||-2|0|10|||46|2|||1|596332|-1|4|3|44
502073665|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-21|2016-02-04|Followup|2014-05-21|2014-05-21|Complete|Done|4|4|4|1|4|4|3.5|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||1|5|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Red||Child/Family: Moved|32.5||2|2|1|1|F|Black||13|No|Mother|29732|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|F|White||31|28226|Bachelors Degree|Single|Medical: Healthcare Worker|28211|0|3|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013781|502074089|31|0|2|503245956|1|0|2|500696434|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|598082||4|3|45
502278991|BBBS of Greater Charlotte|Main Office|C|Active|2010-12-03|NaT|Followup|2013-12-03|2014-01-16|Complete|Done|4|3|3|2|4|4|3.33|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|||75.4||1|1|1|1|F|Black||12|No|Mother|28213|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||40|28269|Bachelors Degree|Married|Tech: Management|28255|1|9|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502279417|31|0|2|502263116|31|0|2|500494784|2||-2||2|1|||-2|500000294|-2|6854|8|||6247|12|||1|598704||4|3|45
500724632|BBBS of Greater Charlotte|Main Office|C|Active|2007-03-07|NaT|Followup|2014-03-07|2014-05-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||120.3||1|1|1|1|F|Black||17||Mother|28213|One Parent: Female|Less than $10,000|Y|No||School|General Community||Match Support|F|Black||32|28214|Bachelors Degree|Married|Architect|28270|0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|500724899|31|0|2|500803551|31|0|2|500164708|2||-2||2|1|||-2||-2|0|4|||46|2|||1|598731||4|0|45
502982301|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-22|2015-08-06|Followup|2014-05-22|2014-07-23|Declined|Late||||||||4|4|4|4|4|4|4|||||||||2|3|3|4|4|4|3.33||||||4|4|4|4|||||||2|4|4|4|3.5||||||||||4|4|4|4|3|4|3|3.71||||||3|4|2|3|||||4|4|4||||2|2||||4|4||Green||Child/Family: Lost contact with volunteer/agency|26.5||1|1|2|2|M|Black||18|No|Mother|28215|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||54|28262|Bachelors Degree|Married|Business||7|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|502983753|31|0|1|503442370|31|0|1|500695892|2||-2||4|1|||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|599124|590573|4|1|45
501599416|BBBS of Greater Charlotte|Main Office|C|Active|2009-04-28|NaT|Followup|2014-04-28|2014-07-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||94.6||1|1|1|1|M|White||14|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||46|28078|Masters Degree|Single|Retail: Mgt|28207|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501599736|1|0|1|500188567|1|0|1|500357914|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|599567||4|0|45
503379566|BBBS of Greater Charlotte|Main Office|C|Active|2013-05-23|NaT|Followup|2014-05-23|2014-05-23|Complete|Done|4|4|4|4|4|4|4|4|3|4|2|4|4|3.5|14.29|4|4|4|3|3|4|3.67|3|4|4|3|4|4|3.67|0|4|4|4|4|4|4|4|4|0|4|4|4|2|3.5|4|4|4|5|4.25|-17.65|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|Cabarrus County||45.8||1|1|1|1|M|Black||16||Mother|28027|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||51|28269|Bachelors Degree|Married|Business: Sales||6|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|503381423|31|0|1|503407492|1|0|1|500697331|2||500016307||2|1|500016374|500016374|-2|500016374|-2|34|2|||46|2|||1|599778|596320|4|3|45
502549826|BBBS of Greater Charlotte|Main Office|C|Inactive|2013-05-28|NaT|Followup|2014-05-28|2014-05-28|Complete|Done|3|4|2|4|1|3|2.83|3|2|3|2|3|4|2.83|0|2|3|3|4|2|3|2.83|2|4|4|3|3|3|3.17|-10.73|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|3|3|3|3|3|8.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|3|3|3.33|3|4|4|3.67|-9.26|3|2|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Green|||45.6||4|4|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||38|28215|Bachelors Degree|Single|Business: Mgt, Admin|28210|11|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|2|503431300|31|0|2|500693780|2||-2||3|1||500014505, 500015184|-1||-2|0|4|||7464|9|||1|602066|285796|4|3|45
502966254|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-04|2015-03-18|Followup|2014-05-04|2014-06-16|Complete|Done|3|3|3|4|1|4|3|2|3|2|4|2|3|2.67|12.36|2|4|3|1|4|3|2.83|2|4|3|2|2|3|2.67|5.99|4|4|4|4|4|3|4|3.67|8.99|3|1|3|5|3|3|4|2|2|2.75|9.09|4|4|4|4|3|4|3|3.71|4|4|4|4|4|4|3|3.86|-3.89|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Lost contact with child/agency|34.4||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Self|General Community||Match Support|F|Black||48|28217|Bachelors Degree|Divorced|Medical: Admin|28232|11|5|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|500784955|31|0|2|502895517|31|0|2|500609631|2||-2||4|2|||-2||-2|0|10|||7438|1|||1|602849|423139|4|3|45
502829894|BBBS of Greater Charlotte|Main Office|C|Active|2013-05-31|NaT|Followup|2014-05-31|2014-06-11|Complete|Done|4|2|3|3|3|4|3.17|3|1|2|1|2|3|2|58.5|2|4|2|2|2|3|2.5|1|2|2|2|2|2|1.83|36.61|3|3|3|3|4|2|3|3|0|4|3|3|4|3.5|2|3|3|3|2.75|27.27|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Yellow|||45.5||2|2|1|1|F|Hispanic||14|No|Mother|28269|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Hispanic||41|28079|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|502831178|3|0|2|503443998|3|0|2|500696822|2||-2||2|2|||-2||-2|0|4|||7464|9|||1|606121|391151|4|3|45
502794252|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-31|2014-08-29|Followup|2014-05-31|2014-07-15|Complete|Done|3|2|3|3|3|3|2.83|||||||||2|4|2|2|3|3|2.67|||||||||4|3|2|3||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|2|2|||||2|2||||4|4||||Red||Volunteer: Time constraint|14.9||2|2|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|White||30|28202|Bachelors Degree|Single|Business|28203|1|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502129968|31|0|2|503351102|1|0|2|500696692|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|607209||4|3|45
503023832|BBBS of Greater Charlotte|Main Office|C|Active|2013-05-31|NaT|Followup|2014-05-31|2014-07-15|Complete|Done|3|4|3|2|4|3|3.17|4|2|2|2|2|2|2.33|36.05|1|4|3|2|3|3|2.67|2|3|3|2|2|3|2.5|6.8|4|4|4|4|3|3|3|3|33.33|3|3|3|3|3|3|3|3|3|3|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|1|1|100|4|4|4|4|0|Green|||45.5||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|White||33|28278|Bachelors Degree|Single|Arts, Entertainment, Sports|28269|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|503025372|31|0|1|503139766|1|0|1|500692957|2||-2||2|1|||-2||-2|0|10|||7671|13|||1|607367|484219|4|3|45
502845758|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-19|2015-09-16|Followup|2014-04-19|2014-06-03|Complete|Done|4|4|4|3|4|4|3.83|4|2|4|2|3|4|3.17|20.82|3|4|4|4|4|4|3.83|1|3|3|2|2|4|2.5|53.2|4|4|4|4|4|3|3|3.33|20.12|4|3|3|3|3.25|3|4|4|2|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|2|3|2.5|2|1|1.5|66.67|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|40.9||1|1|1|1|M|Black||15|No|Mother|28202|One Parent: Male|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28277||Single|Business||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502847118|31|0|1|502944923|1|0|1|500606912|2||-2||4|3|||-2||-2|34|2|||7464|9|||1|609309|417837|4|3|45
503405468|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-30|2015-10-01|Baseline|2013-06-05|2013-07-30|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|2|3|3|3|3|2.67|||||||||3|2|2|2.33||||||4|3|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|26.1||2|2|2|2|F|White||13|No|Father|28211|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||58|28277|High School Graduate|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503407325|1|0|2|502944301|1|0|2|500699540|2||-2||4|2||500014681|-2||-2|0|10|||7464|9|||1|611443|-1|4|3|44
503425373|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-24|2014-06-25|Baseline|2013-06-05|2013-06-24|Complete|Done|4|4|4|4|4|3|3.83|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Red||Child/Family: Moved|12||1|1|2|2|M|Multi-race (Black & White)||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||60|28269|Bachelors Degree|Married|Business: Sales|28079|9|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500013781|503427238|36|0|1|500967139|31|0|1|500699541|2||-2||4|3|||-2||-2|0|10|||4748|14|||1|611461|-1|4|3|44
502868969|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-18|NaT|Baseline|2013-06-05|2013-12-16|Complete|Done|2|4|4|4|3|4|3.5|||||||||2|4|4|1|3|3|2.83|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|4|3|||||2|2||||4|4||||Green|||38.9||1|1|1|1|F|Black||17|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||26|11237||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020753|502870370|31|0|2|503574667|1|0|2|500736904|2||-2||2|1|||-2|500000294|-2|0|10|||46|2|||1|611488|-1|4|3|44
500740295|BBBS of Greater Charlotte|Main Office|C|Completed|2007-06-12|2014-07-11|Followup|2014-06-12|2014-07-11|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Feels incompatible with child/family|85||1|1|1|1|M|Black||18||Mother|28216|One Parent: Female|$20,000 to $24,999||No||Therapist/Counselor|General Community||Match Support|M|White||55|28216|Bachelors Degree|Divorced|Tech: Engineer||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|500740560|31|0|1|500794907|1|0|1|500179696|2||-2||4|2|||-2||-2|0|5|||46|2|||1|611772||4|1|45
502402515|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-17|2015-12-28|Followup|2014-05-17|2014-05-16|Complete|Done|3|3|4|2|3|4|3.17|3|1|3|1|1|4|2.17|46.08|2|4|3|2|2|3|2.67|1|4|3|1|3|4|2.67|0|4|4|4|4|4|4|4|4|0|4|4|2|4|3.5|3|2|2|2|2.25|55.56|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|3|3.67|8.99|4|4|4|4|3|3.5|14.29|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|55.4||1|1|1|1|M|Black||16|No|Mother|28215|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28215||Single|Law: Police Officer||14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502402953|31|0|1|502537081|31|0|1|500535130|2||-2||4|1|500005291|500005291|-2||-2|34|2|||7464|9|||1|611844|276236|4|3|45
501722052|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-11|2015-01-30|Followup|2014-05-11|2014-07-26|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Time constraint|56.7||2|2|1|1|F|White||13|Yes|GrandMother|28083|Grandparents|Unknown||No||Self|General Community||Enrollment|F|White||40|28027||Single|Customer Service|28027|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501227925|1|0|2|502030533|1|0|2|500450450|2||-2||4|1|500000294||-2||-2|0|10|||7464|9|12|3|1|612074||4|0|45
503326540|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-24|2014-08-18|Baseline|2013-06-05|2013-06-24|Complete|Done|4|4|3|3|4|4|3.67|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|3|3|3|3.57||||||||||4|3|4|3.67||||||2|4|3|||||1|1||||4|4||||Red||Volunteer: Time constraint|13.8||2|2|1|1|F|Black||16|No|Mother|28215|Two Parent|$50,000 to $59,999||No||Self|General Community||Match Support|F|Black||30|28213|Some College|Single|Child/Day Care Worker||2|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|503328374|31|0|2|503459688|31|0|2|500699638|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|612165|-1|4|3|44
502813513|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-06|2016-05-04|Followup|2014-06-06|2014-06-09|Complete|Done|4|2|2|1|4|4|2.83|||||||||2|3|4|1|2|4|2.67|||||||||4|4|4|4||||||5|3|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green||Child: Lost interest|34.9||1|2|1|2|F|White||13|No|Non-Relative: Other|28164|Other/Unknown|Unknown||Yes||School|General Community||Match Support|F|White||39|28031|Bachelors Degree|Single|Arts, Entertainment, Sports|28031|5|6|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500020752|502814790|1|0|2|502915648|1|0|2|500697560|2||-2||4|1|||-2||-2|0|4|||7439|1|||1|612650||4|3|45
502287066|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-03|2014-09-04|Followup|2014-05-03|2014-06-26|Complete|Late|4|4|4|4|4|4|4|||||||||2|3|3|1|3|3|2.5|||||||||4|3|3|3.33||||||2|3|4|3|3|||||||4|4|4|4|2|3|1|3.14||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|40.1||2|2|1|1|M|Black||15||GrandMother|28227|One Parent: Female|Unknown|Y|Yes|AARTF|BBBS Board/Staff|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28215|Associate Degree|Married|Medical: Nurse||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502287498|31|0|1|502501212|1|0|1|500532817|2||-2||4|1|500005291|500005291|-2||-2|7294|13|||7464|9|||1|613758||4|3|45
502530227|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-04|2014-10-20|Followup|2014-05-04|2014-06-26|Declined|Late||||||||4|1|1|2|4|4|2.67|||||||||2|4|4|2|3|4|3.17||||||4|4|4|4|||||||5|5|4|5|4.75||||||||||4|4|4|3|4|3|4|3.71||||||3|4|3|3.33|||||2|4|3||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|41.6||1|1|1|1|F|Hispanic||15|No|Mother|28213|One Parent: Female|$10,000 to $14,999||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||30|28210|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502530676|3|0|2|502531485|3|0|2|500532078|2||-2||4|3|500005291|500005291|-2||-2|0|4|||7464|9|||1|613972|268895|4|1|45
502045254|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-08|2015-10-09|Followup|2014-06-08|2014-07-22|Complete|Done|2|4|4|4|4|4|3.67|2|4|4|4|3|4|3.5|4.86|3|4|4|3|2|4|3.33|2|4|3|2|2|3|2.67|24.72|4|4|4|4|4|4|4|4|0|2|5|3|3|3.25|2|4|3|3|3|8.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|2|3|33.33|4|4|4|3|3|3|33.33|2|2|1|1|100|4|4||||Yellow||Child: Graduated|64||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502171015|31|0|2|500454926|2||-2||4|2|||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1|613995|134736|4|3|45
502908460|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-07|2014-09-04|Followup|2014-06-07|2014-07-31|Declined|Late||||||||4|4|1|3|4|4|3.33|||||||||2|2|2|2|1|3|2||||||4|2|2|2.67|||||||1|5|3|3|3||||||||||4|4|4|4|3|4|2|3.57||||||4|4|3|3.67|||||4|1|2.5||||1|1||||4|4||Yellow||Volunteer: Lost contact with child/agency|26.9||1|1|1|1|F|Hispanic||18|No|Mother|28227|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||40|28079|Bachelors Degree|Single|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502909871|3|0|2|502938939|1|0|2|500616222|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|613999|434253|4|1|45
502552443|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-08|2014-12-30|Followup|2014-06-08|2014-06-13|Complete|Done|4|4|4|4|3|4|3.83|4|4|4|2|3|4|3.5|9.43|2|4|4|2|4|4|3.33|4|4|4|4|2|4|3.67|-9.26|4|4|4|4|4|4|4|4|0|3|4|5|4|4|5|4|4|5|4.5|-11.11|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|3|3.71|4.04|3|4|3|3.33|3|4|3|3.33|0|2|1|1.5|2|2|2|-25|2|2||||4|4||||Green|Project Big|Child: Graduated|42.7||1|1|1|1|F|Multi-race (Black & Hispanic)||20|No|GrandMother|28208|Grandparents|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28209|Bachelors Degree|Single|Medical|28209|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502552891|38|0|2|502471967|1|0|2|500537261|2||-2||4|1|500004640|500004640, 500005291|-2||-2|0|4|||7496|10|||1|614007|286064|4|3|45
502551092|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-20|2015-10-29|Followup|2014-05-20|2014-07-10|Complete|Late|3|4|4|4|1|3|3.17|3|3|4|1|4|4|3.17|0|3|4|3|4|2|4|3.33|2|4|3|1|2|4|2.67|24.72|4|4|4|4|4|4|4|4|0|4|4|5|5|4.5|3|4|5|3|3.75|20|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|2|3.71|4.04|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Yellow|Project Big, 2010-2012 OJJDP JJI|Volunteer: Feels incompatible with child/family|53.3||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||42|28210||Single|Business: Human Resources||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|502551545|31|0|2|502366844|1|0|2|500536172|2||-2||4|2|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||10326|3|460|3|1|614018|280274|4|3|45
502495501|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-20|NaT|Followup|2014-05-20|2014-07-17|Declined|Late||||||||3|1|4|2|2|2|2.33|||||||||2|3|3|1|2|3|2.33||||||4|4|4|4|||||||5|3|2|3|3.25||||||||||4|4|4|4|3|4|3|3.71||||||4|4|3|3.67|||||2|1|1.5||||1|1||||4|4||Green|2010-2012 OJJDP JJI||69.9||1|1|1|1|M|White||15|No|Mother|28226|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||55|28210|Bachelors Degree|Married|Finance|28203|1|6|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500018851|502495950|1|0|1|502508181|1|0|1|500531873|2||-2||2|1|500005291|500005291|-2|500005291|-2|0|10|||7464|9|||1|614023|268809|4|1|45
501919423|BBBS of Greater Charlotte|Main Office|C|Active|2010-03-24|NaT|Followup|2014-03-24|2014-02-10|Complete|Early|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|4|3|4|3.67|3|4|4|3|4|4|3.67|0|4|4|4|4|4|4|4|4|0|5|5|5|4|4.75|4|5|4|3|4|18.75|4|4|4|4|1|3|3|3.29|4|4|4|4|4|4|4|4|-17.75|4|4|4|4|4|4|3|3.67|8.99|4|3|3.5|4|3|3.5|0|2|2|1|1|100|4|4||||Green|Project Big||83.7||1|1|1|1|M|Multi-race (Black & Hispanic)||17|No|Mother|28214|One Parent: Female|Unknown||No|TV|Media|General Community|Project Big|Match Support|M|White||34|28164|Masters Degree||Finance|28210|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501919819|38|0|1|502034798|1|0|1|500442066|2||500004641||2|1|500004640|500004640|-2||-2|56|1|||7464|9|||1|614596|36152|4|3|45
502882034|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-13|NaT|Followup|2014-06-13|2014-06-11|Complete|Done|3|2|2|2|2|3|2.33|||||||||2|4|3|3|2|4|3|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green|||57.1||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||27|28208|Bachelors Degree|Single|Business: Mgt, Admin|28213|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501390617|31|0|2|502983700|31|0|2|500615277|2||-2||2|1||500000294|-2||-2|0|10|||7464|9|||1|614969||4|3|45
500186245|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-24|NaT|Followup|2014-05-24|2014-06-19|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|4|4|4|4|4|3.67|||||||||4|3|4|3.67||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|1|1.5|||||2|2||||4|4||||Green|Amachi||57.7||2|3|1|1|M|Black||16|Yes|Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|M|White||34|28203|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500187840|31|0|1|502989318|1|0|1|500614903|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|615130||4|3|45
503469072|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-24|2015-02-10|Baseline|2013-06-10|2013-06-24|Complete|Done|4|4|4|1|2|2|2.83|||||||||4|2|1|1|2|4|2.33|||||||||1|4|4|3||||||4|3|3|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|4|3.5|||||2|2||||4|4||||Red||Volunteer: Time constraint|19.6||2|2|1|1|M|White||13||GrandMother|28210|One Parent: Female|Unknown|Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||35|28217||Married|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503470938|1|0|1|503478672|1|0|1|500700143|2||-2||4|3||500014681|-2||-2|0|10|||7464|9|||1|615797|-1|4|3|44
502979757|BBBS of Greater Charlotte|Main Office|C|Completed|2013-02-28|2017-02-28|Followup|2014-02-28|2014-04-11|Complete|Done|4|3|3|2|4|4|3.33|||||||||2|4|4|4|3|4|3.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|2|3|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|48||1|1|1|1|M|Black||12|No|Mother|28211|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||31|28210|Bachelors Degree|Single|Business: Engineer||5|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502981210|31|0|1|503161988|1|0|1|500682191|2||-2||4|3|||-2||-2|0|10|||17161|11|||1|615823||4|3|45
503452382|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-28|2013-09-12|Baseline|2013-06-11|2013-06-28|Complete|Done|2|4|2|4|4|4|3.33|||||||||2|4|4|4|3|4|3.5|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|3|4|3.86||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|2.5||1|1|1|1|F|Multi-race (Black & White)||17|No|Mother|28269|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||25|28262|Some College|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500004169|503454248|36|0|2|503401641|1|0|2|500700156|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|616013|-1|4|3|44
501611456|BBBS of Greater Charlotte|Main Office|C|Active|2010-05-28|NaT|Followup|2014-05-28|2014-06-19|Complete|Done|3|2|4|1|4|4|3|||||||||2|3|3|4|2|4|3|||||||||4|4|4|4||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||81.6||1|1|1|1|M|Black||15|No|Mother|28262|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black|Other African|32|28262||Married|Law: Police Officer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501611776|31|0|1|501876475|31|31|1|500450969|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|616524||4|3|45
501142903|BBBS of Greater Charlotte|Main Office|C|Active|2008-06-05|NaT|Followup|2014-06-05|2014-06-17|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi||105.3||1|1|1|1|M|Black||14|Yes|GrandMother|28208|One Parent: Female|Less than $10,000||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|M|White||53|28204|Juris Doctorate (JD)|Married|Law: Lawyer|28244|16|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501143177|31|0|1|501236825|1|0|1|500268808|2||500003586||2|1|500000294|500000294|-2|500000294|-2|7294|13|||2238|7|||1|616587||4|3|45
502234905|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-05|2015-08-25|Followup|2013-12-05|2013-12-04|Complete|Done|4|2|4|1|4|4|3.17|||||||||2|3|4|2|4|3|3|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|44.6||3|3|1|1|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28083|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|M|White||36|28097|Masters Degree|Divorced|Finance|28026|7|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|502777258|38|0|1|502799047|1|0|1|500583119|2||-2||4|1|500000294|500000294, 500014681, 500016374|-2||-2|0|10|||7671|13|||1|616590||4|3|45
502763968|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2016-09-08|Followup|2014-04-30|2014-04-30|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Red||Volunteer: Moved|52.3||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Enrollment|M|White||38|28206|Bachelors Degree|Divorced|Business: Mgt, Admin|28164|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|502764880|31|0|1|502939016|1|0|1|500608284|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|617417||4|3|45
503149009|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-13|2015-07-28|Followup|2014-06-13|2014-07-28|Complete|Done|3|3|4|3|4|4|3.5|4|4|4|4|4|4|4|-12.5|3|4|4|3|3|4|3.5|2|4|2|3|2|3|2.67|31.09|4|4|4|4|4|4|4|4|0|2|4|4|3|3.25|2|4|4|3|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|2|3|4|2|3|0|2|2|2|2|0|4|4|4|4|0|Red||Child/Family: Lost contact with volunteer/agency|25.5||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|$15,000 to $19,999|Y|Yes|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||37|28269|Masters Degree|Single|Business: Human Resources|28262|1|3|Recruitment Event|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|503150686|31|0|2|503199095|31|0|2|500696674|2||-2||4|3|||-2||-2|6855|8|||7460|12|||1|617688|593541|4|3|45
502866475|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-23|NaT|Followup|2014-05-23|2014-07-17|Complete|Late|4|3|4|3|3|4|3.5|4|4|4|4|4|4|4|-12.5|2|4|3|2|3|3|2.83|3|4|4|2|4|4|3.5|-19.14|4|4|4|4|4|4|4|4|0|4|3|5|2|3.5|5|3|3|4|3.75|-6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|3|3.33|4|4|3|3.67|-9.26|4|4|4|4|4|4|0|2|2|1|1|100|4|4|4|4|0|Green|||57.8||1|1|1|1|M|Black||16|No|Mother|28270|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|M|White||29|28203|Bachelors Degree||Finance: Accountant||1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502867876|31|0|1|502961396|1|0|1|500614954|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|617925|418831|4|3|45
502566108|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-24|2014-09-08|Followup|2014-05-24|2014-07-17|Declined|Late||||||||3|2|4|1|3|4|2.83|||||||||2|3|3|2|2|3|2.5||||||4|3|4|3.67|||||||4|1|4|4|3.25||||||||||4|4|4|4|4|4|4|4||||||4|3|4|3.67|||||3|4|3.5||||1|1||||4|4||Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|39.5||1|1|1|1|F|Hispanic||17|No|Mother|28213|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||33|28209||Single|Student: College||0|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502566562|3|0|2|502562271|1|0|2|500535933|2||-2||4|1|500005291|500005291|-2|500005291|-2|0|4|||7464|9|||1|617958|279328|4|1|45
502320003|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2014-09-24|Followup|2014-04-30|2014-06-14|Complete|Done|4|2|3|2|3|3|2.83|4|2|4|4|3|4|3.5|-19.14|2|3|3|3|3|3|2.83|2|3|4|1|2|4|2.67|5.99|4|3|3|3.33|4|4|4|4|-16.75|2|3|3|2|2.5|4|3|5|4|4|-37.5|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|3|3|3|4|4|4|4|-25|2|3|2.5|4|1|2.5|0|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Moved|28.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||30|28216||Single|Tech: Research/Design||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502320438|31|0|2|502810883|31|0|2|500606071|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|618612|416362|4|3|45
502828137|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-06-29|Followup|2014-04-30|2014-06-14|Complete|Done|4|4|4|3|4|4|3.83|3|1|1|3|1|1|1.67|129.34|3|4|4|3|3|4|3.5|1|2|2|2|1|3|1.83|91.26|4|4|4|4|4|4|4|4|0|4|4||4||2|2|4|2|2.5||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|2|2|2|3|3|3|-33.33|2|2|2|2|0|4|4|4|4|0|Green||Child/Family: Moved|37.9||1|1|1|1|F|Multi-Race (None of the above)||16|No|Father|28214|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher|28078|0|8|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502829415|7|0|2|502446364|31|0|2|500607445|2||-2||4|1|||-2|500004640|-2|0|10|||7464|9|||1|618616|419338|4|3|45
500545470|BBBS of Greater Charlotte|Main Office|C|Completed|2007-04-30|2016-01-25|Followup|2014-04-30|2014-05-19|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|4|2|2|4|3|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|104.9||1|1|1|1|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||34|29708|Bachelors Degree|Single|Self-Employed, Entrepreneur|29708|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501750989|31|0|1|500815012|1|0|1|500173957|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|3|||2238|7|||1|618684||4|3|45
502879621|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-15|2014-11-13|Followup|2014-05-15|2014-07-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|30||1|1|2|2|F|Black||12|No|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|F|White||47|28078|Juris Doctorate (JD)|Single|Law: Lawyer|28203|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502881024|31|0|2|502295287|1|0|2|500603216|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|618689||4|1|45
501213488|BBBS of Greater Charlotte|Main Office|C|Active|2008-05-19|NaT|Followup|2014-05-19|2014-07-03|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||105.9||1|1|1|1|F|White||14|No|Father|28207|One Parent: Male|Unknown||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Finance: Banking|28255|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|501213764|1|0|2|501225276|1|0|2|500262655|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|619307||4|3|45
502319972|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-08-19|Followup|2014-04-30|2014-06-14|Complete|Done|4|3|2|3|3|3|3|4|4|4|1|4|4|3.5|-14.29|2|3|3|3|3|3|2.83|4|4|4|3|4|4|3.83|-26.11|4|4|4|4|4|4|4|4|0|2|2|3|3|2.5|4|4|3|4|3.75|-33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|||4|4|4|4||3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Moved|39.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Less than $10,000||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||32|28214|Bachelors Degree|Married|Self-Employed, Entrepreneur|29715|0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502320407|31|0|1|502911091|1|0|1|500607368|2||-2||4|2||500005291|-2||-2|6854|8|||7464|9|||1|619445|418896|4|3|45
502319984|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-30|2015-03-24|Followup|2014-04-30|2014-06-14|Complete|Done|3|2|2|2|2|2|2.17|3|3|4|4|4|4|3.67|-40.87|2|3|2|2|3|2|2.33|2|4|3|2|2|4|2.83|-17.67|3|2|2|2.33|4|4|4|4|-41.75|3|2|2|||3|3|4|4|3.5||4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|4|4|4|4|-25|2|3|2.5|4|3|3.5|-28.57|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Time constraint|34.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Bachelors Degree|Single|Finance|28216|3|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502320419|31|0|1|502290677|1|0|1|500607367|2||-2||4|3||500005291|-2||-2|6854|8|||17161|11|||1|619448|418895|4|3|45
502868925|BBBS of Greater Charlotte|Main Office|C|Completed|2012-04-25|2014-09-24|Followup|2014-04-25|2014-07-10|Expired|Late||||||||3|1|2|1|3|3|2.17|||||||||2|4|4|1|2|3|2.67||||||4|3|3|3.33|||||||3|4|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|3|2.5||||2|2||||4|4||Red||Child/Family: Lost contact with volunteer/agency|29||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||35|28262|Bachelors Degree|Divorced|Finance: Banking||2|6|Charlotte Cares|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502870324|31|0|2|502885744|31|0|2|500607510|2||-2||4|3|||-2||-2|0|4|||11246|6|||1|619450|419518|4|0|45
502183053|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-28|NaT|Followup|2014-06-28|2014-07-23|Complete|Done|2|2|3|1|1|2|1.83|3|1|2|1|1|2|1.67|9.58|3|4|3|1|1|3|2.5|4|2|4|2|3|4|3.17|-21.14|4|4|4|4|4|4|3|3.67|8.99|5|4|5|||4|4|4|4|4||4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|4|4|4|3|2|2.5|60|2|2|2|2|0|4|4|4|4|0|Green|||56.6||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||46|28134|Bachelors Degree|Married|Finance|28105|1|6|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|502183482|31|0|1|503073638|31|0|1|500621039|2||-2||2|1|||-2|500014681|-2|0|10|||4748|14|633|1|1|619801|414734|4|3|45
500934908|BBBS of Greater Charlotte|Main Office|C|Active|2010-06-18|NaT|Followup|2014-06-18|2014-06-20|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Green|Amachi||80.9||2|2|1|1|M|Black||16|Yes|Aunt|28216|One Parent: Female|Less than $10,000|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||34|20175|Bachelors Degree|Single|Business: Sales|28211|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|500935173|31|0|1|502107314|1|0|1|500456443|2||500003586||2|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|619858||4|3|45
500185778|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-17|2016-06-23|Followup|2014-06-17|2014-06-23|Complete|Done|3|1|3|1|2|3|2.17|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||1|4|2.5|||||1|1||||4|4||||Green||Child: Graduated|144.2||1|1|1|1|M|Black||18||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||42|27514||Married|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500187368|31|0|1|500188776|1|0|1|500036776|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|620556||4|3|45
503396873|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-09|2014-01-31|Baseline|2013-06-19|2013-08-08|Complete|Done|3|3|1|2|2|4|2.5|||||||||2|3|4|4|3|3|3.17|||||||||3|4|4|3.67||||||5|3|2|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green||Child: Lost interest|5.7||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||33|28202|Masters Degree|Single|Arts, Entertainment, Sports||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500008321|503398730|31|0|1|503381783|1|0|1|500701243|2||-2||4|1|||-2||-2|0|10|||46|2|||1|620785|-1|4|3|44
501143674|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-08|2016-08-05|Followup|2014-05-08|2014-06-20|Declined|Done||||||||3|4|3|3|1|3|2.83|||||||||2|2|2|3|2|4|2.5||||||2|3|3|2.67|||||||2|4|3|3|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|2|2||||2|2||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|50.9||3|3|1|1|F|Black||16||Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||28|28211|Bachelors Degree|Single|Human Services||2|0|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|277|60|598|500000170|500008321|501143948|31|0|2|502958999|1|0|2|500612879|2||500004641||4|2|||-2||-2|0|10|||132|8|||1|620865|17126|4|1|45
502583662|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-30|2014-06-19|Baseline|2013-06-20|2013-08-30|Complete|Done|4|1|2|1|3|4|2.5|||||||||1|3|4|2|3|2|2.5|||||||||3|4|4|3.67||||||3|4|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Red||Volunteer: Time constraint|9.6||3|3|1|1|F|Black||14|No|GrandMother|28215|Grandparents|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|F|Black||45|28204|Some College|Married|Finance: Banking|29715|4|0|Big For A Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500013781|502584168|31|0|2|503515217|31|0|2|500706497|2||-2||4|3|||-2||-2|0|4|||16422|8|||1|621292|-1|4|3|44
502583660|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-26|2014-06-26|Baseline|2013-06-20|2013-06-26|Complete|Done|4|1|4|1|4|4|3|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||4|3|5|3|3.75|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||4|1|2.5|||||2|2||||4|4||||Red||Volunteer: Time constraint|12||2|2|1|1|F|Black||14|No|GrandMother|28215|Grandparents|$30,000 to $34,999|Y|Yes||School|General Community||RTBM|F|White||32|28211|Bachelors Degree|Single|Business|28211|3|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502584168|31|0|2|503286709|1|0|2|500701403|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|621328|-1|4|3|44
501194563|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-20|NaT|Followup|2014-06-20|2014-06-19|Complete|Done|3|3|4|1|4|4|3.17|||||||||2|4|4|4|2|3|3.17|||||||||4|4|4|4||||||3|5|2|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||44.8||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$40,000 to $44,999||Yes||Self|General Community||Match Support|M|Black||30|28205|Bachelors Degree|Single|Self-Employed, Entrepreneur|28206|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501194837|31|0|1|503477116|31|0|1|500700141|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|621349||4|3|45
501224282|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-20|NaT|Followup|2014-06-20|2014-06-19|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||44.8||2|2|1|1|F|Black||15|Yes|Mother|28270|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||35|28205|Bachelors Degree|Married|Business: Mgt, Admin|28217|5|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501224558|31|0|2|503347558|1|0|2|500700583|2||-2||2|1|500000294|500000294|-2||-2|5635|9|||46|2|||1|621452||4|3|45
503024102|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-21|2014-09-30|Followup|2014-06-21|2014-07-16|Complete|Done|4|3|3|3|3|4|3.33|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|15.3||2|2|1|1|F|Black||13|No|Mother|28227|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|F|White||28|28212|Bachelors Degree|Single|Finance|28217|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501001116|31|0|2|503465770|1|0|2|500700716|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|621785||4|3|45
503216769|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-21|2017-02-28|Followup|2014-06-21|2014-08-04|Complete|Done|3|3|3|2|3|3|2.83|4|4|4|4|4|3|3.83|-26.11|3|3|3|3|2|3|2.83|2|3|3|3|2|3|2.67|5.99|4|3|3|3.33|4|3|3|3.33|0|4|4|4|4|4|3|4|4|4|3.75|6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|3|3|3|3|4|2|3|0|3|4|3.5|3|4|3.5|0|2|2|2|2|0|4|4|4|4|0|Red||Child/Family: Moved|44.3||1|1|2|2|F|Black||18|No|Mother|28262|Two Parent|$75,000 to $99,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||25|28269|Bachelors Degree|Single|Education: Teacher|28210|0|4|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503218550|31|0|2|503344849|31|0|2|500698465|2||-2||4|3|||-2||-2|34|2|||46|2|||1|621919|592542|4|3|45
502370669|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-22|NaT|Followup|2014-06-22|2014-06-23|Complete|Done|3|2|3|2|4|4|3|4|3|3|3|4|4|3.5|-14.29|4|1|3|2|2|4|2.67|3|4|4|3|3|3|3.33|-19.82|3|4|3|3.33|4|4|4|4|-16.75|5|4|5|4|4.5|2|4|4|4|3.5|28.57|3|4|4|3|4|4|3|3.57|4|4|4|4|4|4|4|4|-10.75|4|4|2|3.33|4|4|4|4|-16.75|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|||44.8||2|2|1|1|M|Black||18|No|Mother|28269|One Parent: Female|$40,000 to $44,999|Y|Yes||Self|General Community||Match Support|M|White||57|28277|Some College|Married|Business: Sales||28|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502371107|31|0|1|503472866|1|0|1|500700192|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|622104|362162|4|3|45
502513881|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-21|2014-09-22|Followup|2014-06-21|2014-08-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Lost contact with child/agency|27||2|2|3|3|F|Hispanic||14|No|Mother|28262|One Parent: Female|Unknown||No||School|General Community||Enrollment|F|Black||49|28213|Juris Doctorate (JD)|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502514330|3|0|2|502393006|31|0|2|500615307|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|622356||4|1|45
502527168|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-19|2016-08-29|Followup|2014-06-19|2014-07-30|Complete|Done|2|2|2|1|2|3|2|2|4|3|3|3|3|3|-33.33|2|4|4|3|2|3|3|2|4|3|2|3|3|2.83|6.01|4|3|3|3.33|4|4|4|4|-16.75|4|3|1|3|2.75|4|4|3|4|3.75|-26.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|3|4|3.67|3|3|4|3.33|10.21|4|4|4|4|3|3.5|14.29|2|2|2|2|0|4|4|4|4|0|Red||Child: Graduated|50.3||1|1|2|2|M|Hispanic|Mexican|19|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502527621|3|10|1|501646021|3|0|1|500618440|2||-2||4|3||500005291|-2||-2|2203|12|||7464|9|||1|622358|456875|4|3|45
502552438|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-02|2017-02-23|Followup|2014-06-02|2014-06-13|Complete|Done|4|3|3|3|4|4|3.5|4|3|4|1|3|4|3.17|10.41|3|4|3|3|3|4|3.33|4|4|4|2|4|3|3.5|-4.86|4|4|4|4|4|4|4|4|0|4|4|3|5|4|5|4|4|5|4.5|-11.11|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|4|4|3.67|-9.26|1|1|1|2|4|3|-66.67|2|2|2|2|0|4|4|4|4|0|Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|68.8||1|1|1|1|M|Black||16|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||36|28205|Masters Degree|Living w/ Significant Other|Journalist/Media|28202|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|502552891|31|0|1|502549491|1|0|1|500538826|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|10|||7464|9|||1|622362|292098|4|3|45
502552445|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-12|NaT|Followup|2014-06-12|2014-06-23|Complete|Done|3|1|4|1|4|4|2.83|||||||||2|4|3|2|3|3|2.83|||||||||4|4|4|4||||||5|4|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|2|3.33||||||1|2|1.5|||||2|2||||4|4||||Green|Project Big||69.1||1|1|1|1|F|Black||12|No|GrandMother|28208|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community|Project Big|Match Support|F|White||28|28209|Bachelors Degree|Single|Business: Sales|28277|0|9|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502552891|31|0|2|502545537|1|0|2|500539524|2||500004641||2|1|500004640|500004640|-2|500000294, 500004640|-2|0|4|||7464|9|||1|622364||4|3|45
503326540|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-24|2014-08-18|Followup|2014-06-24|2014-06-27|Complete|Done|3|4|4|2|3|4|3.33|4|4|3|3|4|4|3.67|-9.26|2|4|4|4|4|4|3.67|3|3|4|4|4|4|3.67|0|4|4|4|4|4|4|4|4|0|4|4|5|4|4.25|4|5|5|5|4.75|-10.53|4|4|4|4|4|3|3|3.71|4|4|4|4|3|3|3|3.57|3.92|4|4|4|4|4|3|4|3.67|8.99|3|2|2.5|2|4|3|-16.67|1|1|1|1|0|4|4|4|4|0|Red||Volunteer: Time constraint|13.8||2|2|1|1|F|Black||16|No|Mother|28215|Two Parent|$50,000 to $59,999||No||Self|General Community||Match Support|F|Black||30|28213|Some College|Single|Child/Day Care Worker||2|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|503328374|31|0|2|503459688|31|0|2|500699638|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|622444|612165|4|3|45
503469072|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-24|2015-02-10|Followup|2014-06-24|2014-07-19|Complete|Done|4|4|4|1|3|4|3.33|4|4|4|1|2|2|2.83|17.67|4|4|4|2|4|4|3.67|4|2|1|1|2|4|2.33|57.51|4|4|4|4|1|4|4|3|33.33|5|3|3|3|3.5|4|3|3|5|3.75|-6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|3|3.67|0|1|3|2|3|4|3.5|-42.86|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Time constraint|19.6||2|2|1|1|M|White||13||GrandMother|28210|One Parent: Female|Unknown|Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||35|28217||Married|Finance||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503470938|1|0|1|503478672|1|0|1|500700143|2||-2||4|3||500014681|-2||-2|0|10|||7464|9|||1|622471|615797|4|3|45
502549829|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-30|NaT|Followup|2014-06-30|2014-07-08|Complete|Done|4|4|4|4|3|4|3.83|3|1|2|1|2|2|1.83|109.29|2|4|3|2|2|3|2.67|2|3|2|2|2|2|2.17|23.04|4|4|4|4|3|2|2|2.33|71.67|2|2|3|3|2.5|3|2|2|3|2.5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|0|2|2|1|1|100|4|4||||Green|Amachi, Project Big, Project Big AND Amachi||68.5||1|1|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|Amachi, PERL 2014-2016, Project Big, Project Big AND Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Business: Engineer|30357|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|1|502594393|31|0|1|500541795|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901, 500014681|-1||-2|0|4|||7464|9|||1|622808|283404|4|3|45
502933371|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-13|NaT|Followup|2013-07-13|2013-07-12|Complete|Done|3|1|2|1|4|3|2.33|||||||||2|4|3|2|1|3|2.5|||||||||4|3|4|3.67||||||4|3|2|2|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||56.1||2|2|1|1|M|Black||12|No|Mother|28206|One Parent: Female|Less than $10,000|Y|Yes||Self|General Site||Match Support|M|White||37|28209|Bachelors Degree|Married|Unemployed|22202|9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|502934793|31|0|1|503080292|1|0|1|500623322|2||-2||2|1|||-1||-2|0|10|||7496|10|||1|622864||4|3|45
502700505|BBBS of Greater Charlotte|Main Office|C|Active|2012-06-27|NaT|Followup|2014-06-27|2014-08-01|Complete|Done|1|4|4|4|4|4|3.5|4|3|3|3|4|4|3.5|0|2|3|3|1|2|4|2.5|2|3|3|2|2|3|2.5|0|4|4|4|4|4|4|4|4|0|3|3|3|4|3.25|3|2|2|3|2.5|30|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3||||4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|||56.6||1|1|1|1|M|Black||17|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Black||41|28210|Bachelors Degree|Separated|Arts, Entertainment, Sports|28202|2|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502701350|31|0|1|503029324|31|0|1|500619505|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|622923|461562|4|3|45
501626226|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-30|2017-03-14|Followup|2014-06-30|2014-08-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|80.5||2|2|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||33|28203|High School Graduate|Single|Retail: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501622822|31|0|2|502036832|1|0|2|500457771|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|622925||4|1|45
502270499|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-25|NaT|Followup|2014-05-25|2014-07-09|Complete|Done|2|3|3|2|4|4|3|4|2|1|1|3|4|2.5|20|4|4|4|4|4|4|4|2|4|4|2|1|3|2.67|49.81|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3|4|3|4|3.5|42.86|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|4|3.5|4|4|4|-12.5|2|2|2|2|0|4|4||||Green|Amachi||69.7||2|2|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Unknown||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||34|28203|Masters Degree|Single|Business: Mgt, Admin|28273|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502231230|31|0|2|502510107|1|0|2|500536754|2||500003586||2|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|623412|218599|4|3|45
502393980|BBBS of Greater Charlotte|Main Office|C|Active|2012-05-25|NaT|Followup|2014-05-25|2014-07-09|Complete|Done|3|4|4|3|4|4|3.67|3|1|1|1|3|3|2|83.5|3|3|4|3|3|4|3.33|2|3|2|2|2|3|2.33|42.92|4|4|4|4|4|4|4|4|0|4|4|4|5|4.25|2|3|5|5|3.75|13.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|1|4|1|2|100|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Green|Amachi||57.7||2|2|1|1|F|Multi-race (Black & White)||16|Yes|Aunt|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28078|Associate Degree|Married|Tech: Support, Writing|28210|2|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|502394418|36|0|2|502928199|31|0|2|500613992|2||500003586||2|1|500000294|500005291|-2||-2|0|5|||7462|13|||1|623429|254548|4|3|45
502576641|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-25|NaT|Followup|2014-05-25|2014-07-09|Complete|Done|3|3|2|2|4|4|3|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|4|3.33||||||4|4|4|||||2|2||||4|4||||Green|||69.7||1|1|1|1|F|Black||13|No|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|White||41|28207|Masters Degree|Married|Business: Marketing|28202|2|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502577144|31|0|2|502537061|1|0|2|500535114|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|623435||4|3|45
502896719|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-01|2015-08-19|Followup|2014-06-01|2014-07-15|Complete|Done|3|3|3|2|4|4|3.17|4|1|2|1||4|||3|4|3|4|4|4|3.67|2|4|4|2|1|4|2.83|29.68|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|4|5|5|4.75|5.26|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|4|4|4|4|-8.25|4|4|4|2|3|2.5|60|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Moved|38.6||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|F|White||27|28269|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|502898127|31|0|2|502959645|1|0|2|500614239|2||-2||4|2|||-2||-2|0|10|||46|2|||1|623459|411397|4|3|45
501185592|BBBS of Greater Charlotte|Main Office|C|Completed|2008-06-23|2016-03-03|Followup|2014-06-23|2014-06-23|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|2|3|3|3|3|2.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green||Child: Family structure changed|92.3|Y|1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28227|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||45|28211||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|501185866|36|0|1|501255830|1|0|1|500270254|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|623588||4|3|45
502787404|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-26|NaT|Followup|2014-06-26|2014-08-08|Complete|Done|3|2|2|2|3|3|2.5|3|2|1|1|4|4|2.5|0|2|3|3|3|2|3|2.67|1|4|4|2|2|4|2.83|-5.65|3|2|3|2.67|3|4|2|3|-11|4|4|4|4|4|4|5|5|5|4.75|-15.79|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|2|2.67|2|4|4|3.33|-19.82|2|2|2|1|1|1|100|2|2|1|1|100|4|4|4|4|0|Yellow|||44.6||1|1|1|1|M|Black||12|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Black||32|28262|Some College|Single|Business||0|5|United Way|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|502788587|31|0|1|503485414|31|0|1|500701279|2||-2||2|2|||-2||-2|0|10|||16263|6|||1|623684|593927|4|3|45
501721762|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-26|NaT|Followup|2014-06-26|2014-06-26|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|3|3|3|3|2|2.67|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green|||44.6||3|3|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||39|28211||Single|Retail: Sales||0|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501722098|31|0|2|503471102|31|0|2|500700196|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|624015||4|3|45
502436198|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-27|NaT|Followup|2014-06-27|2014-06-27|Complete|Done|3|4|3|3|3|3|3.17|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|3|3||||||2|3|2.5|||||2|2||||4|4||||Green|||44.6||2|2|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28209|Masters Degree|Single|Medical|28207|0|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|502436641|31|0|2|503255826|1|0|2|500701262|2||-2||2|1|||-2||-2|34|2|||7496|10|||1|624148||4|3|45
500408135|BBBS of Greater Charlotte|Main Office|C|Completed|2006-05-25|2015-01-30|Followup|2014-05-25|2014-07-09|Complete|Done|3|3|4|3|4|3|3.33|||||||||2|4|3|4|4|3|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|104.2||1|1|4|4|F|Black||19|Yes|Mother|28083|One Parent: Female|Unknown||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500008321|500408385|31|0|2|500189709|31|0|2|500099932|2||500003586||4|1|500000294|500000294|-2|500000294, 500016374|-2|6854|8|||2230|7|||1|625683||4|3|45
502866443|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-14|2014-09-23|Followup|2014-06-14|2014-07-31|Declined|Late||||||||4|1|2|1|3|4|2.5|||||||||1|3|3|1|2|4|2.33||||||4|2|4|3.33|||||||5|3|5|4|4.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|1|2.5||||2|2||||4|4||Red||Volunteer: Lost contact with child/agency|27.3||1|1|1|1|F|Black||14|No|Mother|28262|One Parent: Female|$30,000 to $34,999|Y|No||Self|General Community||Match Support|F|Black||38|28212|Some College|Single|Business: Mgt, Admin|28270|7|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502867844|31|0|2|502920462|31|0|2|500613414|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|625685|432716|4|1|45
503465438|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-30|2014-10-31|Baseline|2013-07-01|2013-07-30|Complete|Done|3|1|4|4|1|3|2.67|||||||||1|3|4|1|1|4|2.33|||||||||4|4|3|3.67||||||1|5|5|||||||||4|4|3|4|4|4|4|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Red||Volunteer: Lost contact with child/agency|15||1|1|1|1|F|Black||13|No|Mother|28215|One Parent: Female|$35,000 to $39,999||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|Some Other Race||31|28262|Masters Degree|Single|Finance: Accountant|28262|2|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503467304|31|0|2|503422939|41|0|2|500702504|2||-2||4|3|||-2||-2|34|2|||7496|10|||1|626036|-1|4|3|44
500545328|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-02|2016-09-30|Followup|2014-07-02|2014-08-17|Complete|Late|4|2|2|3|3|3|2.83|||||||||2|4|3|3|1|3|2.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|99||3|3|1|1|F|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|F|Black||43|28208|Masters Degree|Single|Business: Sales|28078|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|2|501033808|31|0|2|500274449|2||-2||4|1|||-2||-2|0|10|||46|2|||1|626160||4|3|45
502223076|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-21|NaT|Followup|2013-10-21|2013-11-01|Complete|Done|3|1|2|1|4|3|2.33|||||||||2|4|3|1|3|3|2.67|||||||||4|2|2|2.67||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|||64.8||2|2|1|1|F|Black||12|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Mgt, Admin|28204|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|502223507|31|0|2|502694717|1|0|2|500560829|2||-2||2|1||500004640|-2||-2|0|10|||7464|9|||1|627083||4|3|45
503511553|BBBS of Greater Charlotte|Main Office|C|Active|2013-07-21|NaT|Baseline|2013-07-08|2013-07-19|Complete|Done|3|3|2|2|3|4|2.83|||||||||3|4|3|3|3|4|3.33|||||||||4|4|4|4||||||5|3|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||1|1||||4|4||||Green|||43.8||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|White||28|28273|Bachelors Degree||Business|28217|2|0|Elevation Church|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|503513424|31|0|1|503504991|1|0|1|500702866|2||-2||2|1|||-2||-2|0|10|||16414|7|||1|627225|-1|4|3|44
503484186|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-26|2016-03-08|Baseline|2013-07-08|2013-08-26|Complete|Done|3|3|4|3|3|3|3.17|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Child: Lost interest|30.4||1|1|1|1|M|White||16|No|Mother|28273|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|M|White||63|28226|Masters Degree|Widowed|Business: Marketing||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|503486052|1|0|1|503355490|1|0|1|500706097|2||-2||4|3|||-2||-2|0|10|||7671|13|1561|2|1|627226|-1|4|3|44
503492214|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2013-12-12|Baseline|2013-07-08|2013-10-24|Complete|Done|3|2|3|2|2|4|2.67|||||||||2|4|3|2|2|2|2.5|||||||||4|4|4|4||||||5|5|2|2|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||1|1|1|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|1.6||2|2|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Site|Amachi, mentor2.0, mentor2.0 2016|Match Support|F|White||50|28216|Bachelors Degree|Married|Business: Human Resources|28202|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503494082|31|0|2|503551073|1|0|2|500711788|2||-2||4|3||500000294, 500014505, 500016394|-1||-2|0|10|||7464|9|||1|627227|-1|4|3|44
503472839|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-26|2015-05-29|Baseline|2013-07-08|2013-07-25|Complete|Done|3|4|4|3|3|4|3.5|||||||||3|4|4|3|4|3|3.5|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|4|3|||||1|1||||4|4||||Green||Child/Family: Moved|22.1||1|1|1|1|F|Black||16|Yes|Mother|28214|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||25|28223|Some College|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503474705|31|0|2|503503841|31|0|2|500702872|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|627240|-1|4|3|44
502761742|BBBS of Greater Charlotte|Main Office|C|Active|2013-06-28|NaT|Followup|2014-06-28|2014-08-21|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Cabarrus County||44.6||1|1|2|2|M|Black||12|No|Mother|28083|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||60|28027|Bachelors Degree|Separated|Insurance|28262|24|0|Local Radio|Media|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502762654|31|0|1|503041890|1|0|1|500699565|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|10|||7437|1|||1|627518||4|1|45
502255156|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-24|NaT|Followup|2014-04-24|2014-04-24|Complete|Done|4|4|4|2|4|4|3.67|||||||||2|1|4|2|2|4|2.5|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi||58.7||2|2|1|1|F|Black||14|Yes|Relative: Other|28227|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||35|28277|Masters Degree|Single|Education: Admin||8|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|502255582|31|0|2|502946412|1|0|2|500608992|2||500003586||2|1|500000294|500000294|-2||-2|0|5|||7462|13|||1|627545||4|3|45
500186952|BBBS of Greater Charlotte|Main Office|C|Active|2004-07-15|NaT|Followup|2014-07-15|2014-07-31|Complete|Done|3|4|4|2|4|4|3.5|||||||||2|3|4|4|4|4|3.5|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi||152||1|1|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|White||73|28203||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|500188132|31|0|2|500189723|1|0|2|500037836|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|627638||4|3|45
502537477|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-12|2016-07-14|Followup|2014-05-12|2014-07-23|Declined|Late||||||||3|2|1|1|3|3|2.17|||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||3|5|4|4|4||||||||||4|4|4|4|3|4|3|3.71||||||2|3|2|2.33|||||2|4|3||||2|2||||4|4||Green|Project Big, 2010-2012 OJJDP JJI|Child: Graduated|62.1||1|1|3|4|F|Black||19||Mother|28208|Two Parent|$15,000 to $19,999||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||48|28214|Bachelors Degree|Single|Tech: Management|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Project Big|Enrollment|277|60|598|500000170|500017732|502537922|31|0|2|500189507|31|0|2|500535475|2||-2||4|1|500004640, 500005291|500004640, 500005291|-2|500000294, 500004640|-2|0|4|||2238|7|||1|628022|277756|4|1|45
502185074|BBBS of Greater Charlotte|Main Office|C|Completed|2011-05-12|2016-08-02|Followup|2014-05-12|2014-05-12|Complete|Done|2|2|1|1|2|2|1.67|1|2|1|4|1|1|1.67|0|3|3|3|2|2|2|2.5|3|1|3|1|1|1|1.67|49.7|4|4|4|4|4|4|4|4|0|2|3|3|3|2.75|3|2|4|5|3.5|-21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|2|3|2|2.33|42.92|2|4|3|2|2|2|50|2|2|2|2|0|4|4||||Green|2010-2012 OJJDP JJI|Child: Graduated|62.7||2|2|1|1|F|Black||18|No|GrandMother|28208|Grandparents|Unknown||Yes|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||68|28262|Bachelors Degree|Living w/ Significant Other|Business: Clerical||2|0|Relative|Relative|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017732|502185503|31|0|2|502490418|31|0|2|500533846|2||-2||4|1|500005291|500005291|-2|500000294, 500004640|-2|5635|9|||17161|11|||1|628023|159621|4|3|45
502566369|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-17|NaT|Followup|2014-07-17|2014-10-01|Expired|Late||||||||3|1|4|2|4|4|3|||||||||4|4|4|1|3|4|3.33||||||4|4|4|4|||||||3|5|4|5|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|4|4||||1|1||||4|4||Green|||56||2|2|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||49|28215|Bachelors Degree|Married|Business: Mgt, Admin|28277|13|0|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|502566823|31|0|2|503065299|1|0|2|500622859|2||-2||2|1|||-2||-2|0|10|||7439|1|||1|628059|275023|4|0|45
503328946|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-19|2016-08-09|Baseline|2013-07-10|2013-07-19|Complete|Done|3|1|1|2|2|4|2.17|||||||||1|3|4|1|2|3|2.33|||||||||4|3|4|3.67||||||3|5|3|5|4|||||||4|4|4|3||4|2|||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|36.7||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Enrollment|M|Black||26|28217|Bachelors Degree|Single|Business: Marketing|28217|4|0|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500013781|503330792|31|0|1|503371779|31|0|1|500703253|2||-2||4|1|||-2||-2|0|10|||7447|3|||1|628108|-1|4|3|44
500243491|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-10|NaT|Followup|2014-07-10|2014-08-05|Complete|Done|4|3|4|4|3|4|3.67|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||4|3|3|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||56.2||4|4|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||No||School|General Community|Amachi|Match Support|F|Black||47|28269|Bachelors Degree|Single|Law: Paralegal|28202|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188056|31|0|2|502919490|31|0|2|500619145|2||-2||2|1||500000294|-2||-2|0|4|||7464|9|||1|628115||4|3|45
501240369|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2014-10-09|Followup|2014-07-10|2014-07-07|Complete|Done|4|3|3|3|4|4|3.5|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||5|3|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|Amachi|Child: Graduated|75||1|1|1|1|M|Black||20|Yes|Mother|28214|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|M|White||43|28269|Masters Degree|Single|Business: Mgt, Admin|28202|3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|501240645|31|0|1|501240602|1|0|1|500272039|2||500003586||4|1|500000294|500000294|-2||-2|0|3|||131|1|||1|628118||4|3|45
502067798|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-09|NaT|Followup|2014-07-09|2014-08-14|Complete|Done|4|2|4|2|4|4|3.33|4|1|1|1|1|4|2|66.5|2|4|3|1|2|3|2.5|2|3|4|1|1|4|2.5|0|4|4|4|4|4|4|4|4|0|4|4|4|4|4|1|4|5|2|3|33.33|4|4|4|4|4|4|4|4|3|4|4|4|2|4|3|3.43|16.62|3|4|4|3.67|2|2|3|2.33|57.51|3|3|3|2|4|3|0|2|2|2|2|0|4|4||||Green|||80.2||1|1|1|1|M|Black||17|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|White||52|28270|Bachelors Degree|Married|Business: Mgt, Admin||4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|0|1|502062408|1|0|1|500459576|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|628164|154145|4|3|45
501755470|BBBS of Greater Charlotte|Main Office|C|Active|2010-06-30|NaT|Followup|2014-06-30|2014-07-31|Complete|Done|4|4|4|3|3|4|3.67|||||||||3|3|3|3|1|4|2.83|||||||||4|4|4|4||||||5|3|2|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green|||80.5||2|2|2|2|F|Black||13|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|501755813|31|0|2|502038804|31|0|2|500456645|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|628232||4|3|45
502980958|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-17|NaT|Followup|2014-07-17|2014-07-23|Complete|Done|3|3|4|3|3|4|3.33|3|2|3|3|3|3|2.83|17.67|3|3|3|3|3|3|3|3|3|3|3|3|3|3|0|4|4|4|4|4|3|4|3.67|8.99|3|5|5|3|4|4|4|3|3|3.5|14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|||56||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Sales|28273|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502982410|31|0|1|503008664|1|0|1|500620394|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|628653|463519|4|3|45
502034144|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-20|2014-12-04|Followup|2014-07-20|2014-07-16|Complete|Done|3|2|4|3|3|4|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|2|3.33||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|52.5||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||RTBM|M|Some Other Race||45|28210|Bachelors Degree|Married|Education: Teacher||0|0|CIS/Hidden Valley|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500018987|502034543|31|0|1|502212267|41|0|1|500460434|2||||4|1|||-2||-2|34|2|||11522|6|||1|628659||4|3|45
502933371|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-13|NaT|Followup|2014-07-13|2014-08-13|Complete|Done|3|2|1|1|1|1|1.5|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||5|5|5|||||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|||56.1||2|2|1|1|M|Black||12|No|Mother|28206|One Parent: Female|Less than $10,000|Y|Yes||Self|General Site||Match Support|M|White||37|28209|Bachelors Degree|Married|Unemployed|22202|9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|502934793|31|0|1|503080292|1|0|1|500623322|2||-2||2|1|||-1||-2|0|10|||7496|10|||1|628741||4|3|45
502549830|BBBS of Greater Charlotte|Main Office|C|Active|2011-06-30|NaT|Followup|2014-06-30|2014-07-08|Complete|Done|1|1|4|2|3|4|2.5|||||||||1|3|3|1|1|4|2.17|||||||||4|4|4|4||||||2|3|2|2|2.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||68.5||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Site|Amachi, Project Big, Project Big AND Amachi|Match Support|M|Black||25|28211||Single|Transport: Driver||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502550279|31|0|1|502462453|31|0|1|500538768|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-1||-2|0|4|||7464|9|||1|628961||4|3|45
501129794|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-14|2015-10-29|Followup|2014-06-14|2014-07-01|Complete|Done|3|3|4|2|2|4|3|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|52.5||1|2|1|2|M|Black||14||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|F|Black||45|28273|Masters Degree|Single|Tech: Research/Design||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500017777|501130068|31|0|1|500922570|31|0|2|500540937|2||-2||4|1|||-2||-2|0|4|||46|2|||1|628972||4|3|45
503459852|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-31|2014-09-22|Baseline|2013-07-15|2013-07-31|Complete|Done|3|2|2|1|2|3|2.17|||||||||2|3|3|1|2|3|2.33|||||||||4|4|3|3.67||||||5|2|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|13.7||1|1|1|1|F|Hispanic||16|No|Mother|28078|One Parent: Female|Less than $10,000||Yes|BBBS National Site|Web Link|General Community||RTBM|F|Hispanic||28|28031|Bachelors Degree||Business|28202|0|2|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|503461718|3|0|2|503208612|3|0|2|500703588|2||-2||4|1|||-2||-2|34|2|||46|2|||1|629135|-1|4|3|44
502570396|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-08|Followup|2014-06-30|2014-06-30|Complete|Done|4|4|4|4|4|4|4|3|4|4|4|4|4|3.83|4.44|2|4|3|4|2|4|3.17|4|4|3|4|2|3|3.33|-4.8|3|3|3|3|4|4|4|4|-25|1|3|2|3|2.25|3|5|3|3|3.5|-35.71|4|3|4|4|3|4|3|3.57|4|4|4|4|4|4|4|4|-10.75|3|4|2|3|4|4|4|4|-25|1|1|1|1|3|2|-50|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|51.3||1|1|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28215|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28078|Bachelors Degree|Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018987|502570850|38|0|2|502545897|31|0|2|500539251|2||-2||4|1|500005291|500005291|-2||-2|34|2|||46|2|||1|629215|296321|4|3|45
503047019|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-16|2014-02-27|Followup|2013-11-16|2014-01-31|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Time constraint|15.4||1|1|1|1|F|Hispanic||12|No|Mother|28211|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Hispanic||31|28210|Masters Degree|Single|Business||1|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500011746|503048667|3|0|2|503070946|3|0|2|500655762|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|629420||4|0|45
503255669|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-26|2016-05-25|Baseline|2013-07-16|2013-07-26|Complete|Done|1|4|4|4|4|4|3.5|||||||||3|4|4|3|2|4|3.33|||||||||4|3|3|3.33||||||4|4|3|5|4|||||||4|4|4|4|3|4|2|3.57||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Yellow||Child: Lost interest|34||1|1|2|3|M|Black||17|No|Mother|28216|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|M|Black||40|28202|Bachelors Degree|Single|Consultant|28281|4|5|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013781|503257474|31|0|1|500188812|31|0|1|500703771|2||-2||4|2|||-2|500000294|-2|0|10|||2238|7|||1|629607|-1|4|3|44
503230648|BBBS of Greater Charlotte|Main Office|C|Active|2013-07-17|NaT|Followup|2014-07-17|2014-09-04|Complete|Late|4|4|4|4|4|4|4|3|2|4|4|3|4|3.33|20.12|2|4|4|4|2|3|3.17|2|3|4|4|4|3|3.33|-4.8|4|4|4|4|4|4|4|4|0|3|5|4|5|4.25|3|5|4|5|4.25|0|3|4|4|4|3|4|3|3.57|4|4|4|4|4|4|4|4|-10.75|4|4|4|4|4|4|4|4|0|3|3|3|3|4|3.5|-14.29|1|1|2|2|-50|4|4|4|4|0|Green|||44||1|1|1|1|F|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|Black||39|28214|Bachelors Degree|Single|Govt||1|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502841119|31|0|2|503169561|31|0|2|500700323|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|629879|577620|4|3|45
502537469|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-17|2015-08-07|Followup|2014-07-17|2014-10-01|Expired|Late||||||||4|2|3|4|3|4|3.33|||||||||3|4|3|2|3|3|3||||||3|4|3|3.33|||||||3|3|4|5|3.75||||||||||4|4|4|4|4|4|4|4||||||3|4|4|3.67|||||2|4|3||||2|2||||4|4||Green||Volunteer: Feels incompatible with child/family|24.7||3|3|2|2|F|Black||16|No|Mother|28208|One Parent: Female|$15,000 to $19,999||No||School|General Site||Match Support|F|White||34|28078|Masters Degree|Single|Medical: Doctor, Provider|28001|0|2|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|502537922|31|0|2|503323641|1|0|2|500702088|2||-2||4|1|||-1|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|630063|274447|4|0|45
503187841|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-15|2016-06-20|Baseline|2013-07-19|2014-05-15|Complete|Done|3|4|3|3|1|3|2.83|||||||||1|4|4|4|3|4|3.33|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green||Child/Family: Moved|25.2||1|1|1|1|M|White||16||Mother|28277|One Parent: Female|$40,000 to $44,999|Y|No||Self|General Community||Match Support|M|White||60|28105|Bachelors Degree|Married|Tech: Research/Design|28277|4|0|Recruitment Event|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|503189585|1|0|1|503789478|1|0|1|500762532|2||-2||4|1|||-2||-2|0|10|||7460|12|||1|630563|-1|4|3|44
503328946|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-19|2016-08-09|Followup|2014-07-19|2014-08-04|Complete|Done|4|1|4|2|3|3|2.83|3|1|1|2|2|4|2.17|30.41|2|4|4|1|2|4|2.83|1|3|4|1|2|3|2.33|21.46|4|4|4|4|4|3|4|3.67|8.99|4|5|3|4|4|3|5|3|5|4|0|4|4|4|4|4|4|4|4|4|4|4|3||4|2|||4|4|4|4|3|4|4|3.67|8.99|2|3|2.5|3|2|2.5|0|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|36.7||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Enrollment|M|Black||26|28217|Bachelors Degree|Single|Business: Marketing|28217|4|0|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500013781|503330792|31|0|1|503371779|31|0|1|500703253|2||-2||4|1|||-2||-2|0|10|||7447|3|||1|630583|628108|4|3|45
501609876|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-13|2016-04-29|Followup|2014-07-13|2014-07-14|Complete|Done|1|4|4|4|2|2|2.83|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|4|3|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Child: Graduated|81.5||1|2|1|2|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|Black||38|28269|Masters Degree|Single|Medical: Nurse|28262|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|501610196|31|0|2|501425392|31|0|2|500373716|2||500004641||4|1|500004640|500004640|-2||-2|0|4|||7464|9|||1|630602||4|3|45
503360420|BBBS of Greater Charlotte|Main Office|C|Completed|2014-06-20|2016-03-04|Baseline|2013-07-19|2014-06-20|Complete|Done|2|4|2|2|3|2|2.5|||||||||4|4|4|3|3|4|3.67|||||||||4|4|2|3.33||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|3|3.33||||||2|4|3|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|20.5||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|$40,000 to $44,999||No||Self|General Community||Match Support|M|White||31|28262|Bachelors Degree|Single|Tech: Engineer|28262|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|503362265|31|0|1|503831013|1|0|1|500765209|2||-2||4|2|||-2||-2|0|10|||46|2|||1|630629|-1|4|3|44
503511553|BBBS of Greater Charlotte|Main Office|C|Active|2013-07-21|NaT|Followup|2014-07-21|2014-09-04|Complete|Done|4|3|3|2|4|4|3.33|3|3|2|2|3|4|2.83|17.67|2|4|3|4|4|4|3.5|3|4|3|3|3|4|3.33|5.11|4|3|2|3|4|4|4|4|-25|3|3|3|3|3|5|3|5|4|4.25|-29.41|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|3|3.67|4|4|4|4|-8.25|3|3|3|4|3|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Green|||43.8||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|White||28|28273|Bachelors Degree||Business|28217|2|0|Elevation Church|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|503513424|31|0|1|503504991|1|0|1|500702866|2||-2||2|1|||-2||-2|0|10|||16414|7|||1|630874|627225|4|3|45
500280148|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-13|NaT|Followup|2014-07-13|2014-07-19|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi||80.1||3|3|1|1|F|Black||16|Yes|Mother|28205|One Parent: Female|Unknown||No||Relative|General Community|Amachi|Match Support|F|Black||30|28216|Bachelors Degree|Single|Human Services: Non-Profit|28216|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500188151|31|0|2|502118494|31|0|2|500460767|2||500003586||2|2|500000294|500000294|-2||-2|0|3|||7464|9|||1|630877||4|3|45
500186682|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2015-07-22|Followup|2014-07-20|2014-07-17|Complete|Done|4|4|4|4|4|4|4|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|96.1||3|4|1|1|M|Black||20|Yes|Mother|28227|One Parent: Female|Less than $10,000|Y|No||Self|General Community|Amachi|Match Support|M|Black||57|28262||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|500887363|31|0|1|500184396|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|630878||4|3|45
501716763|BBBS of Greater Charlotte|Main Office|C|Completed|2010-05-07|2016-11-11|Followup|2014-05-07|2014-07-15|Complete|Late|1|1|1|1|2|2|1.33|1|1|1|1|1|1|1|33|1|2|2|1|1|4|1.83|2|1|2|2|3|2|2|-8.5|4|4|4|4|3|3|3|3|33.33|3|4|4|4|3.75|2|3|2|2|2.25|66.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|4|3.33|4|4|4|4|-16.75|2|2|2|4|4|4|-50|2|2|1|1|100|4|4||||Red||Child/Family: Lost contact with volunteer/agency|78.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Amachi, Cabarrus County|Match Support|F|Black||39|28269||Single|Self-Employed, Entrepreneur|28027|7|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501716992|31|0|2|502112513|31|0|2|500449029|2||-2||4|3||500000294, 500016374|-2|500016374|-2|6854|8|||7458|9|||1|630933|30228|4|3|45
501347097|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-30|2014-10-16|Followup|2014-07-30|2014-10-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Time constraint|74.5||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||35|28078|Bachelors Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500011349|501347376|31|0|2|501099568|1|0|2|500278256|2||-2||4|2|||-2||-2|0|10|||46|2|||1|630962||4|0|45
501513669|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-09|2015-02-04|Followup|2014-08-09|2014-10-24|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child/Family: Lost contact with volunteer/agency|29.9||1|2|2|3|F|White||18|No|Mother|28031|Other/Unknown|Unknown||No||School|General Community||Match Support|F|White||68|28036||Divorced|Business: Sales||5|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500011349|501513961|1|0|2|500824400|1|0|2|500626772|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|630967||4|0|45
500896588|BBBS of Greater Charlotte|Main Office|C|Completed|2007-07-20|2016-06-15|Followup|2014-07-20|2014-08-27|Complete|Done|4|3|3|4|3|4|3.5|||||||||2|4|4|3|3|4|3.33|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|2|3|2.67||||||2|3|2.5|||||2|2||||4|4||||Green||Child: Graduated|106.9||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28273|Two Parent|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||36|28269|Masters Degree|Married|Education|28205|6|6|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|500896858|3|15|2|500924445|1|0|2|500183434|2||-2||4|1|||-2||-2|0|10|||7671|13|||1|631127||4|3|45
501253965|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-11|2016-05-17|Followup|2014-06-11|2014-06-30|Complete|Done|4|4|4|4|3|4|3.83|||||||||2|3|4|2|2|3|2.67|||||||||4|4|4|4||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|47.2||3|3|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|Y|No||Self|General Community|Amachi|Enrollment|F|Black||34|28215|Some College|Single|Customer Service||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503287812|31|0|2|502985911|31|0|2|500613577|2||-2||4|1||500000294|-2||-2|0|10|||7464|9|||1|631149||4|3|45
501631140|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-17|2016-03-03|Followup|2014-06-17|2014-08-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|80.5||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Service: Hotel|28202|2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501631463|31|0|1|501628976|1|0|1|500367187|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|631151||4|1|45
500570756|BBBS of Greater Charlotte|Main Office|C|Active|2013-07-22|NaT|Followup|2014-07-22|2014-08-27|Complete|Done|2|3|3|3|3|4|3|||||||||2|4|2|2|3|3|2.67|||||||||4|3|3|3.33||||||2|3|5|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|4|3.5|||||2|2||||4|4||||Green|||43.8||4|5|2|2|F|Black||15||Aunt|28213|Two Parent|Unknown||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||24|28262|Some College|Single|Student: College|28216|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|500214349|31|0|2|502889143|31|0|2|500703847|2||-2||2|1||500004640, 500005291|-2||-2|0|4|||7464|9|||1|631156||4|3|45
501721761|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-25|2015-07-27|Followup|2014-06-25|2014-06-26|Complete|Done|3|2|4|2|4|4|3.17|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|2|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|37||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||RTBM|M|White||31|28210|Bachelors Degree|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501722098|31|0|1|503023854|1|0|1|500618753|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|631219||4|3|45
502506397|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-30|2016-11-01|Followup|2014-06-30|2014-07-31|Complete|Done|2|2|3|3|2|4|2.67|2|1|2|2|3|3|2.17|23.04|3|4|3|3|2|4|3.17|3|3|4|3|2|4|3.17|0|4|4|3|3.67|3|2|2|2.33|57.51|5|5|4|4|4.5|5|4|3|2|3.5|28.57|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|2|2|3|2.33|1|3|3|2.33|0|3|3|3|2|4|3|0|2|2|1|1|100|4|4|4|4|0|Yellow||Child: Severity of challenges|52.1||1|1|1|1|F|White||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||33|28277|Bachelors Degree|Single|Consultant|28202|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502506846|1|0|2|503039829|1|0|2|500619509|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|631222|407242|4|3|45
501157075|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-30|2016-01-21|Followup|2014-06-30|2014-07-31|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Yellow||Child: Lost interest|42.7||3|4|1|1|F|Black||17||Relative: Other|28206|Grandparents|Unknown||Yes||School|General Community|Amachi|Match Support|F|Black||37|28215|Masters Degree|Single|Human Services: Social Worker||2|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020752|501157349|31|0|2|502978065|31|0|2|500619009|2||-2||4|2||500000294|-2||-2|0|4|||7464|9|||1|631223||4|3|45
502207223|BBBS of Greater Charlotte|Main Office|C|Active|2013-07-23|NaT|Followup|2014-07-23|2014-07-22|Complete|Done|3|2|1|1|4|4|2.5|||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||2|3|2|2.33||||||1|4|2.5|||||2|2||||4|4||||Green|||43.8||2|2|1|1|F|Black||13|No|Mother|28216|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||38|28273|Bachelors Degree|Separated|Customer Service|28134|1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502207652|31|0|2|503251424|1|0|2|500703587|2||-2||2|1|||-2||-2|6854|8|||7464|9|||1|631313||4|3|45
501618024|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-26|2016-01-08|Followup|2014-07-26|2014-07-28|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|3|2|4|4|4|3.17|||||||||4|4|4|4||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|41.4||1|2|1|2|M|Hispanic||16||Mother|28031|Other/Unknown|Unknown||No||School|General Community||Match Support|M|White||65|28031|Some College|Married|Tech: Sales, Mktg|4241|5|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017777|501618344|3|0|1|501500078|1|0|1|500626248|2||-2||4|3|||-2||-2|0|4|||7462|13|||1|631678||4|3|45
502588461|BBBS of Greater Charlotte|Main Office|C|Completed|2011-07-22|2016-04-29|Followup|2014-07-22|2014-09-04|Declined|Done||||||||3|3|2|2|2|3|2.5|||||||||3|4|4|3|2|4|3.33||||||4|3|4|3.67|||||||4|5|4|5|4.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||4|4|4||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Child: Graduated|57.3||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||46|28278|Bachelors Degree|Separated|Transport: Pilot|28208|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|502588977|31|0|1|502636478|31|0|1|500546741|2||-2||4|3|500005291|500005291|-2||-2|6854|8|||46|2|||1|631679|319772|4|1|45
502530688|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-25|2016-05-20|Followup|2014-06-25|2014-07-15|Complete|Done|4|3|4|3|4|4|3.67|4|3|2|2|4|4|3.17|15.77|2|4|3|3|3|3|3|3|4|4|2|3|4|3.33|-9.91|4|3|3|3.33|4|4|4|4|-16.75|3|4|3|4|3.5|3|2|4|3|3|16.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|2|2|2|2|2|2|0|2|2|1|1|100|4|4|4|4|0|Yellow||Volunteer: Time constraint|46.8||2|2|3|3|M|Black||17||Mother|28210|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28277|Bachelors Degree|Married|Business||0|0|Michael Baisden|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502531141|31|0|1|502166996|31|0|1|500621632|2||-2||4|2||500005291|-2||-2|0|3|||11272|1|||1|631688|279295|4|3|45
503005868|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-24|2017-02-26|Followup|2014-07-24|2014-07-24|Complete|Done|3|1|3|1|1|3|2|2|2|2|1|2|3|2|0|2|1|3|1|2|3|2|2|2|3|2|2|3|2.33|-14.16|4|4|4|4|4|4|4|4|0|2|4|3|3|3|2|3|3|2|2.5|20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|3|3.67|4|4|4|4|-8.25|3|4|3.5|4|4|4|-12.5|2|2|2|2|0|4|4|4|4|0|Red||Child: Lost interest|55.1||1|1|1|1|M|Multi-race (Black & Hispanic)||15||Mother|28270|One Parent: Female|$25,000 to $29,999|Y|No||Therapist/Counselor|General Community||Match Support|M|White||51|28173|Bachelors Degree|Married|Consultant|28173|1|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020753|503007379|38|0|1|502935610|1|0|1|500623124|2||-2||4|3|||-2||-2|0|5|||7671|13|||1|631693|456253|4|3|45
502303088|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2016-08-29|Followup|2014-06-27|2014-08-12|Complete|Late|2|3|4|1|2|4|2.67|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Project Big|Volunteer: Time constraint|62.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community|Project Big|Enrollment|F|Black||33|28215|Bachelors Degree|Single|Human Services: Social Worker|28217|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500017777|502303520|31|0|2|502445797|31|0|2|500533193|2||-2||4|1|500004640|500004640|-2|500000294, 500004640|-2|6854|8|||7464|9|||1|631696||4|3|45
502813470|BBBS of Greater Charlotte|Main Office|C|Active|2013-07-24|NaT|Followup|2014-07-24|2014-07-24|Complete|Done|4|4|4|4|3|4|3.83|2|3|3|3|2|3|2.67|43.45|4|4|4|4|1|4|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||43.7||1|2|1|2|F|Black||14|No|Mother|28031|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|White||63|28031|Bachelors Degree|Married|Retired||0|0|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500020752|503507249|31|0|2|502889718|1|0|2|500701362|2||-2||2|1|||-2||-2|0|4|||7439|1|||1|631750|401353|4|3|45
503318447|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-27|2017-02-23|Baseline|2013-07-24|2013-09-27|Complete|Done|3|1|3|1|4|3|2.5|||||||||3|4|4|2|4|3|3.33|||||||||3|4|4|3.67||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Green||Agency: Challenges with program/partnership|40.9||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||47|28215|Bachelors Degree|Married|Finance: Banking|28269|13|6|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|503320281|31|0|1|503537303|31|0|1|500709889|2||-2||4|1|||-2||-2|0|10|||7458|9|||1|631862|-1|4|3|44
501402710|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-19|2015-06-17|Followup|2014-06-19|2014-08-04|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|71.9||1|1|1|1|M|Black||18|No|Mother|30058|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28215||Married|Consultant|28285|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501402995|31|0|1|501728845|1|0|1|500368860|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|632130||4|1|45
502578459|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-23|NaT|Followup|2014-07-23|2014-08-04|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Cabarrus County||55.8||1|1|1|1|M|Black||18|No|Mother|28025|One Parent: Female|$35,000 to $39,999||Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||48|28269|Some College|Married|Tech: Management|28204|10|0|AA Task Force|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502578962|31|0|1|502869485|31|0|1|500615803|2||500016307||2|2|500016374|500016374|-2|500016374|-2|6854|8|||9229|13|||1|632149|442607|4|3|45
502171910|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-30|2015-08-25|Followup|2014-07-30|2014-08-22|Complete|Done|3|3|4|2|3|4|3.17|3|1|2|2|2|3|2.17|46.08|2|4|4|2|2|4|3|2|3|3|4|2|4|3|0|4|4|4|4|4|4|4|4|0|3|4|3|5|3.75|4|3|4|3|3.5|7.14|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|4|4|4|4|-8.25|2|4|3|4|4|4|-25|2|2|2|2|0|4|4||||Red|Amachi|Volunteer: Time constraint|60.8||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28214|Some College|Married|Medical||3|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|502172339|31|0|1|502141964|31|0|1|500460627|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|5|||7464|9|||1|632162|156504|4|3|45
500186645|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-03|2016-01-06|Followup|2014-06-03|2014-07-21|Complete|Late|3|3|4|2|4|4|3.33|||||||||4|3|3|3|3|3|3.17|||||||||4|4|4|4||||||5|4|3|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|2|1|2||||||4|3|3.5|||||2|2||||4|4||||Green|Amachi|Child: Graduated|139.1||1|1|1|1|M|Black||18|Yes|Mother|28208|Other/Unknown|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28256|High School Graduate|Married|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500018987|500188043|31|0|1|500189545|31|0|2|500037636|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|632345||4|3|45
502569117|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-31|NaT|Followup|2014-05-31|2014-07-23|Declined|Late||||||||4|2|4|1|3|4|3|||||||||2|4|4|3|4|4|3.5||||||4|4|4|4|||||||5|4|5|3|4.25||||||||||4|4|4|4|4|4|3|3.86||||||4|3|2|3|||||2|2|2||||1|1||||4|4||Green|Amachi, 2010-2012 OJJDP JJI||69.5||1|1|1|1|F|Black||15|Yes|Mother|28206|One Parent: Female|$10,000 to $14,999|Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||40|28269|Masters Degree|Single|Tech: Engineer|77058|6|6|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500017732|502569571|31|0|2|502538689|31|0|2|500536957|2||500003586||2|1|500000294, 500005291|500005291|-2||-2|0|10|||17161|11|||1|632346|284793|4|1|45
503255669|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-26|2016-05-25|Followup|2014-07-26|2014-08-12|Complete|Done|2|4|4|4|4|4|3.67|1|4|4|4|4|4|3.5|4.86|3|4|4|1|3|4|3.17|3|4|4|3|2|4|3.33|-4.8|4|4|4|4|4|3|3|3.33|20.12|3|2|3|1|2.25|4|4|3|5|4|-43.75|4|4|4|4|3|4|4|3.86|4|4|4|4|3|4|2|3.57|8.12|3|4|4|3.67|3|4|4|3.67|0|2|3|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Yellow||Child: Lost interest|34||1|1|2|3|M|Black||17|No|Mother|28216|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|M|Black||40|28202|Bachelors Degree|Single|Consultant|28281|4|5|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500013781|503257474|31|0|1|500188812|31|0|1|500703771|2||-2||4|2|||-2|500000294|-2|0|10|||2238|7|||1|632546|629607|4|3|45
503472839|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-26|2015-05-29|Followup|2014-07-26|2014-09-09|Complete|Done|3|3|4|2|4|4|3.33|3|4|4|3|3|4|3.5|-4.86|3|4|4|4|4|4|3.83|3|4|4|3|4|3|3.5|9.43|4|4|4|4|4|4|4|4|0|3|3|4|4|3.5|3|4|4|5|4|-12.5|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|4|3.67|3|4|4|3.67|0|3|3|3|2|4|3|0|2|2|1|1|100|4|4|4|4|0|Green||Child/Family: Moved|22.1||1|1|1|1|F|Black||16|Yes|Mother|28214|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||25|28223|Some College|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503474705|31|0|2|503503841|31|0|2|500702872|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|632575|627240|4|3|45
503443162|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-20|2015-02-11|Baseline|2013-07-26|2013-08-20|Complete|Done|2|1|4|4|4|3|3|||||||||2|3|3|4|2|3|2.83|||||||||4|4|4|4||||||3|4|3|2|3|||||||4|4|4|3|4|3|2|3.43||||||||||4|3|4|3.67||||||1|1|1|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|17.7||1|1|2|2|M|Black||17|No|Mother|28262|One Parent: Female|$25,000 to $29,999||Yes||Relative|General Community||Match Support|M|Black||34|28213|Bachelors Degree|Single|Finance: Banking|28202|0|2|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503445028|31|0|1|500234684|31|0|1|500705816|2||-2||4|2|||-2||-2|0|3|||7458|9|||1|632640|-1|4|3|44
501314348|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-25|2015-07-31|Followup|2013-08-25|2013-10-18|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|59.2||1|1|1|1|M|Black||12|No|Mother|28210|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||45|28211|Masters Degree|Married|Finance: Banking||11|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|501314626|31|0|1|502205797|1|0|1|500460633|2||-2||4|3|||-2||-2|0|10|||2230|7|||1|632872||4|1|45
501645192|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-21|2016-08-19|Followup|2014-07-21|2014-07-22|Complete|Done|3|4|4|2|4|4|3.5|||||||||4|4|4|2|2|4|3.33|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red||Child: Graduated|85||1|1|2|2|M|Hispanic||19|No|Mother|28025|One Parent: Female|Unknown||Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500020753|501645515|3|0|1|501519306|1|0|1|500374818|2||-2||4|3||500016374|-2|500016374|-2|0|10|||7464|9|||1|633087||4|3|45
503405468|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-30|2015-10-01|Followup|2014-07-30|2014-07-29|Complete|Done|4|4|4|2|1|4|3.17|3|4|4|2|4|4|3.5|-9.43|2|4|3|1|2|3|2.5|2|2|3|3|3|3|2.67|-6.37|4|4|4|4|3|2|2|2.33|71.67|4|3|3|5|3.75|4|3|5|4|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|3|3|3|4|4|4|-25|1|1|2|2|-50|4|4|4|4|0|Yellow||Volunteer: Time constraint|26.1||2|2|2|2|F|White||13|No|Father|28211|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||58|28277|High School Graduate|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503407325|1|0|2|502944301|1|0|2|500699540|2||-2||4|2||500014681|-2||-2|0|10|||7464|9|||1|633337|611443|4|3|45
503465438|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-30|2014-10-31|Followup|2014-07-30|2014-09-12|Complete|Done|3|2|3|2|4|4|3|3|1|4|4|1|3|2.67|12.36|2|3|3|3|3|3|2.83|1|3|4|1|1|4|2.33|21.46|3|3|3|3|4|4|3|3.67|-18.26|2|3|3|3|2.75|1|5|5||||4|4|4|4|4|4|3|3.86|4|4|3|4|4|4|4|3.86|0|3|3|3|3|4|4|3|3.67|-18.26|3|3|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|15||1|1|1|1|F|Black||13|No|Mother|28215|One Parent: Female|$35,000 to $39,999||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|Some Other Race||31|28262|Masters Degree|Single|Finance: Accountant|28262|2|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503467304|31|0|2|503422939|41|0|2|500702504|2||-2||4|3|||-2||-2|34|2|||7496|10|||1|633529|626036|4|3|45
502142541|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-18|2015-07-23|Followup|2014-06-18|2014-07-29|Complete|Done|3|4|4|4|4|4|3.83|3|4|4|3|4|4|3.67|4.36|2|4|3|3|2|3|2.83|3|3|3|3|3|3|3|-5.67|4|4|4|4|4|4|4|4|0|1|4|5|3|3.25|4|4|5|3|4|-18.75|4|4|4|4|3|4|4|3.86|4|4|4|4|3|4|3|3.71|4.04|4|4|4|4|4|4|4|4|0|1|1|1|2|2|2|-50|2|2|2|2|0|4|4||||Green||Child: Graduated|61.1||1|1|2|2|F|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|502142970|31|0|2|501905673|31|0|2|500455759|2||-2||4|1|||-2||-2|0|4|||7496|10|||1|633997|141478|4|3|45
501872144|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-30|NaT|Followup|2014-07-30|2014-08-26|Complete|Done|4|4|4|3|3|4|3.67|4|4|3|1|3|3|3|22.33|4|4|3|3|2|||2|3|2|1|2|2|2||4|4|4|4|2|3|2|2.33|71.67|3|5|4|4|4|2|2|1|2|1.75|128.57|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|3|3.67|8.99|4|2|3|1|1|1|200|2|2|2|2|0|4|4||||Green|||79.5||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown|Y|Yes||Relative|General Community||Match Support|M|White||35|28205|Masters Degree|Married|Tech: Engineer|28115|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501872517|31|31|1|502063676|1|0|1|500460156|2||-2||2|1|||-2||-2|0|3|||46|2|||1|637195|155585|4|3|45
503021552|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-19|2015-10-22|Followup|2014-06-19|2014-06-24|Complete|Done|2|1|4|1|4|4|2.67|3|1|1|4|3|4|2.67|0|4|4|4|4|4|4|4|2|4|4|4|2|4|3.33|20.12|4|4|4|4|4|4|4|4|0|5|4|5|5|4.75|3|4|3|4|3.5|35.71|4|4|4|4|4|4|4|4|4|4|4|4|4|4||||3|3|4|3.33|4|4|3|3.67|-9.26|2|3|2.5|2|3|2.5|0|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Moved|40.1||1|1|1|1|F|Black||14|No|Mother|28270|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Multi-Race (None of the above)||28|28215|Some College|Single|Insurance||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503023091|31|0|2|502951522|7|0|2|500618601|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|637483|457665|4|3|45
503448711|BBBS of Greater Charlotte|Main Office|C|Completed|2014-02-26|2015-11-19|Baseline|2013-08-02|2014-02-20|Complete|Done|3|3|4|3|3|3|3.17|||||||||2|4|3|4|3|3|3.17|||||||||4|4|4|4||||||2|3|2|2|2.25|||||||4|4|4|4|3|4|4|3.86||||||||||2|4|4|3.33||||||2|1|1.5|||||1|1||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|20.7||1|1|1|1|M|Black||17|No|Mother|28226|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|White||34|28210|Masters Degree|Married|Real Estate: Realtor|28202|2|3|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503450577|31|0|1|503576769|1|0|1|500742906|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|637485|-1|4|3|44
502997224|BBBS of Greater Charlotte|Main Office|C|Completed|2012-05-21|2015-04-13|Followup|2014-05-21|2014-06-20|Complete|Done|3|4|4|2|3|4|3.33|||||||||2|4|3|3|2|4|3|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||1|4|1|2||||||2|3|2.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|34.7||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Black||32|28210|Bachelors Degree|Married|Business: Human Resources|28269|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|502998689|31|0|2|502939526|31|0|2|500613729|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|637803||4|3|45
502222545|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-03|2017-01-24|Followup|2014-08-03|2014-08-13|Complete|Done|3|3|4|4|2|2|3|||||||||1|3|4|2|3|3|2.67|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|77.7||1|1|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||School|General Community||Enrollment|F|White||37|28208|Masters Degree|Single|Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502222979|31|0|2|502196116|1|0|2|500462566|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|637822||4|3|45
502183217|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-05|NaT|Followup|2014-08-05|2014-08-05|Complete|Done|4|2|3|2|4|4|3.17|||||||||4|4|4|2|3|4|3.5|||||||||4|4|4|4||||||5|3|5|5|4.5|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green|Amachi||79.3||1|1|2|2|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|Black||50|28078|||Service: Restaurant|28082|0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502183646|31|0|1|501733851|31|0|1|500462588|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7464|9|||1|637825||4|3|45
500186956|BBBS of Greater Charlotte|Main Office|C|Completed|2004-06-21|2015-03-04|Followup|2014-06-21|2014-08-05|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Child: Graduated|128.4||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||54|28203|Bachelors Degree|Married|Law: Lawyer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|500189727|1|0|1|500037841|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|638010||4|1|45
503452963|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-22|2015-01-21|Baseline|2013-08-06|2013-08-22|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|4|2|3|3|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|17||1|1|1|1|M|Black||14|No|Mother|28211|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|M|Black||41|28216|Bachelors Degree|Single|Customer Service|28262|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|503430105|31|0|1|503489818|31|0|1|500705904|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|638157|-1|4|3|44
500826603|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-06|2015-02-11|Followup|2014-08-06|2014-10-21|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|18.2||3|3|2|2|F|Black||16|No|Mother|28226|Two Parent|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|F|Black||34|28215|Some College|Single|Finance: Banking|28270|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|500826861|31|0|2|502672644|31|0|2|500703783|2||-2||4|2|||-2||-2|0|5|||7464|9|||1|638169||4|0|45
502090492|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-13|2013-09-26|Followup|2013-09-13|2013-09-04|Blank|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Feels incompatible with child/family|12.4||1|1|1|1|M|Black||12|No|Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||44|28213|Associate Degree|Single|Laborer|28216|4|6|Local TV|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502090916|31|0|1|503088662|31|0|1|500631918|2||-2||4|3|||-2||-2|0|10|||7438|1|||1|638329||4|3|45
503014417|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-26|2016-08-17|Baseline|2013-08-07|2013-08-24|Complete|Done|4|1|4|2|4|4|3.17|||||||||2|4|4|4|2|3|3.17|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|3|3.67||||||2|1|1.5|||||2|2||||4|4||||Green||Child: Lost interest|35.7||1|1|1|1|F|Black||17|No|Mother|28203|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||29|28110|Masters Degree|Single|Education: Teacher||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|503015947|31|0|2|503518076|1|0|2|500706096|2||-2||4|1|||-2||-2|0|10|||46|2|||1|638535|-1|4|3|44
501726201|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-08|2015-01-30|Followup|2014-07-08|2014-08-22|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Moved|66.8||1|1|1|1|F|Black||17|Yes|Mother|28212|One Parent: Female|Unknown||Yes|YeaGod|Faith Organization|General Community|Amachi|Match Support|F|Black||51|28262|PHD|Married|Real Estate: Realtor||0|0|Weeping Willow|Faith Organization|Big|General Community||Enrollment|277|60|598|500000170|500008321|501726541|31|0|2|501734664|31|0|2|500371036|2||-2||4|3|500000294|500000294|-2||-2|5634|9|||9218|7|||1|638639||4|1|45
501488919|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-09|2015-08-25|Followup|2014-08-09|2014-08-12|Complete|Done|4|2|4|1|4|4|3.17|||||||||2|4|3|2|2|3|2.67|||||||||4|4|3|3.67||||||4|5|5|5|4.75|||||||4|3|3|3|4|3|3|3.29||||||||||3|3|3|3||||||2|4|3|||||2|2||||4|4||||Yellow||Child: Lost interest|36.5||1|2|1|2|F|Black||17||Mother|28031|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||36|28205|Bachelors Degree|Single|Business: Mgt, Admin|28036|0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501489205|31|0|2|501392684|31|0|2|500626771|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|638759||4|3|45
502045258|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-25|2016-08-29|Followup|2014-06-25|2014-08-11|Declined|Late||||||||4|2|4|1|4|4|3.17|||||||||4|4|4|4|4|4|4||||||4|4|4|4|||||||5|5|5|5|5||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||4|3|3.5||||2|2|||||||Green||Volunteer: Lost contact with child/agency|74.2||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||33|28262|Bachelors Degree|Single|Medical: Nurse|28262|4|9|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017777|502045664|31|0|2|502190790|31|0|2|500457916|2||-2||4|1|||-2||-2|0|10|||6247|12|||1|638785|148107|4|1|45
502589865|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-30|2015-10-29|Followup|2014-06-30|2014-07-02|Complete|Done|4|3|3|1|3|4|3|1|4|2|3|1|1|2|50|3|4|4|4|4|4|3.83|3|1|3|4|4|4|3.17|20.82|4|4|4|4|4|4|4|4|0|3|4|5|4|4|5|5|5|5|5|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|3|3.33|20.12|3|4|3.5|1|1|1|250|2|2|2|2|0|4|4|4|4|0|Red|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|52||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Black||40|28037|Bachelors Degree|Married|Medical: Doctor, Provider||2|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502590381|31|0|1|502625828|31|0|1|500544108|2||500004641||4|3|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|638794|291589|4|3|45
502605331|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-13|NaT|Followup|2014-08-13|2014-08-28|Complete|Done|1|1|1|1|1|3|1.33|3|4|4|1|3|3|3|-55.67|2|2|1|1|1|2|1.5|2|4|3|4|4|3|3.33|-54.95|3|3|3|3|4|4|4|4|-25|1|3|3|3|2.5|5|5|5|4|4.75|-47.37|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|3|4|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Red|Cabarrus County||55.1||1|1|1|1|M|Hispanic||13|No|Mother|28027|One Parent: Female|$25,000 to $29,999||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||33|28036|Bachelors Degree|Married|Business||2|5|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502605848|3|0|1|503090281|1|0|1|500627504|2||500016307||2|3|500016374|500016374|-2|500016374|-2|34|2|||7464|9|||1|639409|482204|4|3|45
502813454|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-13|NaT|Followup|2014-08-13|2014-08-13|Complete|Done|3|3|4|2|3|4|3.17|3|1|2|1|4|3|2.33|36.05|2|3|3|1|2|3|2.33|2|3|2|1|1|3|2|16.5|4|4|4|4|4|4|4|4|0|2|3|4|3|3|2|3|3|1|2.25|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|1|1|1|1|300|2|2|2|4|4|4|-50|2|2|1|1|100|4|4|4|4|0|Green|||55.1||1|2|1|2|F|White||14|No|Mother|28031|Two Parent|Unknown||Yes||School|General Community||Match Support|F|White||61|28031|Bachelors Degree|Divorced|Business: Mgt, Admin||5|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500020752|502814731|1|0|2|502855397|1|0|2|500627861|2||-2||2|1|||-2||-2|0|4|||129|1|||1|639430|390213|4|3|45
500771746|BBBS of Greater Charlotte|Main Office|C|Completed|2009-05-29|2016-06-15|Followup|2014-05-29|2014-05-29|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|3|1|2|3|2.33|||||||||4|4|4|4||||||1|2|1|1|1.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|4|3.33||||||1|3|2|||||2|2||||4|4||||Green|Project Big|Child: Graduated|84.6||3|4|1|2|F|Black||19||Mother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|F|White||37|28012|Some College|Married|Finance: Banking|28208|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500772014|31|0|2|500996153|1|0|2|500366437|2||500004641||4|1|500004640||-2||-2|0|4|||7464|9|||1|639717||4|3|45
502478700|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-09|2014-11-13|Followup|2014-08-09|2014-09-24|Declined|Late||||||||4|4|4|2|2|4|3.33|||||||||2|4|4|3|4|4|3.5||||||4|4|4|4|||||||5|4|5|5|4.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||2|2|2||||1|1||||4|4||Red|2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|39.2||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28027|Masters Degree|Single|Business: Engineer|28262|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|277|60|598|500000170|500013781|502881024|31|0|1|502578355|1|0|1|500544505|2||-2||4|3|500005291|500005291|-2|500015184|-1|0|5|||7462|13|||1|639978|315352|4|1|45
503355095|BBBS of Greater Charlotte|Main Office|C|Completed|2013-04-26|2016-05-02|Followup|2014-04-26|2014-06-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|36.2||1|1|1|1|F|Black||12|Yes|Mother|28212|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||36|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28202|5|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018851|503356940|31|0|2|503373533|31|0|2|500691042|2||-2||4|1||500000294|-2||-2|0|10|||7496|10|||1|639986||4|1|45
502619926|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-09|2015-05-05|Followup|2014-08-09|2014-10-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Project Big|Volunteer: Lost contact with child/agency|44.8||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||38|28205|Bachelors Degree|Single|Law: Lawyer|28202|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502620542|31|0|2|502642260|1|0|2|500548116|2||500004641||4|1|500004640||-2||-2|0|10|||7464|9|||1|640176||4|1|45
502637766|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-12|2017-01-24|Followup|2014-07-12|2014-07-23|Complete|Done|4|1|3|1|1|2|2|||||||||1|1|2|1|1|1|1.17|||||||||2|3|3|2.67||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|54.4||1|1|1|1|M|Black||13|No|Mother|28262|One Parent: Female|$50,000 to $59,999||Yes||School|General Community||Match Support|M|Black||34|28269|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500021785|502638462|31|0|1|503016558|31|0|1|500619500|2||-2||4|1|||-2||-2|0|4|||7462|13|||1|640352||4|3|45
502785308|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-16|NaT|Followup|2014-08-16|2014-08-22|Complete|Done|4|4|4|4|4|4|4|3|2|2|2|1|3|2.17|84.33|2|4|4|1|2|4|2.83|2|4|3|1|2|4|2.67|5.99|4|4|4|4|2|2|2|2|100|4|4|4|4|4|2|5|2|5|3.5|14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|Cabarrus County||55||1|2|1|2|F|American Indian or Alaska Native||16|No|Aunt|28027|One Parent: Male|Unknown||Yes||School|General Community|Cabarrus County|Match Support|F|White||49|28027|Bachelors Degree|Married|Business: Marketing|28025|14|0|ACN|Workplace Partner|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|504347632|6|0|2|502736971|1|0|2|500628695|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|4|||13581|3|||1|640423|359572|4|3|45
501195410|BBBS of Greater Charlotte|Main Office|C|Active|2008-08-15|NaT|Followup|2014-08-15|2014-08-29|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|5|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||103||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Asian||35|28210|Bachelors Degree|Married|Business: Sales|28217|5|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501195684|31|0|1|501277677|4|0|1|500278978|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|640578||4|3|45
503503500|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-26|2017-01-17|Baseline|2013-08-16|2013-08-26|Complete|Done|3|3|4|3|4|4|3.5|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|40.7||1|1|1|1|F|Black||15|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|White||37|28078|Bachelors Degree|Single|Medical|46285|6|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|503505371|31|0|2|503390470|1|0|2|500706999|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|640683|-1|4|3|44
502300563|BBBS of Greater Charlotte|Main Office|C|Active|2012-08-09|NaT|Followup|2014-08-09|2014-08-12|Complete|Done|1|4|4|4|3|3|3.17|3|3|4|1|3|4|3|5.67|3|4|3|3|3|4|3.33|4|4|3|4|3|4|3.67|-9.26|4|4|4|4|4|4|4|4|0|4|4|4|5|4.25|4|4|5|5|4.5|-5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|3|4|4|3.67|4|4|3|3.67|0|3|1|2|2|3|2.5|-20|2|2|1|1|100|4|4||||Green|||55.2||1|2|1|2|M|Black||15|No|Mother|28031|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Black||53|28078|PHD|Married|Medical|28078|2|0|AA Task Force|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020753|502300995|31|0|1|502101059|31|0|1|500626773|2||-2||2|1|||-2||-2|0|4|||11098|8|||1|641434|177594|4|3|45
503443162|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-20|2015-02-11|Followup|2014-08-20|2014-10-27|Declined|Late||||||||2|1|4|4|4|3|3|||||||||2|3|3|4|2|3|2.83||||||4|4|4|4|||||||3|4|3|2|3||||||||||4|4|4|3|4|3|2|3.43||||||4|3|4|3.67|||||1|1|1||||2|2||||4|4||Yellow||Child/Family: Lost contact with volunteer/agency|17.7||1|1|2|2|M|Black||17|No|Mother|28262|One Parent: Female|$25,000 to $29,999||Yes||Relative|General Community||Match Support|M|Black||34|28213|Bachelors Degree|Single|Finance: Banking|28202|0|2|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503445028|31|0|1|500234684|31|0|1|500705816|2||-2||4|2|||-2||-2|0|3|||7458|9|||1|641586|632640|4|1|45
502902247|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-11|NaT|Followup|2014-07-11|2014-08-29|Declined|Late||||||||2|4|4|2||2||||||||||3|4|3|3|3|3|3.17||||||4|4|4|4|||||||4|5|3|5|4.25||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||3|3|3||||1|1||||4|4||Green|||56.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||30|28203|Bachelors Degree|Single|Business: Marketing|28117|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502903657|31|0|2|502801082|1|0|2|500619356|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|641850|422744|4|1|45
503071350|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-22|2015-05-13|Followup|2014-08-22|2014-08-21|Complete|Done|4|2|4|2|4|4|3.33|||||||||2|3|3|4|2|4|3|||||||||4|4|4|4||||||4|5|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Time constraint|20.7||3|3|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||36|28210|Masters Degree|Divorced|Medical|28209|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|503073009|31|0|2|503421602|1|0|2|500705806|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|642060||4|3|45
503452963|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-22|2015-01-21|Followup|2014-08-22|2014-10-03|Declined|Done||||||||3|4|4|4|4|4|3.83|||||||||2|4|3|4|2|3|3||||||4|4|4|4|||||||5|4|4|4|4.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Red||Volunteer: Time constraint|17||1|1|1|1|M|Black||14|No|Mother|28211|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|M|Black||41|28216|Bachelors Degree|Single|Customer Service|28262|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500013781|503430105|31|0|1|503489818|31|0|1|500705904|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|642197|638157|4|1|45
502920377|BBBS of Greater Charlotte|Main Office|C|Completed|2012-06-29|2017-02-28|Followup|2014-06-29|2014-08-13|Declined|Done||||||||3|2|2|2|2|3|2.33|||||||||2|3|2|3|3|3|2.67||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||3||||||2|2||||4|4||Green||Volunteer: Lost contact with child/agency|56||1|1|1|1|F|Black||14|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||31|28211|Bachelors Degree|Single|Real Estate: Realtor|19137|2|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502921794|31|0|2|502942994|1|0|2|500620441|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|642612|439883|4|1|45
503014417|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-26|2016-08-17|Followup|2014-08-26|2014-08-26|Complete|Done|4|2|4|4|4|4|3.67|4|1|4|2|4|4|3.17|15.77|2|4|4|2|4|4|3.33|2|4|4|4|2|3|3.17|5.05|4|4|4|4|4|4|4|4|0|4|4|2|4|3.5|3|4|4|4|3.75|-6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|3|4|4|3.86|0|4|4|4|4|4|4|3|3.67|8.99|3|3|3|2|1|1.5|100|1|1|2|2|-50|4|4|4|4|0|Green||Child: Lost interest|35.7||1|1|1|1|F|Black||17|No|Mother|28203|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||29|28110|Masters Degree|Single|Education: Teacher||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|503015947|31|0|2|503518076|1|0|2|500706096|2||-2||4|1|||-2||-2|0|10|||46|2|||1|642883|638535|4|3|45
503484186|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-26|2016-03-08|Followup|2014-08-26|2014-08-26|Complete|Done|2|3|4|3|4|3|3.17|3|3|4|3|3|3|3.17|0|3|4|3|4|3|4|3.5|3|3|4|4|4|4|3.67|-4.63|4|4|4|4|4|4|4|4|0|5|5|4|5|4.75|5|5|5|4|4.75|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|4|4|-8.25|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Red||Child: Lost interest|30.4||1|1|1|1|M|White||16|No|Mother|28273|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|M|White||63|28226|Masters Degree|Widowed|Business: Marketing||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|503486052|1|0|1|503355490|1|0|1|500706097|2||-2||4|3|||-2||-2|0|10|||7671|13|1561|2|1|642966|627226|4|3|45
503503500|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-26|2017-01-17|Followup|2014-08-26|2014-09-05|Complete|Done|3|2|3|3|3|4|3|3|3|4|3|4|4|3.5|-14.29|3|4|3|3|3|4|3.33|3|3|4|4|4|4|3.67|-9.26|4|4|4|4|4|4|4|4|0|3|3|3|||5|4|5|5|4.75||4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|3|3.67|3|4|3|3.33|10.21|3|2|2.5|3|3|3|-16.67|||2|2||4|4|4|4|0|Green||Volunteer: Moved|40.7||1|1|1|1|F|Black||15|No|Mother|28216|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|White||37|28078|Bachelors Degree|Single|Medical|46285|6|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|503505371|31|0|2|503390470|1|0|2|500706999|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|642974|640683|4|3|45
501825910|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-24|2016-09-23|Followup|2014-08-24|2014-08-28|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|3|4|4|4|3.83|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Volunteer: Lost contact with child/agency|85||1|1|1|1|M|Black||16|Yes|Mother|28213|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|M|White||51|28214|Masters Degree|Married|Business: Sales|94108|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500188141|31|0|1|501196986|1|0|1|500380446|2||500003586||4|2|500000294|500000294|-2|500000294|-2|0|10|||7496|10|||1|643233||4|3|45
502601023|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-31|2016-08-11|Followup|2014-08-31|2014-08-21|Complete|Done|3|2|3|2|3|3|2.67|3|2|3|1|3|4|2.67|0|2|4|3|2|2|4|2.83|3|3|4|2|2|3|2.83|0|4|4|4|4|4|4|4|4|0|3|3|4|4|3.5|3|3|4|5|3.75|-6.67|4|4|4|4|4|4|3|3.86|4|2|4|4|3|4|3|3.43|12.54|3|4|3|3.33|3|4|2|3|11|2|3|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child: Graduated|59.4||1|1|1|1|F|Black||19||Mother|28216|Two Parent|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||51|28277|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502601540|31|0|2|502546883|1|0|2|500550809|2||-2||4|1|500005291|500005291|-2||-2|6854|8|||7464|9|||1|643347|331012|4|3|45
502591898|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-18|NaT|Followup|2014-07-18|2014-09-04|Declined|Late||||||||3|3|4|2|3|4|3.17|||||||||4|3|4|2|4|4|3.5||||||4|4|4|4|||||||5|5|4|5|4.75||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Green|||55.9||2|2|1|1|F|Black||16|No|Mother|28214|Two Parent|$40,000 to $44,999|Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28210|Masters Degree|Single|Medical: Healthcare Worker||1|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|502592415|31|0|2|503002003|31|0|2|500620503|2||-2||2|1||500004640, 500005291|-2||-2|0|4|||7496|10|||1|643866|294647|4|1|45
502255223|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-11|NaT|Followup|2014-08-11|2014-09-25|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||79.1||1|1|1|1|F|Hispanic||14|No|Mother|28212|One Parent: Female|Unknown|Y|No|Spanish Radio|Media|General Community||Match Support|F|White||33|28209||Single|Education: Teacher||0|0||High School Partner|Big|General Community||Match Support|277|60|598|500000170|500020753|502255655|3|0|2|501823103|1|0|2|500463922|2||-2||2|1|||-2||-2|7068|1|||0|4|||1|643903||4|1|45
503512877|BBBS of Greater Charlotte|Main Office|C|Completed|2014-07-11|2016-11-10|Baseline|2013-08-29|2014-07-11|Complete|Done|3|2|4|1|4|4|3|||||||||1|4|4|1|1|4|2.5|||||||||4|3|3|3.33||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|28||1|1|1|1|M|Black||12|No|Mother|28211|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|M|White||27|28226|Bachelors Degree|Single|Tech: Research/Design|28269|0|8|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500021785|503514748|31|0|1|503893014|1|0|1|500766726|2||-2||4|1|||-2||-2|0|10|||17101|1|||1|644026|-1|4|3|44
501994951|BBBS of Greater Charlotte|Main Office|C|Completed|2010-06-15|2014-09-18|Followup|2014-06-15|2014-07-29|Complete|Done|4|4|4|3|4|4|3.83|3|3|3|1|4|4|3|27.67|3|4|4|3|1|4|3.17|4|4|3|4|4|4|3.83|-17.23|4|3|3|3.33|4|4|4|4|-16.75|3|4|4|3|3.5|4|5|5|4|4.5|-22.22|4|4|4|4|4|3|3|3.71|4|4|4|3|3|3|3|3.43|8.16|3|4|3|3.33|3|3|3|3|11|2|2|2|3|1|2|0|2|2|1|1|100|4|4||||Yellow||Volunteer: Lost contact with child/agency|51.1||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|Unknown||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||36|28078||Single|Customer Service||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|501843047|31|0|2|502048623|31|0|2|500455478|2||-2||4|2|||-2||-2|7294|13|||7464|9|||1|644347|139614|4|3|45
502990571|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-30|2016-08-11|Followup|2014-08-30|2014-08-28|Complete|Done|2|1|2|2|2|2|1.83|3|3|2|1|2|1|2|-8.5|2|1|2|3|2|2|2|3|3|4|3|4|4|3.5|-42.86|4|4|4|4|4|4|4|4|0|1|4|3|4|3|5|4|4|5|4.5|-33.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|2|2|3|2.33|4|4|4|4|-41.75|3|3|3|3|2|2.5|20|2|2|1|1|100|4|4|4|4|0|Red||Child/Family: Moved|35.4||2|2|1|1|F|Multi-race (Black & Hispanic)||15|Yes|Mother|28217|Two Parent|$35,000 to $39,999||Yes||Self|General Community||Match Support|F|Black||28|28269|Bachelors Degree|Single|Business||0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502992028|38|0|2|503400909|31|0|2|500707095|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|644408|460382|4|3|45
501288021|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-27|2016-02-01|Followup|2014-08-27|2014-08-25|Complete|Done|4|4|4|4|3|4|3.83|||||||||2|3|3|3|2|4|2.83|||||||||4|4|4|4||||||4|5|2|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Moved|89.2||1|1|1|1|F|Black||16|No|Mother|28211|Two Parent|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28027|PHD|Single|Education: College Professor|27411|1|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|501288299|31|0|2|501249338|31|0|2|500281778|2||-2||4|1|||-2||-2|0|10|||46|2|||1|644472||4|3|45
502245343|BBBS of Greater Charlotte|Main Office|C|Active|2011-05-05|NaT|Followup|2014-05-05|2014-06-19|Complete|Done|3|3|3|2|3|3|2.83|||||||||2|3|3|2|3|3|2.67|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|Amachi||70.4||1|1|1|1|M|Black||12|Yes|Mother|28216|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|M|White||32|28104|Bachelors Degree|Single|Business|28216|5|3|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502245774|31|0|1|502526001|1|0|1|500532810|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||17161|11|||1|644826||4|3|45
503044619|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-03|2016-09-15|Followup|2014-08-03|2014-09-18|Declined|Late||||||||3|1|4|1|2|2|2.17|||||||||4|4|4|4|4|4|4||||||3|2|4|3|||||||4|5|3|5|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||1|4|2.5||||2|2||||4|4||Green||Child/Family: Moved|49.4||1|1|1|1|M|Black||15|No|Mother|28205|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance: Banking|28202|0|7|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020910|503046265|31|0|1|503021454|1|0|1|500624634|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|644969|474027|4|1|45
502252828|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-03|2015-10-13|Followup|2014-08-03|2014-09-17|Complete|Done|3|2|4|2|4|4|3.17|4|1|4|4|1|2|2.67|18.73|3|4|4|2|2|4|3.17|1|2|1|2|2|2|1.67|89.82|4|4|4|4|1|1|1|1|300|4|4|3|4|3.75|4|3|2|1|2.5|50|4|4|4|4|3|4|4|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|2|2|3|2.33|71.67|3|3|3|4|3|3.5|-14.29|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Volunteer: Time constraint|50.3||1|1|1|1|M|Black||15||GrandMother|28227|Grandparents|Unknown||No||Self|General Community|PERL 2014-2016|RTBM|M|White||27|28205|Associate Degree|Single|Law: Police Officer||0|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|277|60|598|500000170|500017777|502253254|31|0|1|502602451|1|0|1|500547383|2||-2||4|1|500005291|500014681|-2|500005291|-2|0|10|||7496|10|||1|644970|320066|4|3|45
502431187|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-17|2016-01-07|Followup|2014-08-17|2014-09-30|Complete|Done|3|1|3|2|3|2|2.33|3|2|4|1|3|4|2.83|-17.67|2|3|3|3|3|3|2.83|2|3|3|2|3|3|2.67|5.99|4|4|4|4|2|4|4|3.33|20.12|3|2|3|3|2.75|4|3|5|3|3.75|-26.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|3|3.33|3|2|3|2.67|24.72|3|2|2.5|2|3|2.5|0|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Time constraint|40.7||2|2|1|1|F|Black||17|No|GrandMother|28208|One Parent: Female|Unknown||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|RTBM|F|White||41|28105|Bachelors Degree|Divorced|Business|28112|1|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|502431630|31|0|2|503015009|1|0|2|500627361|2||-2||4|2||500005291|-2||-2|0|5|||46|2|||1|644973|272216|4|3|45
502000252|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-22|NaT|Followup|2014-08-22|2014-08-22|Complete|Done|3|3|4|2|4|4|3.33|||||||||2|3|3|2|3|3|2.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||3|4|4|3.67||||||3|1|2|||||2|2||||4|4||||Green|||78.8||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500020910|502000651|31|0|1|502127058|1|0|1|500465318|2||-2||2|1|||-2||-2|0|10|||130|1|||1|644976||4|3|45
503496889|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-25|2015-05-29|Baseline|2013-09-03|2013-09-25|Complete|Done|3|4|4|4|3|4|3.67|||||||||2|4|2|2|2|4|2.67|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Moved|20.1||1|1|1|1|M|Black||16|No|Mother|28273|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|White||28|28207|Bachelors Degree|Single|Education: Teacher||1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503498757|31|0|1|503490051|1|0|1|500708903|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|645105|-1|4|3|44
501809541|BBBS of Greater Charlotte|Main Office|C|Active|2009-08-07|NaT|Followup|2014-08-07|2014-10-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||91.3||1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|M|White||49|28031|Bachelors Degree|Married|Transport: Pilot|40223|9|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501809896|36|0|1|501620528|1|0|1|500375025|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|645151||4|1|45
502593613|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-19|2017-02-28|Followup|2014-08-19|2014-11-03|Expired|Late||||||||3|2||1|2|2||||||||||3|3|3|3|3|3|3||||||4|4|4|4|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|4|4||||||4|3|3|3.33|||||3|3|3||||2|2||||4|4||Yellow||Volunteer: Lost contact with child/agency|66.4||1|1|1|1|F|Black||16|No|Mother|28208|Two Parent|$35,000 to $39,999|Y|Yes||Relative|General Community||Match Support|F|Hispanic||26|28217|Bachelors Degree|Single|Service: Restaurant||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502594130|31|0|2|502601730|3|0|2|500547881|2||-2||4|2|||-2||-2|0|3|||7464|9|||1|645153|322561|4|0|45
500881634|BBBS of Greater Charlotte|Main Office|C|Active|2008-07-14|NaT|Followup|2014-07-14|2014-07-25|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|2|4|4|3.67|||||||||4|3|3|3.33||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|||104||1|2|1|2|M|Black||18||Mother|28213|Other/Unknown|Unknown||No||School|General Community||Match Support|F|Black||38|28213||Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|500881903|31|0|1|500816190|31|0|2|500277615|2||-2||2|1|||-2||-2|0|4|||46|2|||1|645154||4|3|45
500186435|BBBS of Greater Charlotte|Main Office|C|Completed|2003-07-23|2015-08-20|Followup|2014-07-23|2014-07-24|Complete|Done|3|4|4|4|3|1|3.17|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|144.9||1|1|1|1|M|Black||20||Mother|28216|One Parent: Female|Unknown||No|Brochure|Media|General Community||Match Support|M|White||45|28226|Bachelors Degree|Married|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187988|31|0|1|500189358|1|0|1|500037395|2||-2||4|1|||-2||-2|51|1|||7496|10|||1|645157||4|3|45
500395038|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-01|2015-02-20|Followup|2014-08-01|2014-10-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|102.7||1|1|1|1|M|White||20||Mother|28226|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|M|White||39|28211|Masters Degree|Married|Law: Lawyer|28204|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500395288|1|0|1|500392006|1|0|1|500104016|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|645158||4|1|45
500835156|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-10|2016-11-10|Followup|2014-07-10|2014-07-17|Complete|Done|2|4|4|4|4|4|3.67|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|100||1|2|1|2|M|Black||17||Mother|28217|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Multi-Race (None of the above)||38|29710|Bachelors Degree|Single|Architect||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500835425|31|0|1|500466903|7|0|1|500277232|2||-2||4|1|||-2||-2|0|4|||46|2|||1|645190||4|3|45
500915359|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-10|2014-12-18|Followup|2014-08-10|2014-10-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|28.3||3|3|1|1|F|Black||19|No|Mother|28227|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28204|Bachelors Degree|Single|Medical: Nurse||0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500915629|31|0|2|503044413|1|0|2|500622861|2||-2||4|2|||-2||-2|34|2|||7496|10|||1|645191||4|1|45
502215233|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-16|2014-12-17|Baseline|2013-09-04|2013-09-16|Complete|Done|3|3|2|2|4|3|2.83|||||||||2|3|3|3|4|3|3|||||||||4|4|4|4||||||3|4|3|2|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|15||2|2|1|1|F|Hispanic|Other South American|14|No|Mother|28212|Two Parent|Unknown||Yes|Big|Neighbor/Friend|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|White||34|28270||Married|Unknown|28236|1|0|Big For A Day|Special Event|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500017777|502215660|3|15|2|503558339|1|0|2|500709090|2||-2||4|3||500011312, 500014681|-2|500000294|-2|6854|8|||16422|8|||1|645412|-1|4|3|44
501721760|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-22|2016-11-01|Followup|2014-06-22|2014-06-26|Complete|Done|4|2|4|2|4|4|3.33|||||||||2|4|3|1|1|3|2.33|||||||||4|4|3|3.67||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Infraction of match rules/agency policies|88.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||59|28269|Masters Degree|Married|Clergy||0|0|Coca Cola|Workplace Partner|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|501722098|31|0|1|501755476|1|0|1|500368545|2||-2||4|1|||-2|500000294|-2|0|10|||9610|3|||1|645940||4|3|45
500910037|BBBS of Greater Charlotte|Main Office|C|Active|2009-06-22|NaT|Followup|2014-06-22|2014-07-07|Complete|Done|2|3|4|4|2|3|3|||||||||2|4|3|2|2|3|2.67|||||||||4|4|4|4||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|2|3||||||4|4|4|||||2|2||||4|4||||Green|||92.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|M|White||46|28277||Married|Business: Mgt, Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|500910307|31|0|1|500856100|1|0|1|500368834|2||-2||2|1|||-2||-2|0|10|||46|2|||1|645941||4|3|45
501160242|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-09|2016-11-07|Followup|2014-08-09|2014-09-03|Complete|Done|3|2|1|2|1|2|1.83|||||||||2|3|3|3|2|3|2.67|||||||||3|3|3|3||||||2|3|3|5|3.25|||||||4|4|4|4|4|4|4|4||||||||||2|3|2|2.33||||||2|4|3|||||2|2||||4|4||||Red|Cabarrus County|Volunteer: Lost contact with child/agency|51||3|4|1|2|F|White||17|No|GrandFather|28147|Grandparents|Unknown||No||School|General Community|Cabarrus County|Match Support|F|White||29|28078||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501160516|1|0|2|502325100|1|0|2|500626774|2||500016307||4|3|500016374|500016374|-2|500016374|-2|0|4|||7496|10|||1|646163||4|3|45
501641325|BBBS of Greater Charlotte|Main Office|C|Completed|2009-06-24|2015-08-03|Followup|2014-06-24|2014-09-08|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|73.3||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Multi-race (Asian & White)||34|28205|Bachelors Degree|Single|Tech: Research/Design|28255|3|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|1|501715652|37|0|1|500366872|2||-2||4|1||500000294|-2|500000294|-2|6854|8|||7464|9|||1|646315||4|0|45
501721579|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-24|2016-06-17|Followup|2014-07-24|2014-09-08|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Volunteer: Moved|82.8||2|2|1|1|F|Multi-Race (None of the above)||14|No|Mother|28211|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||50|28227|Some College|Single|Human Services: Social Worker||2|5|St. Paul Baptist|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501721919|7|0|2|501687513|31|0|2|500375006|2||500003586||4|3|500000294|500000294|-2|500000294|-2|5635|9|||9609|7|||1|646361||4|1|45
503421607|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-26|2017-02-28|Baseline|2013-09-09|2013-09-25|Complete|Done|2|2|1|1|2|4|2|||||||||3|3|3|2|1|4|2.67|||||||||4|3|3|3.33||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||2|2||||4|4||||Green||Child: Family structure changed|41.1||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28214|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|F|Black||49|28273|Associate Degree|Single|Finance: Accountant|28273|7|0|Agency Sponsored|Special Event|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503423471|36|0|2|503520561|31|0|2|500711787|2||-2||4|1|||-2|500000294|-2|0|10|||16426|8|||1|646424|-1|4|3|44
500465506|BBBS of Greater Charlotte|Main Office|C|Active|2006-08-21|NaT|Followup|2014-08-21|2014-08-20|Complete|Done|3|4|4|4|3|4|3.67|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|5|3|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Yellow|Amachi||126.8||1|1|1|1|M|Black||16|Yes|Mother|28262|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||54|28226|Bachelors Degree|Married|Arts, Entertainment, Sports||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500465757|31|0|1|500496966|1|0|1|500118121|2||500003586||2|2|500000294|500000294|-2|500000294|-2|0|4|||2238|7|||1|646483||4|3|45
502907527|BBBS of Greater Charlotte|Main Office|C|Completed|2012-08-23|2014-11-21|Followup|2014-08-23|2014-09-02|Complete|Done|4|2|4|2|4|4|3.33|4|1|4|1|4|4|3|11|2|4|3|4|2|3|3|4|4|4|4|1|4|3.5|-14.29|4|4|4|4|4|4|4|4|0|3|5|4|4|4|3|5|3|3|3.5|14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|3|3.5|4|4|4|-12.5|2|2|2|2|0|4|4|4|4|0|Yellow||Volunteer: Moved|26.9||1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community|Amachi|Match Support|M|White||55|28202|Associate Degree|Married|Business||30|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502908938|31|0|1|502996593|1|0|1|500624606|2||-2||4|2||500000294|-2||-2|0|10|||7464|9|||1|646538|473967|4|3|45
503476243|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-20|2015-04-23|Baseline|2013-09-10|2013-09-20|Complete|Done|3|3|2|4|3|3|3|||||||||3|3|4|3|4|4|3.5|||||||||4|4|4|4||||||3|5|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|3|3|3.33||||||1|3|2|||||1|1||||4|4||||Red||Child: Lost interest|19.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|White||63|28210|Bachelors Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|503478109|31|0|1|503334174|1|0|1|500710120|2||-2||4|3|||-2||-2|0|10|||7671|13|1561|2|1|646966|-1|4|3|44
503472232|BBBS of Greater Charlotte|Main Office|C|Completed|2013-06-17|2016-08-08|Followup|2014-06-17|2014-07-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|37.7||1|1|1|1|M|Black||12||Mother|28217|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||48|28273|Some College|Divorced|Transport: Driver|29730|3|0|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|503474098|31|0|1|503444888|31|0|1|500700046|2||-2||4|3|||-2||-2|34|2|||130|1|||1|647079||4|1|45
501842678|BBBS of Greater Charlotte|Main Office|C|Completed|2011-06-27|2015-06-19|Followup|2014-06-27|2014-07-29|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|3|3.67||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|3|3|||||2|2|||||||||Yellow||Volunteer: Feels incompatible with child/family|47.7||2|2|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown|Y|No||Self|General Community||Match Support|M|White||53|28117|Bachelors Degree|Married|Real Estate: Realtor|28031|0|0|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|277|60|598|500000170|500015820|501843047|31|0|1|502335257|1|0|1|500542227|2||-2||4|2|||-2|500000294, 500004901|-2|0|10|||7464|9|||1|647117||4|3|45
503361148|BBBS of Greater Charlotte|Main Office|C|Active|2013-09-24|NaT|Baseline|2013-09-11|2013-09-24|Complete|Done|3|2|4|2|3|4|3|||||||||2|3|3|2|3|2|2.5|||||||||2|2|2|2||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|2|3|||||2|2||||4|4||||Green|||41.7||1|1|2|2|M|Multi-race (Black & Hispanic)||14|No|Mother|28273|One Parent: Female|$50,000 to $59,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|503362993|38|0|1|502459922|1|0|1|500710308|2||-2||2|1|||-2|500004640|-2|34|2|||7464|9|||1|647241|-1|4|3|44
503497835|BBBS of Greater Charlotte|Main Office|C|Active|2013-09-19|NaT|Baseline|2013-09-11|2013-09-19|Complete|Done|3|1|2|1|3|2|2|||||||||1|2|2|2|1|2|1.67|||||||||4|3|2|3||||||2|4|4|5|3.75|||||||4|4|4|4|4|3|2|3.57||||||||||3|3|4|3.33||||||3|2|2.5|||||1|1||||4|4||||Green|||41.9||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|F|Black||26|28209|Bachelors Degree|Single|Retail: Sales|28210|0|10|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|503499703|31|0|2|503507978|31|0|2|500710423|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|647341|-1|4|3|44
502179379|BBBS of Greater Charlotte|Main Office|C|Completed|2010-07-25|2015-07-31|Followup|2014-07-25|2014-09-09|Declined|Late||||||||4|4|4|4|2|4|3.67|||||||||1|4|4|1|2|4|2.67||||||4|4|4|4|||||||3|3|5|5|4||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||1|2|1.5||||2|2|||||||Red|Project Big|Volunteer: Lost contact with child/agency|60.2||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|Black||34|28269||Single|Student: College||0|0|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|502179808|31|0|2|502161458|31|0|2|500461681|2||-2||4|3|500004640|500004640|-2||-2|0|10|||9221|5|||1|648207|158340|4|1|45
502234504|BBBS of Greater Charlotte|Main Office|C|Active|2010-07-28|NaT|Followup|2014-07-28|2014-09-12|Complete|Late|4|2|2|2|3|4|2.83|4|4|4|4|2|4|3.67|-22.89|2|4|4|2|3|3|3|1|4|4|1|2|4|2.67|12.36|4|4|4|4|4|4|4|4|0|3|3|3|3|3|3|3|5|5|4|-25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|4|3.67|8.99|3|3|3|1|3|2|50|2|2|2|2|0|4|4||||Yellow|Project Big||79.6||1|1|2|2|F|Black||16|No|GrandMother|28208|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|Project Big|Match Support|F|Black||37|28216|Bachelors Degree|Single|Customer Service||8|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|277|60|598|500000170|500008321|502234935|31|0|2|502129464|31|0|2|500463451|2||500004641||2|2|500004640|500004640|-2||-1|0|4|||11247|3|1204|3|1|648209|155881|4|3|45
502863781|BBBS of Greater Charlotte|Main Office|C|Completed|2012-07-31|2015-01-30|Followup|2014-07-31|2014-09-14|Complete|Done|3|4|4|3|4|4|3.67|3|4|3|2|3|4|3.17|15.77|2|3|3|3|3|3|2.83|2|4|3|2|1|2|2.33|21.46|4|4|4|4|4|4|4|4|0|2|3|3|2|2.5|2|3|3|2|2.5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|4|3|3.33|0|2|3|2.5|4|4|4|-37.5|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Time constraint|30||1|1|1|1|M|Black||18|No|Mother|28031|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|M|White||26|28031|High School Graduate|Single|Personal Trainer/Coach|28117|0|4|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500008321|502865175|31|0|1|503002010|1|0|1|500621061|2||-2||4|3|||-2||-2|0|10|||17161|11|||1|648210|465050|4|3|45
502863776|BBBS of Greater Charlotte|Main Office|C|Active|2012-07-31|NaT|Followup|2014-07-31|2014-09-14|Complete|Done|3|2|3|2|4|4|3|2|2|3|4|3|4|3|0|2|3|3|4|4|3|3.17|2|3|3|3|3|3|2.83|12.01|4|4|4|4|4|4|4|4|0|3|5|4|4|4|3|5|3|4|3.75|6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|3|4|3|3.33|0|2|2|2|1|1|1|100|2|2|1|1|100|4|4|4|4|0|Green|||55.5||1|1|1|1|F|Black||14|No|Mother|28031|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Mgt, Admin|28078|1|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502865175|31|0|2|503029273|1|0|2|500622877|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|648211|434619|4|3|45
500958307|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-19|NaT|Followup|2014-09-19|2014-09-19|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|1|4|3|2.83|||||||||4|4|4|4||||||3|3|2|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi, Cabarrus County||113.9|Y|1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$40,000 to $44,999|Y|No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|Black||62|28213||Married|Finance: Economist||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|277|60|598|500000170|500022817|500958577|31|0|1|500876132|31|0|1|500193868|2||500003586||2|1|500000294, 500016374|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|648556||4|3|45
502215233|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-16|2014-12-17|Followup|2014-09-16|2014-12-01|Expired|Late||||||||3|3|2|2|4|3|2.83|||||||||2|3|3|3|4|3|3||||||4|4|4|4|||||||3|4|3|2|3||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Red||Volunteer: Feels incompatible with child/family|15||2|2|1|1|F|Hispanic|Other South American|14|No|Mother|28212|Two Parent|Unknown||Yes|Big|Neighbor/Friend|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|White||34|28270||Married|Unknown|28236|1|0|Big For A Day|Special Event|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500017777|502215660|3|15|2|503558339|1|0|2|500709090|2||-2||4|3||500011312, 500014681|-2|500000294|-2|6854|8|||16422|8|||1|648766|645412|4|0|45
503425736|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-16|2016-06-15|Baseline|2013-09-17|2013-09-28|Complete|Done|3|3|4|2|4|4|3.33|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4|3|2|3|3|||||||2|2|2|2|2|2|2|2||||||||||1|2|2|1.67||||||4|2|3|||||1|1||||4|4||||Green||Child: Graduated|32||1|1|1|1|F|Black||18|No|GrandMother|28213|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|White||29|28211|Juris Doctorate (JD)|Married|Law|28202|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|503427601|31|0|2|503519747|1|0|2|500711543|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|649102|-1|4|3|44
502529397|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-11|NaT|Followup|2014-08-11|2014-08-12|Complete|Done|3|4|4|3|1|3|3|||||||||2|4|3|4|3|3|3.17|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|Project Big||67.2||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||48|28216|Bachelors Degree|Married|Finance: Banking|28255|8|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502529850|31|0|1|500188946|31|0|1|500548763|2||500004641||2|1|500004640||-2||-2|6854|8|||7464|9|||1|649406||4|3|45
502455004|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-20|NaT|Followup|2014-09-20|2014-10-19|Complete|Done|4|4|4|2|4|4|3.67|4|2|4|1|1|4|2.67|37.45|2|4|4|2|2|1|2.5|4|4|4|2|4|4|3.67|-31.88|4|4|4|4|4|4|4|4|0|5|4|3|4|4|5|5|4|5|4.75|-15.79|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||65.8||1|1|1|1|M|Black|Other African|15|No|Mother|29732|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|29720|Bachelors Degree|Married|Business: Sales|28134|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502074089|31|31|1|502680045|1|0|1|500553363|2||-2||2|1|500005291|500005291|-2||-2|0|4|||7464|9|||1|649638|336027|4|3|45
503497835|BBBS of Greater Charlotte|Main Office|C|Active|2013-09-19|NaT|Followup|2014-09-19|2014-09-16|Complete|Done|4|4|4|4|4|3|3.83|3|1|2|1|3|2|2|91.5|3|4|4|3|3|4|3.5|1|2|2|2|1|2|1.67|109.58|4|4|4|4|4|3|2|3|33.33|4|4|4|5|4.25|2|4|4|5|3.75|13.33|3|4|4|4|4|4|3|3.71|4|4|4|4|4|3|2|3.57|3.92|4|4|4|4|3|3|4|3.33|20.12|3|3|3|3|2|2.5|20|2|2|1|1|100|4|4|4|4|0|Green|||41.9||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|F|Black||26|28209|Bachelors Degree|Single|Retail: Sales|28210|0|10|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|503499703|31|0|2|503507978|31|0|2|500710423|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|649845|647341|4|3|45
503476243|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-20|2015-04-23|Followup|2014-09-20|2014-10-02|Complete|Done|3|4|4|2|4|3|3.33|3|3|2|4|3|3|3|11|4|4|3|4|2|4|3.5|3|3|4|3|4|4|3.5|0|4|4|4|4|4|4|4|4|0|2|5|4|5|4|3|5|4|3|3.75|6.67|4|4|4|4|3|4|4|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|3|3|3.33|20.12|3|2|2.5|1|3|2|25|2|2|1|1|100|4|4|4|4|0|Red||Child: Lost interest|19.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|White||63|28210|Bachelors Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|503478109|31|0|1|503334174|1|0|1|500710120|2||-2||4|3|||-2||-2|0|10|||7671|13|1561|2|1|650217|646966|4|3|45
502347820|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-20|2016-02-08|Followup|2013-12-20|2014-03-06|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Moved|49.6||3|3|2|2|F|Black||12|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Some Other Race||75|28213|Some College|Widowed|Human Services||20|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020990|502348258|31|0|2|502419409|41|0|2|500588112|2||500003586||4|2|500000294|500000294|-2||-2|0|10|||7464|9|||1|650496||4|0|45
502789637|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-23|2015-08-25|Followup|2014-09-23|2014-09-23|Complete|Done|4|4|4|4|1|4|3.5|||||||||1|1|2|4|4|4|2.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|23||4|4|2|2|F|Black||12|No|Mother|28081|One Parent: Female|Less than $10,000||Yes||School|General Community|Cabarrus County|Match Support|F|Black||30|28027|Masters Degree|Married|Unemployed|28027|2|5|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500012459|502790820|31|0|2|503542037|31|0|2|500708902|2||-2||4|2||500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||7464|9|||1|650729||4|3|45
501604443|BBBS of Greater Charlotte|Main Office|C|Active|2009-07-10|NaT|Followup|2014-07-10|2014-08-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||92.2||1|1|1|1|M|Black||18|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||35|28209|Bachelors Degree|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501729878|1|0|1|500371104|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|651073||4|1|45
503361148|BBBS of Greater Charlotte|Main Office|C|Active|2013-09-24|NaT|Followup|2014-09-24|2014-11-07|Complete|Done|3|2|4|2|3|4|3|3|2|4|2|3|4|3|0|2|4|3|3|4|4|3.33|2|3|3|2|3|2|2.5|33.2|4|4|||2|2|2|2||3|3|3|4|3.25|3|2|4|4|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|3|3|3|11|3|3|3|4|2|3|0|2|2|2|2|0|4|4|4|4|0|Green|||41.7||1|1|2|2|M|Multi-race (Black & Hispanic)||14|No|Mother|28273|One Parent: Female|$50,000 to $59,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|503362993|38|0|1|502459922|1|0|1|500710308|2||-2||2|1|||-2|500004640|-2|34|2|||7464|9|||1|651217|647241|4|3|45
501261979|BBBS of Greater Charlotte|Main Office|C|Completed|2008-07-22|2014-10-13|Followup|2014-07-22|2014-07-22|Complete|Done|1|4|4|2|3|4|3|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Moved|74.7||1|1|3|3|F|Black||15|No|Mother|28134|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|Black||55|28173||Married|Human Services: Non-Profit|28205|0|0|Coworker|Workplace Partner|Big|General Community|VOL - Maximizing Match Impact|Match Support|277|60|598|500000170|500011349|501262256|31|0|2|500418936|31|0|2|500278634|2||-2||4|1|||-2|500011314|-2|0|10|||7447|3|||1|651299||4|3|45
500961274|BBBS of Greater Charlotte|Main Office|C|Active|2007-08-27|NaT|Followup|2014-08-27|2014-08-26|Complete|Done|4|3|4|2|4|4|3.5|||||||||3|4|4|4|2|4|3.5|||||||||4|4|4|4||||||3|4|4|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi||114.6||1|1|2|2|F|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||51|28216|Bachelors Degree|Divorced|Business: Clerical|28204|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500934638|31|0|2|500403000|31|0|2|500186952|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|651361||4|3|45
503496889|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-25|2015-05-29|Followup|2014-09-25|2014-11-07|Complete|Done|4|3|3|2|4|4|3.33|3|4|4|4|3|4|3.67|-9.26|3|4|4|4|3|4|3.67|2|4|2|2|2|4|2.67|37.45|4|3|3|3.33|4|4|4|4|-16.75|4|4|5|5|4.5|4|4|5|5|4.5|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|4|4|4|2|2|2|100|2|2|2|2|0|||4|4||Green||Volunteer: Moved|20.1||1|1|1|1|M|Black||16|No|Mother|28273|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|White||28|28207|Bachelors Degree|Single|Education: Teacher||1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503498757|31|0|1|503490051|1|0|1|500708903|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|651486|645105|4|3|45
503524258|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-30|2016-01-26|Baseline|2013-09-25|2013-09-28|Complete|Done|3|4|4|1|1|3|2.67|||||||||1|1|4|1|1|4|2|||||||||3|4|4|3.67||||||5|3|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||2|4|1|2.33||||||4|4|4|||||1|1||||4|4||||Green||Volunteer: Moved|27.9||1|1|3|3|F|Black||14|No|Mother|28217|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Black||34|28273|Bachelors Degree|Single|Retail: Mgt|28217|5|6|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|503526133|31|0|2|500497043|31|0|2|500713184|2||-2||4|1||500000294|-2||-2|34|2|||6247|12|||1|651722|-1|4|3|44
503575828|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-28|2014-12-17|Baseline|2013-09-25|2013-09-28|Complete|Done|3|3|4|4|3|4|3.5|||||||||4|4|4|3|2|4|3.5|||||||||4|3|3|3.33||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Green||Volunteer: Moved|14.6||3|3|1|1|M|Hispanic||13|No|Mother|28206|One Parent: Female|Unknown||Yes|Spanish Radio|Media|General Community|PERL 2014-2016|Match Support|M|White||26|28203|Bachelors Degree|Single|Finance: Banking|28202|0|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|503577713|3|0|1|503576000|1|0|1|500713280|2||-2||4|1||500014681|-2|500000294|-2|7068|1|||7464|9|||1|651809|-1|4|3|44
503207102|BBBS of Greater Charlotte|Main Office|C|Inactive|2014-04-11|NaT|Baseline|2013-09-25|2014-04-11|Complete|Done|2|1|1|1|1|1|1.17|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||3|5|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|||35.2||1|1|1|1|M|Multi-race (Black & Hispanic)||12|No|Mother|28270|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|White||54|28110|Some College|Married|Self-Employed, Entrepreneur|28110|11|6|Relative|Relative|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|277|60|598|500000170|500017777|503208876|38|0|1|503688236|1|0|1|500757797|2||-2||3|1|||-2|500011312|-2|0|10|||17161|11|||1|651875|-1|4|3|44
502245129|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-22|NaT|Followup|2014-08-22|2014-08-21|Complete|Done|4|4|4|4|3|3|3.67|4|3|4|2|3|3|3.17|15.77|2|4|3|3|3|4|3.17|1|4|3|2|4|3|2.83|12.01|4|4|3|3.67|4|3|2|3|22.33|4|5|3|5|4.25|5|4|3|2|3.5|21.43|4|4|4|4|4|4|2|3.71|4|3|4|3|2|4|3|3.29|12.77|4|4|4|4|4|4|3|3.67|8.99|3|2|2.5|4|3|3.5|-28.57|2|2|1|1|100|4|4|4|4|0|Green|Amachi||66.8||1|1|1|1|M|Multi-race (Black & Hispanic)||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||28|28262|High School Graduate|Single|Laborer||0|8|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020752|502245570|38|0|1|502670839|31|0|1|500551050|2||-2||2|1|500000294||-2||-2|0|10|||7671|13|||1|651947|331272|4|3|45
502221847|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-27|NaT|Followup|2014-09-27|2014-09-29|Complete|Done|4|2|4|1|4|4|3.17|3|1|2|1|4|2|2.17|46.08|4|3|4|4|3|4|3.67|4|4|4|2|4|4|3.67|0|4|1|1|2|4|4|4|4|-50|4|3|2|3|3|5|4|5|5|4.75|-36.84|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|2|3|1|2|3|4|4|3.67|-45.5|3|3|3|2|4|3|0|2|2|2|2|0|4|4||||Green|Amachi||65.6||2|2|1|1|F|Black||16|Yes|GrandMother|28213|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||24|28027|Some College|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502222278|31|0|2|502654877|31|0|2|500556560|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|652149|154081|4|3|45
501831581|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-29|NaT|Followup|2014-09-29|2014-10-02|Complete|Done|4|4|4|4|2|3|3.5|||||||||3|3|3|3|4|3|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi||89.5||1|1|2|3|F|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||38|28273||Single|Tech: Engineer||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|501831944|31|0|2|500715453|31|0|2|500387624|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||46|2|||1|652153||4|3|45
501604440|BBBS of Greater Charlotte|Main Office|C|Completed|2009-07-23|2014-11-19|Followup|2014-07-23|2014-10-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|63.9||1|1|1|1|M|Black||20|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||38|28269||Married|Govt||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|501604760|31|0|1|501758365|3|0|1|500373108|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|652157||4|0|45
502634923|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-16|2015-02-20|Followup|2014-08-16|2014-10-07|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|42.2||1|1|1|1|F|Black||13|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community||Match Support|F|Black||42|28210|Masters Degree|Single|Business: Clerical|28036|3|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|502635617|31|0|2|501197016|31|0|2|500548227|2||-2||4|1|||-2||-2|0|3|||46|2|||1|652158||4|1|45
503421607|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-26|2017-02-28|Followup|2014-09-26|2014-12-11|Expired|Late||||||||2|2|1|1|2|4|2|||||||||3|3|3|2|1|4|2.67||||||4|3|3|3.33|||||||3|5|5|5|4.5||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|4|4||||2|2||||4|4||Green||Child: Family structure changed|41.1||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28214|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|F|Black||49|28273|Associate Degree|Single|Finance: Accountant|28273|7|0|Agency Sponsored|Special Event|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503423471|36|0|2|503520561|31|0|2|500711787|2||-2||4|1|||-2|500000294|-2|0|10|||16426|8|||1|652257|646424|4|0|45
503552498|BBBS of Greater Charlotte|Main Office|C|Active|2014-01-30|NaT|Baseline|2013-09-26|2014-01-30|Complete|Done|2|1|1|1|2|4|1.83|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|||37.5||1|1|1|1|F|Black||13|No|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi|Match Support|F|White||29|28210|Bachelors Degree|Single|Business: Marketing|28277|1|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503554371|31|0|2|503538554|1|0|2|500744965|2||-2||2|1||500000294|-2||-2|0|10|||7464|9|||1|652321|-1|4|3|44
503318447|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-27|2017-02-23|Followup|2014-09-27|2014-09-25|Complete|Done|4|1|4|1|4|4|3|3|1|3|1|4|3|2.5|20|3|4|4|4|4|4|3.83|3|4|4|2|4|3|3.33|15.02|4|4|4|4|3|4|4|3.67|8.99|4|5|3|5|4.25|4|5|3|5|4.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|3|3|1|1|1|200|2|2|2|2|0|4|4|4|4|0|Green||Agency: Challenges with program/partnership|40.9||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||47|28215|Bachelors Degree|Married|Finance: Banking|28269|13|6|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|503320281|31|0|1|503537303|31|0|1|500709889|2||-2||4|1|||-2||-2|0|10|||7458|9|||1|652942|631862|4|3|45
503575828|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-28|2014-12-17|Followup|2014-09-28|2014-10-28|Complete|Done|3|2|4|3|3|4|3.17|3|3|4|4|3|4|3.5|-9.43|3|3|4|4|3|3|3.33|4|4|4|3|2|4|3.5|-4.86|4|4|3|3.67|4|3|3|3.33|10.21|4|4|5|4|4.25|3|3|4|4|3.5|21.43|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|4|4|4|4|4|4|0|3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Moved|14.6||3|3|1|1|M|Hispanic||13|No|Mother|28206|One Parent: Female|Unknown||Yes|Spanish Radio|Media|General Community|PERL 2014-2016|Match Support|M|White||26|28203|Bachelors Degree|Single|Finance: Banking|28202|0|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|503577713|3|0|1|503576000|1|0|1|500713280|2||-2||4|1||500014681|-2|500000294|-2|7068|1|||7464|9|||1|653133|651809|4|3|45
501300101|BBBS of Greater Charlotte|Main Office|C|Completed|2008-08-14|2015-05-11|Followup|2014-08-14|2014-09-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|80.9||1|1|4|4|F|Black||19|Yes|GrandMother|28273|Grandparents|Unknown||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501300379|31|0|2|500346193|31|0|2|500281421|2||500003586||4|2|500000294|500000294|-2||-2|7294|13|||46|2|||1|653326||4|1|45
502421176|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-30|2017-03-09|Followup|2014-09-30|2014-12-15|Expired|Late||||||||3|3|3|2|3|2|2.67|||||||||2|2|4|2|4|4|3||||||4|4|4|4|||||||4|5|5|5|4.75||||||||||4|4|4|4|4|4|4|4||||||4|4|3|3.67|||||4|4|4||||1|1||||4|4||Green||Volunteer: Time constraint|41.3||2|2|1|1|F|Black||18|No|GrandMother|28214|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||26|28078|Masters Degree|Single|Education: Teacher|28212|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502421614|31|0|2|503497451|31|0|2|500710577|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|653432|244394|4|0|45
503524258|BBBS of Greater Charlotte|Main Office|C|Completed|2013-09-30|2016-01-26|Followup|2014-09-30|2014-10-14|Complete|Done|4|4|4|2|4|4|3.67|3|4|4|1|1|3|2.67|37.45|2|4|4|4|4|4|3.67|1|1|4|1|1|4|2|83.5|4|4|4|4|3|4|4|3.67|8.99|4|4|5|4|4.25|5|3|5|4|4.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|2|4|1|2.33|71.67|4|2|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Moved|27.9||1|1|3|3|F|Black||14|No|Mother|28217|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Black||34|28273|Bachelors Degree|Single|Retail: Mgt|28217|5|6|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|503526133|31|0|2|500497043|31|0|2|500713184|2||-2||4|1||500000294|-2||-2|34|2|||6247|12|||1|653567|651722|4|3|45
501234606|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-16|NaT|Followup|2014-09-16|2014-10-20|Complete|Done|3|2|4|1|3|4|2.83|||||||||2|3|3|2|2|3|2.5|||||||||3|2|3|2.67||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||2|2|2|2||||||4|4|4|||||2|2||||4|4||||Green|||101.9||1|1|1|1|F|Black||16|No|Mother|28216|Grandparents|Unknown||No|TV|Media|General Community||Match Support|F|Black||42|28212|Bachelors Degree|Single|Unknown|28202|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501234882|31|0|2|501233675|31|0|2|500287478|2||-2||2|1|||-2||-2|56|1|||7464|9|||1|653758||4|3|45
503016111|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-30|2017-02-23|Followup|2014-09-30|2014-10-28|Complete|Done|4|4|4|4|4|4|4|3|3|4|3|4|4|3.5|14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|4|4|5|5|4.5|5|5|5|4|4.75|-5.26|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|1|3.57|8.12|3|4|4|3.67|4|4|3|3.67|0|3|3|3|2|2|2|50|2|2|2|2|0|4|4|4|4|0|Red||Volunteer: Time constraint|52.8||1|1|1|1|M|Black||14|Yes|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|M|Black||32|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503013381|31|0|1|503135600|31|0|1|500636811|2||500003586||4|3||500000294|-2|500000294|-2|0|10|||7496|10|||1|653928|496032|4|3|45
502391396|BBBS of Greater Charlotte|Main Office|C|Active|2013-05-15|NaT|Followup|2014-05-15|2014-06-12|Complete|Done|3|4|4|4|3|||||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green|Cabarrus County||46||2|2|1|1|F|Black||12|Yes|Mother|28052|One Parent: Female|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|White||40|28052|Bachelors Degree|Single|Transport: Pilot||1|1|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502391834|31|0|2|503228398|1|0|2|500690843|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|10|||7464|9|||1|654269||4|3|45
500784687|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-01|2016-01-05|Followup|2014-10-01|2014-10-27|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Red||Volunteer: Time constraint|27.1||2|2|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|No||Therapist/Counselor|General Community||Match Support|M|Black||32|28277|Bachelors Degree|Single|Construction|28211|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|500784955|31|0|1|503531111|31|0|1|500709609|2||-2||4|3|||-2||-2|0|5|||7464|9|||1|654325||4|3|45
501332658|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-01-19|Followup|2014-09-29|2014-10-31|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|4|3|4|1|4|3|||||||||4|4|4|4||||||4|4|4|||||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi|Child: Severity of challenges|87.7||1|1|1|1|M|Black||15|Yes|GrandMother|28213|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||46|28227|High School Graduate|Single|Medical: Healthcare Worker|28269|4|0|Coworker|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|277|60|598|500000170|500020752|501332937|31|0|1|501814288|1|0|1|500384166|2||-2||4|1|500000294|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||7447|3|||1|654328||4|3|45
501332660|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2015-04-08|Baseline|2013-10-02|2013-10-21|Complete|Done|3|4|4|4|3|1|3.17|||||||||2|4|3|2|2|4|2.83|||||||||4|3|4|3.67||||||4|4|2|5|3.75|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green||Volunteer: Moved|17.4||2|2|1|1|M|Black||13||GrandMother|28213|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||42|28212|Bachelors Degree|Married|Arts, Entertainment, Sports|28202|2|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|501332937|31|0|1|503579743|31|0|1|500715179|2||-2||4|1||500000294|-2||-2|6854|8|||7464|9|||1|654823|-1|4|3|44
503052850|BBBS of Greater Charlotte|Main Office|C|Active|2012-09-30|NaT|Followup|2014-09-30|2014-11-17|Declined|Late||||||||4|1|2|1|2|3|2.17|||||||||2|2|2|2|1|3|2||||||2|3|1|2|||||||3|4|2|3|3||||||||||4|4|4|4|4|3|4|3.86||||||4|4|4|4|||||3|3|3||||2|2||||4|4||Green|||53.5||1|1|1|1|F|Hispanic||13|No|Mother|28277|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||31|28210|Bachelors Degree|Single|Education: Teacher|29710|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020753|503027860|3|0|2|503028888|1|0|2|500626321|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|655087|476823|4|1|45
503470435|BBBS of Greater Charlotte|Main Office|C|Completed|2014-03-31|2014-06-30|Baseline|2013-10-03|2014-03-31|Complete|Done|3|4|3|2|3|4|3.17|||||||||1|3|3|2|1|3|2.17|||||||||3|2|2|2.33||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|1|2.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|3||1|1|1|1|M|White||14|No|Mother|28214|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||40|28205|Bachelors Degree|Separated|Construction|28205|4|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503472301|1|0|1|503597172|1|0|1|500757513|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|655446|-1|4|3|44
503580303|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-15|2014-06-18|Baseline|2013-10-03|2013-10-15|Complete|Done|4||4||4|4||||||||||4|4|3|3|2|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|8.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|M|White||42|28212|Bachelors Degree|Single|Business: Engineer||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503582180|31|0|1|503487684|1|0|1|500715761|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|655448|-1|4|3|44
502255210|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-27|NaT|Followup|2014-09-27|2014-10-22|Complete|Done|3|4|4|2|1|2|2.67|||||||||3|4|4|2|3|3|3.17|||||||||4|4|4|4||||||4|3|1|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||77.6||1|1|1|1|M|Black||14|No|Mother|28214|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||29|28210|Bachelors Degree|Married|Business: Mgt, Admin|97224|6|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|500910307|31|0|1|502255794|1|0|1|500470233|2||-2||2|1|||-2|500000294|-2|0|10|||7496|10|||1|655490||4|3|45
501641337|BBBS of Greater Charlotte|Main Office|C|Completed|2009-08-07|2015-03-13|Followup|2014-08-07|2014-10-22|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Moved|67.2||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||31|28269|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500011349|501641648|31|0|2|500835981|31|0|2|500373972|2||-2||4|1||500000294|-2|500000294|-2|0|10|||46|2|||1|655497||4|0|45
501597228|BBBS of Greater Charlotte|Main Office|C|Active|2009-09-04|NaT|Followup|2014-09-04|2014-09-08|Complete|Done|2|1|4|4|4|4|3.17|||||||||4|4|1|4|4|4|3.5|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|Amachi||90.3||1|1|1|1|F|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||40|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28204|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501597548|31|0|2|501397328|31|0|2|500379964|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|655503||4|3|45
503556265|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-18|2014-07-31|Baseline|2013-10-04|2013-10-18|Complete|Done|2|4|4|1|4|4|3.17|||||||||1|3|4|4|4|3|3.17|||||||||4|4|4|4||||||3|5|3|5|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|9.4||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Enrollment|F|Black||42|28216|Bachelors Degree|Single|Business: Mgt, Admin|28210|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503558140|31|0|2|503498990|31|0|2|500715926|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|655734|-1|4|3|44
500399844|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-20|2017-02-24|Followup|2014-08-20|2014-09-23|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Child: Graduated|114.2||1|2|1|2|F|Black||16||Mother|28208|One Parent: Female|Unknown||No||School|General Site||Match Support|F|White||35|28210|Bachelors Degree|Single|Business: Mgt, Admin|29715|0|0|Radio|Media|Big|General Site||Match Support|277|60|598|500000170|500008321|500400094|31|0|2|500188569|1|0|2|500190707|2||-2||4|3|||-1||-1|0|4|||131|1|||1|655992||4|3|45
502445356|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-04|2016-06-20|Followup|2014-10-04|2014-10-31|Complete|Done|4|1|4|1|4|4|3|4|1|3|4|4|4|3.33|-9.91|1|4|4|1|1|4|2.5|4|4|4|4|4|4|4|-37.5|4|4|4|4|4|4|4|4|0|4|4|4|4|4|5|4|3|3|3.75|6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|3|3.67|8.99|3|3|3|3|3|3|0|2|2|2|2|0|4|4||||Green||Child: Lost interest|44.5||1|2|4|5|F|Black||16|Yes|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community|Amachi|Match Support|F|Black||52|28216|Some College|Divorced|Business: Clerical|28202|16|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|502445803|31|0|2|501026290|31|0|2|500641693|2||-2||4|1||500000294|-2||-2|0|4|||46|2|||1|656238|244170|4|3|45
502236953|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-17|2015-01-30|Followup|2014-08-17|2014-09-22|Complete|Done|3|2|4|4|4|4|3.5|||||||||2|3|4|2|4|1|2.67|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Red||Volunteer: Time constraint|53.5||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Black||50|28212|Some College|Married|Law: Police Officer||2|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502237384|31|0|1|502232559|31|0|1|500464143|2||-2||4|3|||-2|500000294|-2|0|10|||7464|9|||1|656242||4|3|45
502290745|BBBS of Greater Charlotte|Main Office|C|Active|2012-04-26|NaT|Followup|2014-04-26|2014-06-09|Complete|Done|3|2|3|2|1|2|2.17|||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||2|5|2|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|||58.6||1|2|2|3|M|Black||12|No|Mother|28215|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||52|28207||Married|Medical: Doctor, Provider||0|0|Omega Psi Phi|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500020752|502291177|31|0|1|501944716|31|0|1|500611964|2||-2||2|1|||-2||-2|34|2|||8694|14|||1|656795||4|3|45
503533026|BBBS of Greater Charlotte|Main Office|C|Active|2013-10-19|NaT|Baseline|2013-10-09|2013-10-18|Complete|Done|1|3|4|2|3|2|2.5|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||5|4|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||40.9||1|1|2|2|F|Black||17|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|503534897|31|0|2|502485670|31|0|2|500717656|2||-2||2|1|||-2||-2|0|10|||7462|13|1204|3|1|657756|-1|4|3|44
502064627|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-20|NaT|Followup|2014-08-20|2014-08-18|Complete|Done|3|3|4|2|3|4|3.17|2|2|4|2|3|4|2.83|12.01|2|3|3|3|2|3|2.67|3|3|4|3|2|4|3.17|-15.77|4|3|4|3.67|4|3|2|3|22.33|4|4|2|3|3.25|5|3|3|4|3.75|-13.33|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|3|2|3|2.67|37.45|3|3|3|2|3|2.5|20|2|2|1|1|100|4|4||||Green|||78.9||1|1|2|2|M|Black||16|No|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|502065051|31|0|1|500773055|3|14|1|500462574|2||-2||2|1|||-2||-2|0|10|||46|2|||1|658102|159373|4|3|45
502721278|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-12|NaT|Followup|2014-10-12|2014-11-06|Complete|Done|3|4|4|4|4|4|3.83|||||||||1|4|4|4|4|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|1|3.57||||||||||3|4|3|3.33||||||1|3|2|||||2|2||||4|4||||Green|Amachi, Cabarrus County||65.1||1|1|1|1|M|White||13|Yes|Mother|28025|One Parent: Female|Unknown||Yes||School|General Community|Cabarrus County|Match Support|M|White||47|28025||Single|Tech: Support, Writing|28026|0|2|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501938680|1|0|1|502701096|1|0|1|500560499|2||500003586||2|1|500000294, 500016374|500016374|-2|500016374|-2|0|4|||7464|9|||1|658109||4|3|45
502471024|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-09|2016-08-01|Followup|2014-09-09|2014-09-12|Complete|Done|4|3|1|2|4|4|3|||||||||3|4|3|3|4|4|3.5|||||||||4|4|4|4||||||5|5|3|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Feels incompatible with child/family|58.7|Y|1|1|1|1|M|Black||13|Yes|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||51|28205|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502471471|31|0|1|502685747|1|0|1|500552890|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|658457||4|3|45
503587461|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-30|2015-06-17|Baseline|2013-10-11|2013-10-30|Complete|Done|3|2|3|2|3|4|2.83|||||||||4|4|3|2|2|4|3.17|||||||||4|4|4|4||||||5|4|2|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||1|1||||4|4||||Green||Child/Family: Time constraints|19.5||1|1|1|1|F|Black||14|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Finance|28202|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503587387|31|0|2|503541106|1|0|2|500718377|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|658777|-1|4|3|44
502172536|BBBS of Greater Charlotte|Main Office|C|Active|2010-10-13|NaT|Followup|2014-10-13|2014-10-20|Complete|Done|2|4|4|4|4|4|3.67|3|2|4|3|1|1|2.33|57.51|3|4|4|3|3|4|3.5|2|4|4|2|2|4|3|16.67|4|4|4|4|4|4|4|4|0|3|4|5|5|4.25|5|4|4|4|4.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|3|4|4|3.67|-18.26|3|3|3|4|2|3|0|2|2|2|2|0|4|4||||Green|||77.1||1|1|1|1|F|Black||17|No|Mother|28269|Two Parent|Unknown||Yes||Relative|General Community||Match Support|F|Multi-race (Asian & White)||33|28205|Masters Degree|Married|Finance: Economist|28223|7|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|502172965|31|0|2|501279665|37|0|2|500475431|2||-2||2|1|||-2||-2|0|3|||129|1|||1|659194|184611|4|3|45
502097843|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-29|2016-08-11|Followup|2014-08-29|2014-08-25|Complete|Done|3|4|4|4|3|3|3.5|3|2|2|1|4|3|2.5|40|4|4|4|4|4|4|4|2|3|3|2|3|3|2.67|49.81|4|4|4|4|4|4|4|4|0|3|5|5|5|4.5|3|3|3|4|3.25|38.46|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|3|3|3|33.33|3|3|3|3||||2|2|2|2|0|4|4|4|4|0|Green|2010-2012 OJJDP JJI|Child: Lost interest|59.4||1|1|2|2|M|Black||17|No|Mother|28078|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500021785|502098263|31|0|1|502643791|3|0|1|500550390|2||-2||4|1|500005291||-2||-2|0|10|||7496|10|||1|659429|330290|4|3|45
503590328|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-27|2016-09-28|Baseline|2013-10-14|2014-08-27|Complete|Done|3|2|4|1|4|4|3|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|25.1||1|1|1|1|M|Hispanic||12|No|Mother|28277|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|Some Other Race||31|28270|Bachelors Degree|Married|Real Estate: Realtor|28110|0|5|Man Up Campaign|Media|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|277|60|598|500000170|500008321|503592205|3|0|1|503874645|41|0|1|500771736|2||-2||4|3|||-2|500011312|-2|0|10|||17101|1|||1|659454|-1|4|3|44
503506115|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-23|2016-09-27|Baseline|2013-10-14|2013-10-23|Complete|Done|3|1|3|1|3|2|2.17|||||||||2|3|2|4|1|3|2.5|||||||||3|4|3|3.33||||||2|4|3|5|3.5|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|3|3.67||||||1|4|2.5|||||2|2||||4|4||||Red||Child: Family structure changed|35.2||1|1|1|1|M|Black||13|No|Mother|28215|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Asian||54|28211|Masters Degree|Married|Self-Employed, Entrepreneur|28211|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503507986|31|0|1|503552068|4|0|1|500718774|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|659462|-1|4|3|44
503490571|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-20|2015-05-14|Baseline|2013-10-14|2013-12-19|Complete|Done|3|4|4|3|3|3|3.33|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|3|4|4|4|4|4|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|VOL - Mentoring Hispanic Youth|Child/Family: Lost contact with volunteer/agency|16.8||1|1|1|1|F|Hispanic|Mexican|16|No|Mother|28208|Two Parent|Unknown|Y|Yes|Spanish Radio|Media|General Community||Match Support|F|White||35|28214|Bachelors Degree|Single|Transport: Flight Attendant|85034|0|3|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|503492439|3|10|2|503645850|1|0|2|500738556|2||-2||4|3|500011312||-2|500000294|-2|7068|1|||7464|9|||1|659479|-1|4|3|44
503533022|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2015-03-03|Baseline|2013-10-14|2013-10-18|Complete|Done|4|2|3|3|4|3|3.17|||||||||4|4|4|3|4|3|3.67|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|4|3|||||1|1||||4|4||||Green||Volunteer: Moved|16.3||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||RTBM|M|Black||27|28216|Bachelors Degree|Single|Business: Engineer|28202|0|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503534897|31|0|1|503534544|31|0|1|500718872|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|659547|-1|4|3|44
501529924|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-27|2017-02-28|Followup|2014-08-27|2014-08-27|Complete|Done|3|4|4|3|4|4|3.67|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|78.1||2|2|1|1|F|Black||15|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||30|28209|Bachelors Degree|Single|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|501530213|31|0|2|502199360|1|0|2|500465517|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|660631||4|3|45
503425736|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-16|2016-06-15|Followup|2014-10-16|2014-10-20|Complete|Done|3|3|4|3|3|3|3.17|3|3|4|2|4|4|3.33|-4.8|3|4|4|3|2|3|3.17|3|4|3|3|3|3|3.17|0|4|4|4|4|4|4|4|4|0|4|5|4|3|4|4|3|2|3|3|33.33|4|3|4|4|3|4|3|3.57|2|2|2|2|2|2|2|2|78.5|2|1|1|1.33|1|2|2|1.67|-20.36|3|2|2.5|4|2|3|-16.67|2|2|1|1|100|4|4|4|4|0|Green||Child: Graduated|32||1|1|1|1|F|Black||18|No|GrandMother|28213|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|White||29|28211|Juris Doctorate (JD)|Married|Law|28202|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|503427601|31|0|2|503519747|1|0|2|500711543|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|660783|649102|4|3|45
502436202|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-02|2015-07-13|Followup|2014-09-02|2014-11-17|Expired|Late||||||||3|2|2|1|3|3|2.33|||||||||3|3|3|4|2|4|3.17||||||4|4|4|4|||||||2|5|5|5|4.25||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||2|4|3||||1|1||||4|4||Green||Child: Graduated|46.3||1|1|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|Masters Degree|Single|Finance: Banking||0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|502436645|31|0|1|502642999|1|0|1|500549046|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|661151|327937|4|0|45
502034298|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-19|2015-08-31|Followup|2014-10-19|2014-12-06|Declined|Late||||||||3|4|4|2|4|4|3.5|||||||||2|4|3|4|3|4|3.33||||||4|4|4|4|||||||5|5|5|4|4.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||2|4|3||||1|1|||||||Red||Volunteer: Time constraint|34.4||2|3|4|6|M|White||16|Yes|Mother|28146|One Parent: Female|Unknown||Yes||School|General Community|Amachi|Match Support|M|White||41|28078|Bachelors Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502034697|1|0|1|500188638|1|0|1|500631278|2||-2||4|3||500000294|-2|500000294|-2|0|4|||7464|9|||1|661714|27853|4|1|45
503523387|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-29|2014-11-21|Baseline|2013-10-18|2013-10-29|Complete|Done|3|1|2|1|3|3|2.17|||||||||2|4|4|2|2|3|2.83|||||||||4|4|4|4||||||4|3|4|5|4|||||||4|4|4|4|4|4|2|3.71||||||||||2|4|4|3.33||||||3|4|3.5|||||2|2||||4|4||||Green||Child/Family: Moved|12.7||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||29|28262|Juris Doctorate (JD)|Single|Law: Lawyer||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|503525262|31|0|2|503537943|31|0|2|500720846|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|661917|-1|4|3|44
501314348|BBBS of Greater Charlotte|Main Office|C|Completed|2010-08-25|2015-07-31|Followup|2014-08-25|2014-11-09|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Volunteer: Lost contact with child/agency|59.2||1|1|1|1|M|Black||12|No|Mother|28210|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||45|28211|Masters Degree|Married|Finance: Banking||11|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500008321|501314626|31|0|1|502205797|1|0|1|500460633|2||-2||4|3|||-2||-2|0|10|||2230|7|||1|662145||4|0|45
500474486|BBBS of Greater Charlotte|Main Office|C|Completed|2006-08-23|2015-08-18|Followup|2014-08-23|2014-11-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|107.8||1|1|1|1|M|Black||20||Mother|28214|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||38|28209|Bachelors Degree|Single|Construction|28247|0|2|Coworker|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500474735|31|0|1|500491064|31|0|1|500118168|2||-2||4|3|||-2||-2|34|2|||7447|3|||1|662147||4|0|45
503533026|BBBS of Greater Charlotte|Main Office|C|Active|2013-10-19|NaT|Followup|2014-10-19|2014-12-23|Declined|Late||||||||1|3|4|2|3|2|2.5|||||||||3|4|4|3|4|4|3.67||||||4|4|4|4|||||||5|4|3|4|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||3|3|3||||1|1||||4|4||Green|||40.9||1|1|2|2|F|Black||17|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|503534897|31|0|2|502485670|31|0|2|500717656|2||-2||2|1|||-2||-2|0|10|||7462|13|1204|3|1|662348|657756|4|1|45
501253195|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-24|NaT|Followup|2014-10-24|2014-10-24|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|4|4|2|2|3|3.17|||||||||4|4|4|4||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|Amachi||100.7||1|1|2|2|M|Black||15|Yes|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||37|28203|Masters Degree|Single|Medical: Doctor, Provider|28211|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|501253471|31|0|1|500395148|1|0|1|500282924|2||500003586||2|1|500000294||-2||-2|0|10|||7464|9|||1|662456||4|3|45
501254255|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-23|2017-02-28|Followup|2014-09-23|2014-10-20|Complete|Done|4|4|4|4|3|4|3.83|||||||||4|4|4|2|4|3|3.5|||||||||4|3|4|3.67||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|3|2|||||2|2||||4|4||||Green||Volunteer: Moved|101.2||1|1|1|1|F|Black||14|No|Mother|28230|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||34|28205|Masters Degree|Single|Finance: Banking|28217|0|4|Yahoo!|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|501254531|31|0|2|501356688|1|0|2|500282157|2||-2||4|1|||-2|500000294|-2|0|10|||32|2|||1|662457||4|3|45
500185723|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-05|2015-06-25|Followup|2014-09-05|2014-11-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child: Graduated|81.6||2|2|1|1|M|Black||19||Mother|28214|One Parent: Female|Unknown||No|AARTF|Neighbor/Friend|General Community||Match Support|M|Black||36|28214|Bachelors Degree|Single|Tech: Computer/Programmer|28147|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187335|31|0|1|501310677|31|0|1|500284133|2||-2||4|3|||-2||-2|6855|8|||7464|9|||1|662474||4|1|45
501010684|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-22|2017-02-23|Followup|2014-10-22|2014-10-20|Complete|Done|1|1|1|1|4|1|1.5|4|2|1|3|3|1|2.33|-35.62|1|4|3|4|1|4|2.83|1|2|3|1|3|1|1.83|54.64|4|4|4|4|4|4|4|4|0|5|3|4|4|4|4|5|3|3|3.75|6.67|4|4|4|4|4|4|4|4|1|4|4|3|4|4|3|3.29|21.58|4|4|3|3.67|3|4|2|3|22.33|3|3|3|1|2|1.5|100|2|2|1|1|100|4|4|4|4|0|Green||Volunteer: Time constraint|40.1||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Less than $10,000||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|White||41|28269|Bachelors Degree|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503560069|31|0|1|503491643|1|0|1|500710107|2||-2||4|1||500005291|-2||-2|7016|11|||7464|9|||1|663317|327911|4|3|45
503398288|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-31|2014-12-23|Followup|2014-08-31|2014-11-15|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Moved|15.7||1|1|1|1|M|Hispanic|Mexican|12|No|Mother|28206|One Parent: Female|$15,000 to $19,999|Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||28|28202|Masters Degree|Single|Consultant||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|503400145|3|10|1|503473834|1|0|1|500707156|2||-2||4|2|||-2|500000294|-2|0|5|||7496|10|||1|663837||4|0|45
503506115|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-23|2016-09-27|Followup|2014-10-23|2014-12-05|Complete|Done|3|2|3|3|3|3|2.83|3|1|3|1|3|2|2.17|30.41|3|3|3|3|3|3|3|2|3|2|4|1|3|2.5|20|3|3|3|3|3|4|3|3.33|-9.91|2|3|3|3|2.75|2|4|3|5|3.5|-21.43|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3|3.71|7.82|4|4|4|4|4|4|3|3.67|8.99|3|3|3|1|4|2.5|20|2|2|2|2|0|4|4|4|4|0|Red||Child: Family structure changed|35.2||1|1|1|1|M|Black||13|No|Mother|28215|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Asian||54|28211|Masters Degree|Married|Self-Employed, Entrepreneur|28211|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503507986|31|0|1|503552068|4|0|1|500718774|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|664460|659462|4|3|45
501309634|BBBS of Greater Charlotte|Main Office|C|Active|2008-09-12|NaT|Followup|2014-09-12|2014-09-19|Complete|Done|3|4|3|2|3|3|3|||||||||3|4|3|2|3|3|3|||||||||4|4|4|4||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|Amachi||102.1||1|1|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Match Support|F|Black||46|27704|Associate Degree|Divorced|Medical: Admin||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|501309912|31|0|2|501046221|31|0|2|500281317|2||500003586||2|1|500000294|500000294|-2|500000294|-2|0|10|||7462|13|||1|664846||4|3|45
502129650|BBBS of Greater Charlotte|Main Office|C|Active|2012-10-26|NaT|Followup|2014-10-26|2014-10-27|Complete|Done|4|3|4|4|3|4|3.67|4|4|4|4|4|4|4|-8.25|3|3|4|4|3|4|3.5|1|4|3|4|1|4|2.83|23.67|4|4|4|4|4|4|4|4|0|5|5|4|5|4.75|5|4|5|4|4.5|5.56|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|2|2|4|4|4|-50|2|2|2|2|0|4|4||||Green|Cabarrus County||52.6||2|2|2|2|F|Black||17|No|GrandMother|28027|Grandparents|Unknown||No||Self|General Community|Cabarrus County|Match Support|F|Black||42|28213|Bachelors Degree|Single|Finance: Banking|28202|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502130079|31|0|2|502598777|31|0|2|500646243|2||500016307||2|1|500016374|500016374|-2|500016374|-2|0|10|||7464|9|||1|664871|220242|4|3|45
501332660|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2015-04-08|Followup|2014-10-24|2014-10-28|Complete|Done|3|1|4|1|4|4|2.83|3|4|4|4|3|1|3.17|-10.73|4|4|4|1|4|4|3.5|2|4|3|2|2|4|2.83|23.67|4|3|4|3.67|4|3|4|3.67|0|3||3|4||4|4|2|5|3.75||4|4|4|4|4|4|4|4|4|4|4|4|3|4|4|3.86|3.63|1|4|4|3|4|4|4|4|-25|4|4|4|4|2|3|33.33|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|17.4||2|2|1|1|M|Black||13||GrandMother|28213|Grandparents|Unknown||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||42|28212|Bachelors Degree|Married|Arts, Entertainment, Sports|28202|2|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500011349|501332937|31|0|1|503579743|31|0|1|500715179|2||-2||4|1||500000294|-2||-2|6854|8|||7464|9|||1|664930|654823|4|3|45
503492220|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2015-10-20|Baseline|2013-10-24|2013-10-24|Complete|Done|3|1|3|2|4|4|2.83|||||||||2|3|3|2|2|4|2.67|||||||||4|4|4|4||||||2|4|1|2|2.25|||||||4|4|4|4|3|4|2|3.57||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|23.9||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||27|28205|Bachelors Degree|Single|Business: Clerical|28277|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503494082|31|0|2|503521240|1|0|2|500711792|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|665105|-1|4|3|44
503492220|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2015-10-20|Followup|2014-10-24|2015-01-08|Expired|Late||||||||3|1|3|2|4|4|2.83|||||||||2|3|3|2|2|4|2.67||||||4|4|4|4|||||||2|4|1|2|2.25||||||||||4|4|4|4|3|4|2|3.57||||||3|4|3|3.33|||||4|4|4||||2|2||||4|4||Yellow||Child/Family: Lost contact with volunteer/agency|23.9||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||27|28205|Bachelors Degree|Single|Business: Clerical|28277|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503494082|31|0|2|503521240|1|0|2|500711792|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|665108|665105|4|0|45
503533022|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2015-03-03|Followup|2014-10-24|2014-12-23|Declined|Late||||||||4|2|3|3|4|3|3.17|||||||||4|4|4|3|4|3|3.67||||||4|4|4|4|||||||5|5|4|4|4.5||||||||||4|4|4|4|4|4|3|3.86||||||3|4|3|3.33|||||2|4|3||||1|1||||4|4||Green||Volunteer: Moved|16.3||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||RTBM|M|Black||27|28216|Bachelors Degree|Single|Business: Engineer|28202|0|1|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503534897|31|0|1|503534544|31|0|1|500718872|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|665113|659547|4|1|45
502969236|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-24|2015-07-23|Followup|2014-10-24|2014-10-27|Complete|Done|3|2|2|2|4|3|2.67|||||||||1|1|4|1|2|3|2|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|20.9||2|2|1|1|F|Some Other Race||13||Mother|28277|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||30|29730|Bachelors Degree|Single|Finance: Accountant|28273|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502970672|41|0|2|503567563|1|0|2|500718760|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|665398||4|3|45
503530345|BBBS of Greater Charlotte|Main Office|C|Completed|2013-08-13|2016-11-07|Followup|2014-08-13|2014-08-13|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|1|2|4|2.83|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|2|2|||||2|2||||4|4||||Red|Cabarrus County|Volunteer: Lost contact with child/agency|38.8||1|1|2|2|F|Black||12|No|Mother|28025|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County|RTBM|F|Black||43|28027|Masters Degree||Education: Teacher|28027|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501204816|31|0|2|502460114|31|0|2|500704946|2||500016307||4|3|500016374|500016374|-2|500016374|-2|0|10|||7464|9|||1|665594||4|3|45
502763586|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-06|2017-02-28|Followup|2014-09-06|2014-09-02|Complete|Done|4|1|1|1|2|2|1.83|3|2|3|2|4|3|2.83|-35.34|3|4|4|3|3|4|3.5|2|3|2|2|2|3|2.33|50.21|4|4|4|4|4|4|4|4|0|5|5|5|5|5|3|3|2|2|2.5|100|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|2|2|2|2|100|1|4|2.5|3|3|3|-16.67|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Moved|53.7||1|2|5|6|M|Black||16||Mother|28208|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Black|Other African|53|28277||Married|Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502764498|31|0|1|500189754|31|31|1|500632648|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|667290|358930|4|3|45
502551048|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-19|2015-01-15|Followup|2014-10-19|2014-10-30|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|3|2|1|2|3|2.17|||||||||4|3|4|3.67||||||4|5|5|3|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Yellow||Volunteer: Moved|38.9||1|1|2|2|F|Hispanic||13|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Enrollment|F|Black||52|30080|Bachelors Degree|Single|Consultant|2451|3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502551498|3|0|2|501472128|31|0|2|500554178|2||-2||4|2|||-2||-2|0|4|||7464|9|||1|667306||4|3|45
503523387|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-29|2014-11-21|Followup|2014-10-29|2014-10-30|Complete|Done|3|3|4|3|4|4|3.5|3|1|2|1|3|3|2.17|61.29|2|4|3|3|3|3|3|2|4|4|2|2|3|2.83|6.01|4|4|4|4|4|4|4|4|0|2|5|2|3|3|4|3|4|5|4|-25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|2|3.71|4.04|2|2|2|2|2|4|4|3.33|-39.94|3|3|3|3|4|3.5|-14.29|2|2|2|2|0|4|4|4|4|0|Green||Child/Family: Moved|12.7||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||29|28262|Juris Doctorate (JD)|Single|Law: Lawyer||0|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|503525262|31|0|2|503537943|31|0|2|500720846|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|667340|661917|4|3|45
502374716|BBBS of Greater Charlotte|Main Office|C|Active|2013-10-29|NaT|Followup|2014-10-29|2014-12-29|Declined|Late|4|3|3|2|4|4|3.33|4|4|4|3|2|3|3.33|0|2|4|3|3|2|4|3|2|3|3|2|2|3|2.5|20|4|2|3|3|4|4|4|4|-25|3|3|3|4|3.25|3|3|4|3|3.25|0|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|4|4|3.67|-9.26|2|3|2.5|4|4|4|-37.5|2|2|2|2|0|4|4||||Green|||40.5||2|2|1|1|M|Hispanic|Mexican|16|No|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Hispanic||29|28214|Bachelors Degree|Single|Self-Employed, Entrepreneur|28214|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020753|502375154|3|10|1|503560077|3|0|1|500723012|2||-2||2|1|||-2||-2|0|4|||46|2|||1|667945|199086|4|1|45
503587461|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-30|2015-06-17|Followup|2014-10-30|2015-01-03|Declined|Late||||||||3|2|3|2|3|4|2.83|||||||||4|4|3|2|2|4|3.17||||||4|4|4|4|||||||5|4|2|3|3.5||||||||||4|4|4|4|4|4|4|4||||||3|4|4|3.67|||||3|3|3||||1|1||||4|4||Green||Child/Family: Time constraints|19.5||1|1|1|1|F|Black||14|Yes|Mother|28262|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Finance|28202|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503587387|31|0|2|503541106|1|0|2|500718377|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|668957|658777|4|1|45
500186106|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-18|2015-08-13|Followup|2014-10-18|2014-12-11|Complete|Late|3|2|4|4|3|3|3.17|||||||||4|4|3|3|3|3|3.33|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|93.8||2|2|1|1|F|Black||20||Mother|28217|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||35|28211|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|500187698|31|0|2|500778380|1|0|2|500202993|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|670186||4|3|45
502223076|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-21|NaT|Followup|2014-10-21|2014-10-29|Complete|Done|3|2|3|3|3|3|2.83|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|||64.8||2|2|1|1|F|Black||12|No|Mother|28216|One Parent: Female|Unknown||Yes||Self|General Community|Project Big|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Mgt, Admin|28204|0|9|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|502223507|31|0|2|502694717|1|0|2|500560829|2||-2||2|1||500004640|-2||-2|0|10|||7464|9|||1|670188||4|3|45
502205848|BBBS of Greater Charlotte|Main Office|C|Active|2011-08-18|NaT|Followup|2014-08-18|2014-09-02|Complete|Done|4|1|4|3|4|4|3.33|3|4|3|2|4|4|3.33|0|2|4|3|2|2|4|2.83|3|2|3|4|3|3|3|-5.67|4|4|4|4|4|4|4|4|0|3||2|2||4|4|5|4|4.25||4|4|4|4|4|4|4|4|4|4|4|4|3|4|4|3.86|3.63|4|4|4|4|4|4|3|3.67|8.99|2|1|1.5|2|4|3|-50|2|2|1|1|100|4|4|4|4|0|Green|2010-2012 OJJDP JJI||66.9||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Juris Doctorate (JD)|Single|Student: College|28208|0|0||Law Student Association|Big|General Community||Match Support|277|60|598|500000170|500020753|502206277|31|0|1|502624702|1|0|1|500549350|2||-2||2|1|500005291|500005291|-2||-2|0|10|||0|15|||1|670530|328511|4|3|45
501725162|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-29|2016-10-14|Followup|2014-10-29|2014-12-29|Declined|Late||||||||4|1|2|1|4|4|2.67|||||||||3|4|2|3|3|3|3||||||1|4|4|3|||||||5|1|5|5|4||||||||||4|4|4|4|4|4|3|3.86||||||4|4|2|3.33|||||4|3|3.5||||2|2|||||||Green||Agency: Challenges with program/partnership|83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501724831|39|0|1|501833178|1|0|1|500394157|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|670982|16143|4|1|45
500382177|BBBS of Greater Charlotte|Main Office|C|Completed|2006-09-18|2015-08-25|Followup|2014-09-18|2014-09-18|Complete|Done|4|4|4|4|4|3|3.83|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|107.2||1|1|2|2|M|Black||16||Mother|28215|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||43|28215|Bachelors Degree|Single|Finance: Banking|28262|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500012459|500382427|31|0|1|500188566|31|0|1|500122093|2||-2||4|2|||-2||-2|0|10|||7496|10|||1|671018||4|3|45
503643026|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-26|2014-03-13|Baseline|2013-11-04|2013-11-26|Complete|Done|3|1|2|1|1|2|1.67|||||||||3|4|4|2|2|4|3.17|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|1|1.5|||||1|1||||4|4||||Yellow||Volunteer: Time constraint|3.5||3|3|1|1|F|Black||14|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Business: Human Resources||1|3|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500015820|503644986|31|0|2|503603792|1|0|2|500731516|2||-2||4|2|||-2||-2|0|10|||7671|13|||1|671048|-1|4|3|44
503666553|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-13|2014-10-30|Baseline|2013-11-04|2013-12-13|Complete|Done|4|1|4|1|4|4|3|||||||||2|4|1|2|2|4|2.5|||||||||4|3|4|3.67||||||3|4|5|5|4.25|||||||4|1|4|4|3|4|4|3.43||||||||||4|3|2|3||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|10.5||2|2|1|1|F|Black||13|Yes|Mother|28025|One Parent: Female|$75,000 to $99,999||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||54|28056|PHD|Married|Education: College Professor|28017|4|0|Newspaper|Media|Big|General Community||Match Support|277|60|598|500000170|500015820|503668509|31|0|2|503548907|31|0|2|500727074|2||-2||4|1||500014681, 500016374|-2||-2|0|10|||129|1|||1|671051|-1|4|3|44
503041998|BBBS of Greater Charlotte|Main Office|C|Active|2012-10-16|NaT|Followup|2014-10-16|2014-12-06|Declined|Late||||||||4|2|3|2|3|4|3|||||||||2|3|3|1|2|4|2.5||||||3|4|4|3.67|||||||4|3|5|3|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||2|4|3||||2|2||||4|4||Yellow|||53||1|1|1|1|M|Black||15|No|Mother|28214|One Parent: Female|$45,000 to $49,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28207|Masters Degree|Married|Finance|28273|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503043639|31|0|1|503110820|1|0|1|500638908|2||-2||2|2|||-2||-2|34|2|||7464|9|||1|671300|498892|4|1|45
500826594|BBBS of Greater Charlotte|Main Office|C|Completed|2007-08-21|2016-06-15|Followup|2014-08-21|2014-11-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|105.8||1|1|1|1|M|Black||18|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|M|Some Other Race||36|28209|||Business: Sales||0|0|General|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|1|500920342|41|0|1|500185735|2||-2||4|1|||-2||-2|0|5|||6450|12|||1|671340||4|0|45
502875668|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-31|2015-07-31|Followup|2014-10-31|2014-12-15|Complete|Done|2|2|3|3|3|3|2.67|||||||||2|3|3|2|3|||||||||||3|3|3|3||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3||||||||||4|4||||Red||Volunteer: Time constraint|33||1|1|1|1|M|Black||12|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Asian||39|28262|PHD|Married|Business: Mgt, Admin|28202|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502877071|31|0|1|503114677|4|0|1|500649397|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|672943||4|3|45
502499851|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-11|2015-07-07|Followup|2014-11-11|2014-11-24|Complete|Done|3|3|3|3|3|3|3|3|1|1|1|2|2|1.67|79.64|2|4|3|3|3|3|3|4|4|4|2|2|4|3.33|-9.91|4|4|4|4|4|4|4|4|0|2|3|4|3|3|5|5|5|4|4.75|-36.84|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|4|3.33|3|4|3|3.33|0|2|4|3|2|4|3|0|2|2|2|2|0|4|4|4|4|0|Red||Agency: Concern with Volunteer re: child safety|43.8||1|1|1|1|M|White||18|No|Mother|28210|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|White||39|28210|Masters Degree|Single|Finance|28106|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|502500300|1|0|1|502690262|1|0|1|500562789|2||-2||4|3|||-2||-2|0|10|||46|2|||1|674719|348364|4|3|45
502206673|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-13|2015-06-23|Followup|2014-10-13|2014-10-28|Complete|Done|3|4|4|2|4|4|3.5|3|2|3|2|3|4|2.83|23.67|2|4|4|2|2|3|2.83|2|3|3|3|3|3|2.83|0|4|4|4|4|4|4|4|4|0|3|3|4|3|3.25|4|5|3|3|3.75|-13.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|3|4|4|3.67|8.99|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Red|Amachi|Child: Lost interest|44.3||1|1|1|1|M|Black||17|Yes|GrandMother|28216|Grandparents|Unknown||Yes||Self|General Community|Amachi|Match Support|M|White||47|28216|Bachelors Degree|Married|Business: Engineer|28255|18|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500013781|502207102|31|0|1|502668179|1|0|1|500557233|2||500003586||4|3|500000294|500000294|-2||-2|0|10|||7464|9|||1|674778|341305|4|3|45
501023408|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-05|NaT|Followup|2014-11-05|2014-11-19|Complete|Done|3|2|1|2|3|3|2.33|||||||||3|3|2|4|4|3|3.17|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Green|||100.3||1|1|1|1|M|Hispanic|Other South American|17|No|Mother|28273|One Parent: Female|Less than $10,000||Yes||Self|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|501023677|3|15|1|501356600|1|0|1|500296545|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|675067||4|3|45
503617980|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-25|2016-01-06|Baseline|2013-11-13|2013-11-25|Complete|Done|4|2|4|4|4|4|3.67|||||||||2|4|4|3|4|3|3.33|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||1|3|2|||||2|2||||4|4||||Green||Child/Family: Moved|25.4||1|1|1|1|F|Black||13|No|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|White||25|28134|Some College|Single|Child/Day Care Worker||0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503619857|31|0|2|503573243|1|0|2|500730441|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|675746|-1|4|3|44
503417576|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-09|2015-12-30|Baseline|2013-11-13|2013-12-09|Complete|Done|3|1|2|1|3|3|2.17||||||||||2|2|2|2|1||||||||||3|3|4|3.33||||||2|3|3|2|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|24.7||1|1|1|1|F|White||17|No|Father|28269|Two Parent|$100,000 to $124,999|Y|No||Relative|General Community||Match Support|F|White||29|28205|Some College|Single|Business: Mgt, Admin|29707|3|10|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503419440|1|0|2|503594017|1|0|2|500730510|2||-2||4|3|||-2|500000294|-2|0|3|||7464|9|||1|675823|-1|4|3|44
500545326|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2016-09-02|Followup|2014-10-29|2014-12-10|Complete|Done|4|4|4|4|4|4|4|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||4|1|4|4|3.25|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|118.1|Y|1|1|1|1|M|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|Y|No||Self|General Community||Match Support|M|Black||55|28214||Married|Clergy||12|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500545578|7|0|1|500697845|31|0|1|500134545|2||-2||4|3|||-2||-2|0|10|||2238|7|||1|676193||4|3|45
502987717|BBBS of Greater Charlotte|Main Office|C|Completed|2014-03-19|2015-03-26|Baseline|2013-11-14|2014-03-19|Complete|Done|3|3|2|3|2|3|2.67|||||||||2|3|2|2|2|3|2.33|||||||||4|1|1|2||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green||Child/Family: Moved|12.2||1|1|1|1|F|Black||13|No|Mother|28134|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|White||37|28209|Bachelors Degree|Divorced|Medical|28078|5|6|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|502989174|31|0|2|503559146|1|0|2|500753781|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|676731|-1|4|3|44
503701025|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-25|2016-08-18|Baseline|2013-11-15|2013-11-25|Complete|Done|4|1|4|1|3|4|2.83|||||||||1|1|1|1|1|4|1.5|||||||||4|4|4|4||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|32.8||1|1|1|1|F|Black||12|Yes|Mother|28269|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|White||53|28227|Some College|Married|Customer Service|28105|30|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|501153063|31|0|2|503576358|1|0|2|500731543|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|677325|-1|4|3|44
502485856|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-15|2015-10-13|Followup|2014-11-15|2014-12-08|Complete|Done|3|2|3|1|3|4|2.67|||||||||3|4|3|4|3|4|3.5|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|22.9||2|2|1|1|F|Hispanic|Other South American|13|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community||Enrollment|F|Hispanic||39|28278|Associate Degree|Married|Finance||1|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|502486303|3|15|2|503544124|3|0|2|500726848|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|677439||4|3|45
503597088|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-06|2016-05-03|Baseline|2013-11-15|2013-12-06|Complete|Done|4|1|4|2|4|4|3.17|||||||||3|4|3|2|4|4|3.33|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|4|3.67||||||1|2|1.5|||||2|2||||4|4||||Green||Volunteer: Moved|28.9||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Retail: Sales|28217|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503598965|31|0|2|503642924|1|0|2|500731612|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|677446|-1|4|3|44
502273093|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-01|2015-03-31|Followup|2014-10-01|2014-11-14|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|3|3|3.33||||||4|4|4|||||2|2||||4|4||||Green||Child/Family: Moved|53.9||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|Black||37|28277|PHD|Single|Medical: Healthcare Worker||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502273525|31|0|2|502252422|31|0|2|500471568|2||-2||4|1|||-2|500000294|-2|0|4|||7496|10|||1|677489||4|3|45
500970267|BBBS of Greater Charlotte|Main Office|C|Active|2010-09-29|NaT|Followup|2014-09-29|2014-12-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi||77.5||1|1|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||61|28204||Divorced|Self-Employed, Entrepreneur||0|0|Billboard|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|500970535|31|0|2|502084649|1|0|2|500468192|2||500003586||2|1|500000294|500000294|-2|500000294|-2|5635|9|||125|1|||1|677492|174196|4|1|45
501859854|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-29|2015-09-16|Followup|2014-09-29|2014-12-11|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|Amachi|Volunteer: Lost contact with child/agency|59.6||1|1|1|1|F|Black||13|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||28|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501860227|31|0|2|502044100|31|0|2|500469954|2||500003586||4|1|500000294|500000294|-2||-2|0|10|||7464|9|||1|677493||4|1|45
501237971|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-17|2016-03-03|Followup|2014-11-17|2014-11-21|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|39.5||2|2|3|3|F|Black||18|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|Y|Yes||Self|General Community|Amachi|Match Support|F|Black||41|28269|||Business: Human Resources|28206|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503287812|31|0|2|501598429|31|0|2|500649363|2||-2||4|1||500000294|-2||-2|0|10|||7464|9|||1|677714||4|3|45
501938282|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-17|NaT|Followup|2014-11-17|2014-11-17|Complete|Done|4|3|4|4|3|4|3.67|||||||||1|3|3|1|2|3|2.17|||||||||4|2|2|2.67||||||3|2|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||1|1|1|||||2|2||||4|4||||Green|Amachi, Cabarrus County||75.9||1|1|1|1|F|White||14|Yes|Mother|28025|Two Parent|Unknown|Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||63|28027|High School Graduate|Married|Self-Employed, Entrepreneur|28027|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|501938680|1|0|2|502356100|1|0|2|500493871|2||500016307||2|1|500000294, 500016374|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|677715||4|3|45
500871683|BBBS of Greater Charlotte|Main Office|C|Completed|2007-10-01|2016-02-22|Followup|2014-10-01|2014-10-28|Complete|Done|4|2|1|1|4|3|2.5|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||2|3|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|Amachi|Child: Graduated|100.7||1|1|1|1|M|Black||19|Yes|Aunt|28208|One Parent: Female|Unknown|Y|No||Self|General Community|Amachi|Match Support|M|White||46|28209|Masters Degree|Single|Self-Employed, Entrepreneur|28209|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500871952|31|0|1|500933829|1|0|1|500199601|2||500003586||4|1|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|677733||4|3|45
501989028|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-22|2016-08-30|Followup|2014-10-22|2014-12-17|Complete|Late|3|2|2|3|3|4|2.83|4|1|4|1|4|4|3|-5.67|3|3|3|3|3|3|3|2|3|4|3|4|4|3.33|-9.91|4|4|4|4|4|3|4|3.67|8.99|4|4|3|3|3.5|5|4|4|4|4.25|-17.65|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|3|3|3|2|3|2.5|20|2|2|2|2|0|4|4|4|4|0|Yellow||Child/Family: Moved|46.3||2|2|1|1|M|Black||15|No|Mother|28273|One Parent: Female|Unknown||Yes|AARTF|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28273|Juris Doctorate (JD)|Single|Law: Lawyer||0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017777|502425720|31|0|1|503039778|31|0|1|500641725|2||-2||4|2||500005291|-2||-2|6855|8|||7496|10|635|1|1|677913|251884|4|3|45
500186133|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-14|2016-06-28|Followup|2014-10-14|2014-11-25|Complete|Done|2|2|2|2|2|2|2|||||||||4|4|4|3|4|3|3.67|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|140.5||1|1|1|1|M|White||18||Mother|28273|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||51|28262|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|500187724|1|0|1|500188930|1|0|1|500036930|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|678546||4|3|45
501372080|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-31|2016-04-22|Followup|2014-10-31|2014-12-12|Complete|Done|3|2|2|2|3|3|2.5|||||||||4|4|4|3|1|4|3.33|||||||||4|4|4|4||||||3|3|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Yellow||Child/Family: Moved|41.7||2|2|2|2|M|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community||Match Support|M|White||31|28269|Masters Degree|Single|Insurance|28262|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|501372359|31|0|1|502500246|1|0|1|500640327|2||-2||4|2|||-2||-2|0|3|||7496|10|||1|678548||4|3|45
502338225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-27|2016-05-26|Followup|2014-10-27|2014-12-11|Complete|Done|4|4|4|2|4|4|3.67|3|2|3|1|4|4|2.83|29.68|4|4|4|4|4|4|4|2|3|2|2|3|3|2.5|60|4|4|4|4|3|3|3|3|33.33|4|4|4|5|4.25|2|3|2|3|2.5|70|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|3|3|3|2|3|2.5|20|2|2|1|1|100|4|4||||Yellow|Project Big|Volunteer: Lost contact with child/agency|67||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||Yes||School|General Community|Project Big|Match Support|F|White||33|28227|Bachelors Degree|Single|Unknown||9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500008321|502338658|31|0|2|502312449|1|0|2|500483095|2||500004641||4|2|500004640|500004640|-2|500004640|-2|0|4|||7496|10|||1|678549|194054|4|3|45
502359051|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-28|2017-02-28|Followup|2014-10-28|2014-12-12|Complete|Done|4|4|4|4|4|4|4|||||||||2|3|3|3|2|3|2.67|||||||||3|4|4|3.67||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|76.1||1|1|1|1|F|Black||14|Yes|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||35|28213|Masters Degree|Married|Business: Clerical||3|6|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|502359489|31|0|2|502242295|31|0|2|500483954|2||500004772||4|3|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|10|||131|1|||1|678550||4|3|45
503328958|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-04|NaT|Baseline|2013-11-20|2013-11-26|Complete|Done|3|3|1|3|3|4|2.83|||||||||1|4|3|1|1|4|2.33|||||||||3|3|3|3||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|2|3||||||4|2|3|||||1|1||||4|4||||Green|||39.4||1|1|1|1|M|Black||15|No|Mother|28213|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|White||31|28203||Single|Law|28202|3|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503330792|31|0|1|503574852|1|0|1|500733114|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|679637|-1|4|3|44
503071479|BBBS of Greater Charlotte|Main Office|C|Active|2012-09-30|NaT|Followup|2014-09-30|2014-11-17|Declined|Late||||||||3|3|3|3|2|2|2.67|||||||||3|2|2|3|3|2|2.5||||||4|4|4|4|||||||4|3|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||3|3|3|3|||||||||||2|2||||4|4||Green|||53.5||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|M|White||28|28269|Some College|Single|Business: Clerical||0|3|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500020910|503069483|31|0|1|503051382|1|0|1|500629193|2||-2||2|1|||-2||-2|0|10|||7671|13|||1|680172|485271|4|1|45
502264006|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-22|2017-02-26|Followup|2014-09-22|2014-09-22|Complete|Done|3|3|4|3|3|3|3.17|2|1|3|1|2|3|2|58.5|2|2|3|2|2|4|2.5|1|3|2|2|1|3|2|25|4|4|4|4|4|4|4|4|0|4|5|3|3|3.75|4|2|3|4|3.25|15.38|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|2|3|3|4|3|3.33|-9.91|4|4|4|4|3|3.5|14.29|2|2|1|1|100|4|4||||Red||Child: Lost interest|77.2||1|1|1|1|F|Hispanic||16|No|Mother|28211|One Parent: Female|Unknown||Yes|Spanish Print|Media|General Community||Match Support|F|Hispanic||38|28202|Bachelors Degree|Single|Tech: Engineer|28202|12|0|Big Day|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020753|502264438|3|0|2|502274748|3|0|2|500470897|2||-2||4|3|||-2||-2|7063|1|||7456|8|||1|680173|178842|4|3|45
502353937|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-22|NaT|Followup|2014-11-22|2014-11-26|Complete|Done|3|4|4|2|3|4|3.33|||||||||2|4|3|2|2|3|2.67|||||||||4|3|4|3.67||||||2|4|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||2|4|3|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||75.8||1|1|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown|Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||31|29605|Bachelors Degree|Single|Business: Human Resources|29615|1|0|Local TV|Media|Big|General Community|Project Big AND Amachi|Match Support|277|60|598|500000170|500018851|502354375|31|0|2|501672025|1|0|2|500487322|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500004901|-2|0|4|||7438|1|||1|680419||4|3|45
502008563|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-21|2015-11-19|Followup|2014-11-21|2015-01-06|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Time constraint|23.9||2|2|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28210|Some College||Business||0|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|502008962|31|0|1|503400112|1|0|1|500730792|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|680515||4|1|45
500252077|BBBS of Greater Charlotte|Main Office|C|Completed|2008-11-24|2016-01-20|Followup|2014-11-24|2014-12-10|Complete|Done|3|4|2|1|3|2|2.5|||||||||2|1|4|2|2|3|2.33|||||||||4|3|2|3||||||4|3|2|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|85.8||3|3|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|Unknown||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Tech: Computer/Programmer||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|501750989|31|0|1|501365749|1|0|1|500317108|2||500003586||4|3|500000294|500000294|-2||-2|7295|11|||46|2|||1|680697||4|3|45
501014187|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-07|NaT|Followup|2014-11-07|2014-11-11|Complete|Done|3|4|4|4|3|4|3.67|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|3|2|||||2|2||||4|4||||Green|Amachi||100.2||2|2|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|White||48|28205|Bachelors Degree|Living w/ Significant Other|Human Services: Non-Profit|28205|3|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|500948399|31|0|2|501404007|1|0|2|500306699|2||500003586||2|1|500000294|500000294|-2||-2|0|10|||7671|13|||1|681377||4|3|45
500970495|BBBS of Greater Charlotte|Main Office|C|Completed|2008-09-10|2017-03-09|Followup|2014-09-10|2014-11-25|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Volunteer: Lost contact with child/agency|101.9||3|3|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$35,000 to $39,999||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black|Other African|44|28212||Single|Consultant||1|5|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|500970766|31|0|2|500965698|31|31|2|500285645|2||-2||4|2|||-2||-2|7294|13|||46|2|||1|681767||4|0|45
503617980|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-25|2016-01-06|Followup|2014-11-25|2014-12-11|Complete|Done|3|2|3|4|3|4|3.17|4|2|4|4|4|4|3.67|-13.62|3|2|3|3|3|3|2.83|2|4|4|3|4|3|3.33|-15.02|4|4|4|4|4|4|4|4|0|3|3|3|3|3|4|5|5|5|4.75|-36.84|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|4|4|3|3.67|-18.26|2|2|2|1|3|2|0|2|2|2|2|0|4|4|4|4|0|Green||Child/Family: Moved|25.4||1|1|1|1|F|Black||13|No|Mother|28217|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|White||25|28134|Some College|Single|Child/Day Care Worker||0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503619857|31|0|2|503573243|1|0|2|500730441|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|681979|675746|4|3|45
503701025|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-25|2016-08-18|Followup|2014-11-25|2014-12-11|Complete|Done|3|2|2|3|3|3|2.67|4|1|4|1|3|4|2.83|-5.65|3|2|3|4|4|3|3.17|1|1|1|1|1|4|1.5|111.33|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|4|4|5|5|4.5|-27.78|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|2|2|4|3|3.5|-42.86|2|2|2|2|0|4|4|4|4|0|Green||Volunteer: Time constraint|32.8||1|1|1|1|F|Black||12|Yes|Mother|28269|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|White||53|28227|Some College|Married|Customer Service|28105|30|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|501153063|31|0|2|503576358|1|0|2|500731543|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|681986|677325|4|3|45
502371558|BBBS of Greater Charlotte|Main Office|C|Active|2011-10-31|NaT|Followup|2014-10-31|2014-12-10|Complete|Done|3|3|3|2|3|4|3|3|2|3|3|3|3|2.83|6.01|3|4|3|2|3|3|3|3|4|4|3|2|4|3.33|-9.91|4|4|4|4|4|4|4|4|0|2|3|3|2|2.5|4|4|4|5|4.25|-41.18|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|3|4|3|3.33|4|4|3|3.67|-9.26|2|2|2|4|2|3|-33.33|2|2|1|1|100|4|4|4|4|0|Green|||64.5||1|1|2|2|M|Black||17|No|Mother|28206|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020752|502371997|31|0|1|502528355|1|0|1|500568298|2||-2||2|1||500000294, 500005291|-2||-2|0|10|||132|8|||1|682012|355033|4|3|45
502602958|BBBS of Greater Charlotte|Main Office|C|Completed|2011-09-11|2017-02-23|Followup|2014-09-11|2014-10-28|Declined|Late||||||||4|1|1|2|3|4|2.5|||||||||4|3|4|4|4|4|3.83||||||4|4|4|4|||||||5|3|5|5|4.5||||||||||4|4|4|4|4|4|3|3.86||||||3|4|4|3.67|||||2|3|2.5||||2|2||||4|4||Green|Project Big, 2010-2012 OJJDP JJI|Child/Family: Lost contact with volunteer/agency|65.4||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||52|28207|Masters Degree|Married|Business|28202|0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|501480402|31|0|1|502578040|1|0|1|500552390|2||500004641||4|1|500004640, 500005291|500004640, 500005291|-2||-2|0|4|||7464|9|||1|682445|333955|4|1|45
503021417|BBBS of Greater Charlotte|Main Office|C|Completed|2012-09-11|2015-10-16|Followup|2014-09-11|2014-10-28|Declined|Late||||||||3|3|4|2|3|4|3.17|||||||||3|4|3|2|3|3|3||||||4|4|4|4|||||||4|5|3|4|4||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|3|2.5||||1|1||||4|4||Yellow||Child/Family: Moved|37.1||1|1|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|White||32|28204|Bachelors Degree|Single|Business: Marketing|29730|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|501428579|31|0|2|503115600|1|0|2|500631553|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|682453|489252|4|1|45
500713817|BBBS of Greater Charlotte|Main Office|C|Active|2009-10-30|NaT|Followup|2014-10-30|2014-11-10|Complete|Done|3|3|4|3|3|4|3.33|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|||88.5||2|2|1|1|M|Black||16||Mother|28216|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28078|||Medical: Pharmacist|28210|10|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|500714084|31|0|1|501834795|1|0|1|500396466|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|682513||4|3|45
503569117|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-19|2015-03-12|Baseline|2013-11-27|2013-12-19|Complete|Done|3|2|4|3|3|4|3.17|||||||||2|3|4|3|3|4|3.17|||||||||4|3|4|3.67||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||1|1||||4|4||||Green||Child/Family: Moved|14.7||1|1|1|1|F|Black||15|No|Mother|2649|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||32|28203|Doctor of Medicine (MD)|Living w/ Significant Other|Medical|28112|1|2|other|College Partner|Big|General Community||Enrollment|277|60|598|500000170|500015820|503570990|31|0|2|503583743|1|0|2|500735247|2||-2||4|1|||-2||-2|0|10|||7670|5|||1|683133|-1|4|3|44
501000843|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-17|2015-09-24|Followup|2014-10-17|2015-01-01|Expired|Late||||||||4|3|4|2|4|4|3.5|||||||||2|4|3|2|3|3|2.83||||||4|4|4|4|||||||2|5|3|3|3.25||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|1|1.5||||1|1||||4|4||Red||Child/Family: Lost contact with volunteer/agency|35.2||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$25,000 to $29,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||26|28269|Bachelors Degree|Single|Business|28262|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|501001116|31|0|2|503106526|31|0|2|500632934|2||-2||4|3|||-2||-2|34|2|||7496|10|||1|683966|491461|4|0|45
503594290|BBBS of Greater Charlotte|Main Office|C|Active|2014-01-14|NaT|Baseline|2013-12-02|2014-01-14|Complete|Done|3|2|4|1|4|4|3|||||||||2|2|4|2|3|2|2.5|||||||||3|4|4|3.67||||||4|3|3|2|3|||||||4|4|4|4|4|3|3|3.71||||||||||3|4|4|3.67||||||3|4|3.5|||||1|1||||4|4||||Green|||38||1|1|1|1|M|Multi-Race (None of the above)||13|No|Mother|28134|Other Relative|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|M|Hispanic||26|28205|||Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503596167|7|0|1|503508074|3|0|1|500735488|2||-2||2|1|||-2||-2|0|5|||7464|9|||1|684069|-1|4|3|44
500829028|BBBS of Greater Charlotte|Main Office|C|Active|2010-11-30|NaT|Followup|2014-11-30|2014-12-11|Complete|Done|3|3|3|3|4|3|3.17|||||||||3|4|3|2|4|3|3.17|||||||||4|4|4|4||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||75.5||3|3|2|2|F|Black||17|No|Mother|28209|One Parent: Female|Less than $10,000|Y|No||Self|General Community||Match Support|F|White||39|28210|Masters Degree|Single|Education|28212|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500020910|502254499|31|0|2|501978180|1|0|2|500498594|2||-2||2|1|||-2|500000294, 500004640|-2|0|10|||7464|9|||1|684142||4|3|45
503017622|BBBS of Greater Charlotte|Main Office|C|Inactive|2012-09-19|NaT|Followup|2014-09-19|2014-09-15|Complete|Done|3|4|3|3|3|4|3.33|3|2|2|2|2||||3|3|3|2|3|4|3|3|4|4|3|3|4|3.5|-14.29|4|3|4|3.67|4|4|4|4|-8.25|3|3|3|3|3|4|3|3|3|3.25|-7.69|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|4|4|3.67|-9.26|3|3|3|3|3|3|0|2|2|2|2|0|4|4|4|4|0|Green|||53.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|$30,000 to $34,999|Y|No|BBBS National Site|Web Link|General Community||Match Support|F|White||33|28207|Bachelors Degree|Married|Business||0|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|503019155|31|0|2|503095382|1|0|2|500631726|2||-2||3|1|||-2||-2|34|2|||7464|9|||1|684147|489657|4|3|45
501129781|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-15|2015-01-15|Followup|2014-11-15|2014-12-11|Complete|Done|3|2|2|2|3|3|2.5|||||||||3|2|3|2|3|3|2.67|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||2|2|||||||||Green||Child: Family structure changed|50||1|2|4|6|F|Black||17||Mother|28217|Two Parent|Unknown||No||School|General Community||Match Support|F|Black||48|28273|Bachelors Degree|Married|Business: Mgt, Admin|28273|4|0|Recruitment Event|Neighbor/Friend|Big|General Community||Enrollment|277|60|598|500000170|500018987|501130055|31|0|2|500189245|31|0|2|500494855|2||-2||4|1|||-2||-2|0|4|||7459|10|||1|684158||4|3|45
502510347|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-31|2016-08-30|Followup|2014-10-31|2014-12-29|Declined|Late||||||||4|1|2|1|4|4|2.67|||||||||1|4|2|2|2|2|2.17||||||4|4|4|4|||||||3|4|2|4|3.25||||||||||4|4|4|4|4|4|2|3.71||||||3|2|1|2|||||4|2|3||||1|1||||4|4||Green|2010-2012 OJJDP JJI|Child: Graduated|58||1|1|1|1|F|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28262|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|502510796|31|0|2|502677833|31|0|2|500557844|2||-2||4|1|500005291|500005291|-2||-2|0|5|||7464|9|||1|684174|310349|4|1|45
501604446|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-19|NaT|Followup|2014-09-19|2014-12-02|Declined|Late|2|3|3|3|2|3|2.67|||||||||2|2|2|1|3|2|2|||||||||||||||||||||||||||||3|4|4|4|4|4|3|3.71||||||||||2|4|2|2.67||||||||||||||||||4|4||||Green|2010-2012 OJJDP JJI||65.9||2|2|1|1|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28213|Bachelors Degree|Married|Tech: Support, Writing|28273|11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500017732|501604760|31|0|1|502664359|31|0|1|500555050|2||-2||2|1|500005291|500005291|-2||-2|0|10|||7462|13|||1|685010||4|1|45
502234905|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-05|2015-08-25|Followup|2014-12-05|2014-12-08|Complete|Done|3|4|3|2|2|2|2.67|||||||||2|3|3|3|4|3|3|||||||||3|3|3|3||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Volunteer: Time constraint|44.6||3|3|1|1|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28083|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|M|White||36|28097|Masters Degree|Divorced|Finance|28026|7|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500012459|502777258|38|0|1|502799047|1|0|1|500583119|2||-2||4|1|500000294|500000294, 500014681, 500016374|-2||-2|0|10|||7671|13|||1|685026||4|3|45
503328958|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-04|NaT|Followup|2014-12-04|2014-12-08|Complete|Done|3|3|4|2|3|4|3.17|3|3|1|3|3|4|2.83|12.01|1|4|4|2|2|4|2.83|1|4|3|1|1|4|2.33|21.46|4|4|4|4|3|3|3|3|33.33|3|4|4|3|3.5|4|3|4|4|3.75|-6.67|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|4|3.67|3|4|2|3|22.33|3|3|3|4|2|3|0|2|2|1|1|100|4|4|4|4|0|Green|||39.4||1|1|1|1|M|Black||15|No|Mother|28213|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|White||31|28203||Single|Law|28202|3|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503330792|31|0|1|503574852|1|0|1|500733114|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|685287|679637|4|3|45
500868942|BBBS of Greater Charlotte|Main Office|C|Active|2007-09-20|NaT|Followup|2014-09-20|2014-12-05|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||113.8|Y|1|1|1|1|M|Black||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|M|White||54|28207||Married|Business: Sales||0|0|Recruitment Event|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|500869211|31|0|1|500947018|1|0|1|500195082|2||-2||2|1|||-2||-2|0|10|||7458|9|||1|685513||4|0|45
503441472|BBBS of Greater Charlotte|Main Office|C|Completed|2014-02-21|2016-05-03|Baseline|2013-12-05|2014-02-21|Complete|Done|2|4|4|3|4|3|3.33|||||||||3|3|2|4|2|3|2.83|||||||||4|4|3|3.67||||||3|2|5|4|3.5|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|26.3||1|1|1|1|F|Black||14|No|Mother|28212|One Parent: Female|$20,000 to $24,999|Y|No||School|General Community||Match Support|F|Black||28|28216|Masters Degree|Single|Consultant|28205|0|0|Recruitment Event|Self|Big|General Community||Enrollment|277|60|598|500000170|500021785|501290021|31|0|2|503551607|31|0|2|500738115|2||-2||4|1|||-2||-2|0|4|||7458|9|||1|685870|-1|4|3|44
503606415|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-06|2017-02-28|Baseline|2013-12-05|2014-01-06|Complete|Done|4|3|4|1|4|4|3.33|||||||||2|3|2|3|2|3|2.5|||||||||4|4|4|4||||||2|2|3|2|2.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|37.7||1|1|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|White||32|28270|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503608292|31|0|2|503665457|1|0|2|500736909|2||-2||4|1|||-2||-2|0|4|||7464|9|||1|685873|-1|4|3|44
503597088|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-06|2016-05-03|Followup|2014-12-06|2015-01-27|Declined|Late||||||||4|1|4|2|4|4|3.17|||||||||3|4|3|2|4|4|3.33||||||4|4|4|4|||||||4|3|3|3|3.25||||||||||4|4|4|4|3|4|3|3.71||||||3|4|4|3.67|||||1|2|1.5||||2|2||||4|4||Green||Volunteer: Moved|28.9||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Retail: Sales|28217|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503598965|31|0|2|503642924|1|0|2|500731612|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|686155|677446|4|1|45
503219503|BBBS of Greater Charlotte|Main Office|C|Completed|2014-02-05|2017-01-26|Baseline|2013-12-06|2014-02-05|Complete|Done|3|4|4|4|4|4|3.83|||||||||1|3|3|1|3|3|2.33|||||||||4|4|4|4||||||2|3|4|5|3.5|||||||4|4|4|4|3|4|4|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|35.7||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Multi-race (Hispanic & White)||33|28226|Some College|Single|Tech: Management|28277|1|7|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|503221284|31|0|1|503589945|35|0|1|500746532|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|686234|-1|4|3|44
502813527|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-09|NaT|Followup|2014-12-09|2015-01-15|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||39.2||1|2|1|2|F|Black||12|No|Mother|28031|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|White||62|28031|Masters Degree|Married|Real Estate: Realtor|28031|8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|502814804|31|0|2|502691411|1|0|2|500736806|2||-2||2|1|||-2||-2|0|4|||7496|10|||1|686999||4|3|45
503417576|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-09|2015-12-30|Followup|2014-12-09|2015-01-12|Complete|Done|4|1|2|1|3|3|2.33|3|1|2|1|3|3|2.17|7.37|1|1|1|1|1|3|1.33||2|2|2|2|1|||4|4|4|4|3|3|4|3.33|20.12|4|3|5|4|4|2|3|3|2|2.5|60|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|4|3.67|4|4|4|4|-8.25|3|3|3|2|3|2.5|20|2|2|1|1|100|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|24.7||1|1|1|1|F|White||17|No|Father|28269|Two Parent|$100,000 to $124,999|Y|No||Relative|General Community||Match Support|F|White||29|28205|Some College|Single|Business: Mgt, Admin|29707|3|10|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|503419440|1|0|2|503594017|1|0|2|500730510|2||-2||4|3|||-2|500000294|-2|0|3|||7464|9|||1|687058|675823|4|3|45
502629201|BBBS of Greater Charlotte|Main Office|C|Active|2012-03-22|NaT|Followup|2014-03-22|2014-04-03|Complete|Done|3|4|4|2|1|3|2.83|||||||||4|3|4|2|2|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|||59.8||2|2|1|1|M|White||12|No|Mother|28277|One Parent: Female|$60,000 to $74,999||No||Self|General Community||Match Support|M|White||32|28210|Bachelors Degree|Single|Business: Mgt, Admin|28226|1|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502629856|1|0|1|502893231|1|0|1|500603253|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|687264||4|3|45
503688885|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-18|NaT|Baseline|2013-12-11|2013-12-18|Complete|Done|4|4|4|1|4|4|3.5|||||||||1|4|4|4|4|4|3.5|||||||||4|4|4|4||||||1|5|5|5|4|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||1|2|1.5|||||1|1||||4|4||||Green|||38.9||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||35|28204|Bachelors Degree|Single|Retail: Mgt|28273|1|10|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|503690850|31|0|2|503606993|1|0|2|500738203|2||-2||2|1|||-2||-2|0|10|||46|2|||1|687980|-1|4|3|44
500185907|BBBS of Greater Charlotte|Main Office|C|Completed|2006-10-29|2015-02-18|Followup|2014-10-29|2014-12-14|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|99.7||2|3|1|1|F|Black||19|Yes|Mother|28262|One Parent: Female|Unknown||No||Self|General Community|Amachi|Match Support|F|Black||48|28212||Single|Medical: Healthcare Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|500187470|31|0|2|500697782|31|0|2|500134557|2||500003586||4|3|500000294|500000294|-2|500000294|-2|0|10|||2238|7|||1|688154||4|1|45
500826592|BBBS of Greater Charlotte|Main Office|C|Completed|2009-10-08|2016-10-18|Followup|2014-10-08|2014-12-23|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|84.3||3|3|1|1|F|Black||20|No|Mother|28226|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community||Match Support|F|White||33|28277|Bachelors Degree|Living w/ Significant Other|Unknown|28209|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|500826861|31|0|2|501314246|1|0|2|500382768|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|688708||4|0|45
502674024|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-07|2016-05-17|Followup|2014-12-07|2014-12-10|Complete|Done|4|3|4|4|4|4|3.83|4|4|4|3|4|4|3.83|0|3|4|4|3|1|4|3.17|2|4|4|4|4|3|3.5|-9.43|4|4|4|4|4|4|4|4|0|3|5|3|3|3.5|4|4|4|3|3.75|-6.67|4|4|4|3|4|4|4|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|3|4|3|3.33|20.12|3|1|2|3|3|3|-33.33|2|2|2|2|0|4|4|4|4|0|Green||Child: Lost interest|53.3||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Sales||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018851|502674852|31|0|2|502660051|1|0|2|500581910|2||-2||4|1||500005291|-2||-2|0|10|||7496|10|||1|688817|374331|4|3|45
502183420|BBBS of Greater Charlotte|Main Office|C|Completed|2010-09-28|2015-01-15|Followup|2014-09-28|2014-12-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|Amachi|Volunteer: Time constraint|51.6||2|2|1|1|M|Multi-race (Black & White)||14|Yes|GrandMother|28215|Grandparents|Unknown||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||58|28226|Masters Degree|Married|Tech: Sales, Mktg|28202|6|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500015820|502183840|36|0|1|502264770|1|0|1|500473793|2||500003586||4|2|500000294|500000294|-2||-2|7016|11|||7464|9|||1|688981||4|0|45
500186742|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-08|2016-06-30|Followup|2014-12-08|2014-12-10|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|3|4|4|3|3|3.33|||||||||4|4|4|4||||||2|5|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Green|Amachi|Child: Graduated|66.7||4|4|1|1|M|Black||19|Yes|Mother|28227|One Parent: Female|Unknown|Y|No||School|General Community|Amachi|Match Support|M|Black||52|28227|Masters Degree|Married|Education: Teacher|28227|2|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500013781|500188056|31|0|1|502397541|31|0|1|500501282|2||500003586||4|1|500000294|500000294|-2|500000294, 500004640|-2|0|4|||12183|14|635|1|1|689080||4|3|45
502920861|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-29|2016-04-22|Followup|2014-10-29|2014-12-12|Complete|Done|4|2|3|3|2|3|2.83|4|2|3|3|4|3|3.17|-10.73|1|3|3|2|2|3|2.33|4|2|3|4|4|2|3.17|-26.5|4|4|4|4|4|4|4|4|0|3|3|3|3|3|5|3|5|5|4.5|-33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3|3.71|7.82|4|4|4|4|4|4|3|3.67|8.99|4|4|4|3|3|3|33.33|2|2|1|1|100|4|4|4|4|0|Yellow||Child/Family: Lost contact with volunteer/agency|41.8||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||34|28203|Juris Doctorate (JD)|Single|Law: Lawyer||2|11|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502922278|31|0|1|503097126|1|0|1|500639233|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|689344|499329|4|3|45
500185812|BBBS of Greater Charlotte|Main Office|C|Completed|2012-10-29|2016-05-26|Followup|2014-10-29|2014-12-12|Complete|Done|2|2|3|2|3|3|2.5|||||||||2|3|3|4|4|3|3.17|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green||Child: Graduated|42.9||2|3|2|3|F|Black||18|Yes|Mother|28210|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community|Amachi|Match Support|F|White||41|28214|Bachelors Degree|Single|Human Services: Non-Profit||3|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|500187400|31|0|2|500188912|1|0|2|500648551|2||-2||4|1||500000294|-2||-2|0|10|||7464|9|||1|689345||4|3|45
501771263|BBBS of Greater Charlotte|Main Office|C|Completed|2009-09-29|2017-02-28|Followup|2014-09-29|2014-12-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|89||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|Black||31|28262|Bachelors Degree|Single|Medical: Admin|28216|0|8|Recruitment Event|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|501741899|31|0|2|501622704|31|0|2|500379993|2||-2||4|1|||-2||-2|0|10|||7443|2|||1|689408||4|0|45
503424337|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-19|2016-05-26|Followup|2014-07-19|2014-09-09|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|34.2||1|1|1|1|F|Black||12||Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Match Support|F|Black||30|28173|Masters Degree|Single|Education|28262|0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503426202|31|0|2|503446943|31|0|2|500703604|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|689507||4|1|45
503565123|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-23|2014-03-03|Baseline|2013-12-16|2014-01-23|Complete|Done|4|2|3|4|3|4|3.33|||||||||4|2|2|2|1|3|2.33|||||||||1|4|1|2||||||5|1|3|4|3.25|||||||4|4|4|4|2|1|3|3.14||||||||||4|3|1|2.67||||||2|1|1.5|||||2|2||||4|4||||Green||Volunteer: Moved|1.3||1|1|1|1|M|Black||12|No|Mother|28213|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|White||30|28262|Masters Degree|Single|Tech: Engineer|28078|2|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503566998|31|0|1|503673127|1|0|1|500739078|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|689782|-1|4|3|44
503496815|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-13|2015-06-19|Baseline|2013-12-17|2014-01-10|Complete|Done|3|1|2|1|3|4|2.33|||||||||2|3|4|4|4|4|3.5|||||||||3|4|3|3.33||||||5|4|3|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red||Volunteer: Time constraint|17.1||1|1|1|1|M|Black||13|No|Mother|28034|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||26|28217|Bachelors Degree|Single|Tech: Engineer|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500015820|503773736|31|0|1|503673962|31|0|1|500739342|2||-2||4|3|||-2||-2|0|10|||7496|10|||1|690298|-1|4|3|44
502580335|BBBS of Greater Charlotte|Main Office|C|Active|2011-11-30|NaT|Followup|2014-11-30|2015-02-14|Expired|Late||||||||3|2|1|1|1|3|1.83|||||||||2|4|3|1|4|3|2.83||||||4|4|3|3.67|||||||5|2|4|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||3|2|2.5||||2|2||||4|4||Green|||63.5||1|1|1|1|F|Black||16||GrandMother|28269|Grandparents|Unknown||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28269|Masters Degree|Single|Finance: Banking|28255|15|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|502580838|31|0|2|502677590|31|0|2|500571804|2||-2||2|1||500005291|-2||-2|0|10|||7464|9|||1|690507|355336|4|0|45
502868969|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-18|NaT|Followup|2014-12-18|2014-12-18|Complete|Done|3|2|3|3||3||2|4|4|4|3|4|3.5||3|4|3|3|4|1|3|2|4|4|1|3|3|2.83|6.01|4|3|3|3.33|4|4|4|4|-16.75|3|2|3|3|2.75|5|5|4|4|4.5|-38.89|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|3|4|3|3.33|20.12|3|3|3|2|4|3|0|2|2|2|2|0|4|4|4|4|0|Green|||38.9||1|1|1|1|F|Black||17|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||26|11237||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020753|502870370|31|0|2|503574667|1|0|2|500736904|2||-2||2|1|||-2|500000294|-2|0|10|||46|2|||1|690770|611488|4|3|45
503688885|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-18|NaT|Followup|2014-12-18|2015-03-04|Expired|Late||||||||4|4|4|1|4|4|3.5|||||||||1|4|4|4|4|4|3.5||||||4|4|4|4|||||||1|5|5|5|4||||||||||4|4|4|4|4|4|2|3.71||||||4|4|4|4|||||1|2|1.5||||1|1||||4|4||Green|||38.9||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||35|28204|Bachelors Degree|Single|Retail: Mgt|28273|1|10|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017732|503690850|31|0|2|503606993|1|0|2|500738203|2||-2||2|1|||-2||-2|0|10|||46|2|||1|690922|687980|4|0|45
503689205|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-08|2015-10-20|Baseline|2013-12-18|2014-01-08|Complete|Done|4|3|4|1|4|4|3.33|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|21.4||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|Black||46|28227|Masters Degree|Married|Finance|28202|8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503691170|31|0|2|503689218|31|0|2|500739856|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|691058|-1|4|3|44
502776341|BBBS of Greater Charlotte|Main Office|C|Active|2012-12-14|NaT|Followup|2014-12-14|2014-12-15|Complete|Done|3|4|3|3|3|4|3.33|||||||||3|4|4|2|4|4|3.5|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|||51||1|2|1|2|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||Yes||School|General Community||Match Support|F|White||31|28202|Bachelors Degree|Single|Retail: Mgt|28273|6|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|502777520|31|0|2|502631040|1|0|2|500652764|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|691114||4|3|45
503569117|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-19|2015-03-12|Followup|2014-12-19|2015-01-15|Complete|Done|3|1|3|3|3|4|2.83|3|2|4|3|3|4|3.17|-10.73|3|3|3|1|3|4|2.83|2|3|4|3|3|4|3.17|-10.73|4|4|4|4|4|3|4|3.67|8.99|3|5|4|5|4.25|4|4|5|5|4.5|-5.56|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|3|4|3.67|4|4|4|4|-8.25|4|4|4|2|4|3|33.33|2|2|1|1|100|4|4|4|4|0|Green||Child/Family: Moved|14.7||1|1|1|1|F|Black||15|No|Mother|2649|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||32|28203|Doctor of Medicine (MD)|Living w/ Significant Other|Medical|28112|1|2|other|College Partner|Big|General Community||Enrollment|277|60|598|500000170|500015820|503570990|31|0|2|503583743|1|0|2|500735247|2||-2||4|1|||-2||-2|0|10|||7670|5|||1|691364|683133|4|3|45
502702145|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-21|2016-05-24|Followup|2014-12-21|2014-12-22|Complete|Done|3|4|4|3|4|4|3.67|3|3|4|3|4|4|3.5|4.86|4|4|4|4|4|4|4|3|4|4|4|4|4|3.83|4.44|4|4|4|4|3|3|3|3|33.33|5|5|5|5|5|5|4|2|4|3.75|33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|3|3|3|2|3|2.67|12.36|2|4|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Red||Child: Graduated|53.1||1|1|2|2|F|Black||17|No|Mother|28083|One Parent: Female|$60,000 to $74,999||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500020753|502702991|31|0|2|502204211|31|0|2|500582836|2||-2||4|3|||-2||-2|6854|8|||7464|9|||1|691395|375724|4|3|45
501273088|BBBS of Greater Charlotte|Main Office|C|Completed|2012-11-28|2017-02-28|Followup|2014-11-28|2014-12-29|Complete|Done|3|1|1|1|1|2|1.5|||||||||3|3|3|2|3|4|3|||||||||4|4|4|4||||||3|2|3|2|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|51||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Unknown||Yes||Relative|General Community||Match Support|F|Black||48|28213|Bachelors Degree|Single|Finance: Accountant||8|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|501273365|31|0|2|503079327|31|0|2|500659156|2||-2||4|1|||-2||-2|0|3|||7464|9|||1|691903||4|3|45
503662377|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-31|2017-02-28|Baseline|2013-12-20|2014-01-31|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|2|2|3|2.5|||||||||3|3|3|3||||||4|3|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|36.9||1|1|1|1|F|Black||13|No|Mother|28216|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503664337|31|0|2|503573326|1|0|2|500743531|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|691921|-1|4|3|44
503689574|BBBS of Greater Charlotte|Main Office|C|Completed|2014-03-20|2016-03-09|Baseline|2013-12-20|2014-03-19|Complete|Done|3|4|4|1|1|1|2.33|||||||||1|2|2|3|2|2|2|||||||||4|4|4|4||||||5|3|2|2|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green||Volunteer: Moved|23.7||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Unknown|Y|Yes||Therapist/Counselor|General Community||Enrollment|F|White||33|28210|PHD|Single|Business: Human Resources|28273|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|503691539|31|0|2|503577882|1|0|2|500751079|2||-2||4|1|||-2||-2|0|5|||7464|9|||1|691927|-1|4|3|44
503490571|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-20|2015-05-14|Followup|2014-12-20|2015-01-14|Complete|Done|3|2|3|3|3|3|2.83|3|4|4|3|3|3|3.33|-15.02|2|3|3|3|2|3|2.67|4|4|4|3|4|4|3.83|-30.29|3|3|3|3|4|4|4|4|-25|3|4|4|4|3.75|4|5|5|5|4.75|-21.05|4|4|4|3|3|4|4|3.71|4|3|4|4|4|4|4|3.86|-3.89|3|3|3|3|4|4|4|4|-25|3|3|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Red|VOL - Mentoring Hispanic Youth|Child/Family: Lost contact with volunteer/agency|16.8||1|1|1|1|F|Hispanic|Mexican|16|No|Mother|28208|Two Parent|Unknown|Y|Yes|Spanish Radio|Media|General Community||Match Support|F|White||35|28214|Bachelors Degree|Single|Transport: Flight Attendant|85034|0|3|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|503492439|3|10|2|503645850|1|0|2|500738556|2||-2||4|3|500011312||-2|500000294|-2|7068|1|||7464|9|||1|692105|659479|4|3|45
502180724|BBBS of Greater Charlotte|Main Office|C|Active|2010-12-30|NaT|Followup|2014-12-30|2014-12-29|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|3|2|4|3.17|||||||||4|4|4|4||||||5|1|5|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Amachi, Project Big, Project Big AND Amachi||74.5|Y|2|2|2|2|M|Black||15|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|502181148|31|0|1|502391505|31|0|2|500505039|2||500004772||2|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7438|1|||1|692504||4|3|45
502604900|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-15|2015-05-14|Followup|2014-11-15|2015-01-05|Declined|Late||||||||3|1|1|1|1|1|1.33|||||||||1|1|2|1|1|3|1.5||||||4|4|4|4|||||||4|4|3|3|3.5||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||4|2|3||||1|1||||4|4||Green||Volunteer: Lost contact with child/agency|41.9||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||30|28211|Bachelors Degree|Single|Finance: Accountant|28204|0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502605417|1|0|1|502582742|1|0|1|500577855|2||-2||4|1|||-2|500000294|-2|6854|8|||7464|9|||1|692515|356462|4|1|45
500337327|BBBS of Greater Charlotte|Main Office|C|Active|2006-12-14|NaT|Followup|2014-12-14|2014-12-29|Complete|Done|3|1|4|4|4|1|2.83|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||3|1|3|5|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Green|||123||2|3|4|5|M|Black||16||GrandMother|28208|Grandparents|Unknown||No||School|General Site||Match Support|M|Black||49|28217|Associate Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site||Match Support|277|60|598|500000170|500017732|500251937|31|0|1|500189300|31|0|1|500148262|2||-2||2|1|||-1||-1|0|4|||7464|9|||1|692529||4|3|45
502747706|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-17|2015-10-09|Followup|2014-11-17|2015-01-05|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|46.7||1|1|1|1|F|Multi-Race (None of the above)||13|No|Mother|28229|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Enrollment|F|Black||34|28226|Bachelors Degree|Single|Business: Clerical|28208|0|6|Self|Self|Big|General Community|Project Big|Enrollment|277|60|598|500000170|500017777|502748616|7|0|2|502618438|31|0|2|500566066|2||-2||4|3|||-2|500004640|-2|0|10|||7464|9|||1|692554||4|1|45
502184849|BBBS of Greater Charlotte|Main Office|C|Active|2012-12-18|NaT|Followup|2014-12-18|2014-12-17|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||5|5|4|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|||50.9||2|2|1|1|M|Multi-race (Hispanic & White)||13|No|Mother|28211|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||28|28210|Bachelors Degree|Single|Business: Marketing|28224|1|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|502185278|35|0|1|503145815|1|0|1|500658541|2||-2||2|1|||-2||-2|0|10|||7496|10|||1|692555||4|3|45
502290468|BBBS of Greater Charlotte|Main Office|C|Completed|2012-02-10|2015-09-16|Followup|2014-02-10|2014-03-27|Complete|Done|2|2|2|2|3|3|2.33|||||||||2|3|2|2|2|3|2.33|||||||||3|3|3|3||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child/Family: Moved|43.2||1|1|1|1|M|Black||12|No|Mother|28227|One Parent: Female|Unknown||Yes||School|General Community||Match Support|M|Multi-race (Hispanic & White)||33|28204|PHD||Medical: Doctor, Provider||0|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502290900|31|0|1|502873884|35|0|1|500596681|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|693207||4|3|45
502507408|BBBS of Greater Charlotte|Main Office|C|Completed|2011-10-13|2016-08-22|Followup|2014-10-13|2014-12-28|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow|2010-2012 OJJDP JJI|Volunteer: Lost contact with child/agency|58.3||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Less than $10,000||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||71|28277|Bachelors Degree|Married|Retired||0|0||Relative|Big|General Community||Match Support|277|60|598|500000170|500017732|502507857|31|0|1|502673562|31|0|1|500559678|2||-2||4|2|500005291||-2||-2|34|2|||0|11|||1|693257||4|0|45
502222548|BBBS of Greater Charlotte|Main Office|C|Active|2010-08-24|NaT|Followup|2014-08-24|2014-09-04|Complete|Done|3|1|4|3|3|2|2.67|||||||||2|3|3|3|4|4|3.17|||||||||3|1|1|1.67||||||4|2|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green|||78.7||1|1|1|1|M|Black||12|No|Mother|28216|One Parent: Female|Unknown||No||School|General Community||Match Support|M|White||40|28211|Bachelors Degree|Married|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020753|502222979|31|0|1|502214317|1|0|1|500465659|2||-2||2|1|||-2|500000294|-2|0|4|||7496|10|||1|693429||4|3|45
502308197|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-03|2016-05-09|Followup|2014-12-03|2014-12-18|Complete|Done|3|3|4|2|4|3|3.17|||||||||3|2|3|3|4|4|3.17|||||||||1|1|1|1||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|65.2||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||Yes||Self|General Community|Amachi|Enrollment|F|White||35|28210|Bachelors Degree|Living w/ Significant Other|Business: Sales|18034|2|7|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big AND Amachi|Match Support|277|60|598|500000170|500021785|502308629|31|0|2|502325667|1|0|2|500493122|2||500003586||4|1||500000294|-2|500000294, 500004901|-2|0|10|||7496|10|||1|693537||4|3|45
502367953|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-18|2016-01-26|Followup|2014-08-18|2014-09-29|Complete|Done|4|3|3|4|4|4|3.67|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi|Child/Family: Lost contact with volunteer/agency|53.3||1|1|1|1|M|Black||12|Yes|Mother|28208|One Parent: Female|Unknown|Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||43|28212|Masters Degree|Married|Retail: Mgt||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|502368391|31|0|1|502658210|31|0|1|500548740|2||500003586||4|2|500000294|500000294|-2||-2|6854|8|||46|2|||1|693735||4|3|45
501353940|BBBS of Greater Charlotte|Main Office|C|Active|2011-11-30|NaT|Followup|2014-11-30|2014-11-25|Complete|Done|4|1|4|2|4|4|3.17|||||||||3|4|3|4|3|3|3.33|||||||||4|4|4|4||||||5|3|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Amachi||63.5||3|3|1|1|M|Black||16|No|Relative: Other|28205|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||33|28226|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|10|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500020752|501354219|31|0|1|502710990|1|0|1|500574615|2||500003586||2|1|500000294|500000294, 500005291|-2||-2|34|2|||17161|11|||1|694239||4|3|45
501123191|BBBS of Greater Charlotte|Main Office|C|Completed|2010-10-20|2015-12-21|Followup|2014-10-20|2015-01-04|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|62||2|2|1|1|F|Black||15|No|Mother|28227|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||48|28210|Some College|Single|Human Services||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500017732|500915629|31|0|2|502153920|1|0|2|500478644|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|694542||4|0|45
502728289|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-04|2017-03-09|Followup|2014-11-04|2015-01-19|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|64.1||1|1|1|1|F|Hispanic||13|No|Mother|28278|One Parent: Female|Less than $10,000|Y|Yes||Relative|General Community||Match Support|F|White||32|28211||Married|Finance||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|502729186|3|0|2|502339145|1|0|2|500565493|2||-2||4|1|||-2|500000294|-2|0|3|||7496|10|||1|694545||4|0|45
503556065|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-10|2015-10-09|Baseline|2014-01-06|2014-01-10|Complete|Done|3|3|4|2|4|4|3.33|||||||||4|4|3|2|3|4|3.33|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|20.9||1|1|3|3|M|Black||16|No|Mother|28269|One Parent: Female|$50,000 to $59,999||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017777|503557940|31|0|1|501284751|31|0|1|500741332|2||-2||4|2|||-2|500007920, 500011315, 500011316|-2|34|2|||132|8|||1|694970|-1|4|3|44
503671116|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-10|2017-02-23|Baseline|2014-01-06|2014-01-10|Complete|Done|4|2|4|3|4|4|3.5|||||||||2|3|3|3|2|4|2.83|||||||||4|4|4|4||||||2|5|2|3|3|||||||2|3|2|1|3|2|1|2||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2||||4|4||||Green||Volunteer: Moved|37.5||1|1|1|1|M|White||17|No|GrandMother|28278|One Parent: Female|$20,000 to $24,999||No||Self|General Community||Match Support|M|White||37|29708|Bachelors Degree|Single|Real Estate: Realtor|28273|1|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|503673077|1|0|1|503672609|1|0|1|500741347|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|694988|-1|4|3|44
500496598|BBBS of Greater Charlotte|Main Office|C|Active|2008-10-23|NaT|Followup|2014-10-23|2014-10-24|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|4|4|4|3.67|||||||||4|4|4|4||||||3|4|3|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|Amachi, Cabarrus County||100.7||2|2|1|1|M|White||15|Yes|Mother|28083|One Parent: Female|Unknown||No|BBBS National Site|Web Link|General Community|Amachi, Cabarrus County|Match Support|M|White||35|28083|Masters Degree|Single|Business: Mgt, Admin|28027|2|3|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|500496849|1|0|1|501383928|1|0|1|500299090|2||500003586||2|2|500000294, 500016374|500000294, 500016374|-2|500016374|-2|34|2|||7464|9|||1|695087||4|3|45
503662199|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-17|2016-07-29|Baseline|2014-01-08|2014-01-17|Complete|Done|4|4|4|4|4|3|3.83|||||||||2|3|4|3|2|4|3|||||||||4|4|4|4||||||2|4|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||3|3|3|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|30.4||1|1|1|1|M|Black||17|No|Mother|28270|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|M|White||32|28226|Bachelors Degree|Married|Consultant|28202|4|4|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|503664159|31|0|1|503639494|1|0|1|500741727|2||-2||4|2|||-2|500000294|-2|0|10|||7464|9|||1|695544|-1|4|3|44
502859187|BBBS of Greater Charlotte|Main Office|C|Active|2012-11-24|NaT|Followup|2014-11-24|2014-12-11|Complete|Done|2|3|2|2|3|2|2.33|2|2|4|2|4|4|3|-22.33|3|2|3|2|3|3|2.67|2|3|3|3|3|4|3|-11|4|4|3|3.67|4|4|4|4|-8.25|3|3|2|4|3|4|5|3|3|3.75|-20|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|4|4|4|4|-16.75|3|2|2.5|4|4|4|-37.5|2|2|2|2|0|4|4|4|4|0|Green|VOL - PreMatch||51.7||2|2|1|1|F|Black||15|No|GrandMother|28205|Grandparents|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|White||31|28209|Associate Degree|Married|Retail: Mgt|28134|4|3|UNCC|College Partner|Big|General Community||Match Support|277|60|598|500000170|500008321|500187987|31|0|2|503090888|1|0|2|500658723|2||-2||2|1|500007920||-2||-2|0|10|||9221|5|||1|695701|400467|4|3|45
501252806|BBBS of Greater Charlotte|Main Office|C|Active|2008-11-25|NaT|Followup|2014-11-25|2015-01-09|Complete|Done|3|4|4|2|4|4|3.5|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||99.6||1|1|1|1|M|Black||13|No|Mother|28078|One Parent: Female|Unknown||No||Relative|General Community||Match Support|M|Black||45|28262|Bachelors Degree|Married|Business: Mgt, Admin||0|6|AA Task Force|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|501253082|31|0|1|501320197|31|0|1|500310204|2||-2||2|1|||-2||-2|0|3|||6247|12|||1|695702||4|3|45
502255225|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-08|2016-08-26|Followup|2014-11-08|2014-12-29|Declined|Late||||||||2|2|2|4|1|4|2.5|||||||||2|3|3|2|2|3|2.5||||||4|3|3|3.33|||||||5|3|5|3|4||||||||||4|3|4|4|4|4|4|3.86||||||4|4|4|4|||||1|1|1||||1|1|||||||Red||Volunteer: Moved|69.6||1|1|1|1|M|Hispanic||15||Mother|28212|One Parent: Female|Unknown||No|Spanish Radio|Media|General Community||Match Support|M|White||33|28226|Bachelors Degree|Single|Education: Teacher||3|0|Spanish Print|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|502255655|3|0|1|502312682|1|0|1|500487118|2||-2||4|3|||-2||-2|7068|1|||11662|1|||1|696203|199091|4|1|45
500186260|BBBS of Greater Charlotte|Main Office|C|Completed|2004-10-29|2015-12-17|Followup|2014-10-29|2015-01-13|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|133.6||3|3|1|1|M|Black||19|No|Mother|28025|One Parent: Female|Unknown||No||Self|General Site||Match Support|M|Black||42|28025|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002335|500187857|31|0|1|500189139|31|0|1|500037139|2||-2||4|2|||-1||-2|0|10|||7464|9|||1|696669||4|0|45
503547661|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-23|2015-08-06|Baseline|2014-01-14|2014-01-23|Complete|Done|4|1|3|2|4|4|3|||||||||4|4|3|2|2|4|3.17|||||||||4|4|4|4||||||4|5|3|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green||Child/Family: Moved|18.4||1|1|1|1|M|Black||12|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28277|Bachelors Degree|Divorced|Business|28273|4|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503549536|31|0|1|503731665|1|0|1|500742652|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|697106|-1|4|3|44
503587930|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-27|2015-02-05|Baseline|2014-01-14|2014-01-27|Complete|Done|3|3|4|2|3|3|3|||||||||4|||4|3|4||||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|12.3||1|1|3|3|M|Black||16|No|Mother|28215|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|White||26|28203|Bachelors Degree|Single|Finance: Banking|28213|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503589807|31|0|1|500942257|1|0|1|500742670|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|697130|-1|4|3|44
503163476|BBBS of Greater Charlotte|Main Office|C|Active|2012-11-30|NaT|Followup|2014-11-30|2015-01-14|Complete|Done|2|2|2|2|3|3|2.33|3|1|1|1|1|3|1.67|39.52|2|3|3|3|3|3|2.83|2|3|4|2|3|3|2.83|0|3|3|3|3|3|4|4|3.67|-18.26|3|3|3|3|3|4|5|5|5|4.75|-36.84|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|3|3|4|4|4|4|-25|3|3|3|1|2|1.5|100|2|2|2|2|0|4|4|4|4|0|Green|||51.5||1|1|1|1|M|Black||13|No|Mother|28269|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|Black||32|28217|Masters Degree|Single|Consultant||0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503165154|31|0|1|503119713|31|0|1|500663695|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|697459|530536|4|3|45
503486227|BBBS of Greater Charlotte|Main Office|C|Active|2013-10-31|NaT|Followup|2014-10-31|2014-11-25|Complete|Done|2|4|4|3|3|2|3|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|2|3.33||||||3|3|3|||||2|2||||4|4||||Green|||40.5||1|1|1|1|M|Black||12|No|Mother|28270|One Parent: Female|$30,000 to $34,999||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||32|28210|Bachelors Degree|Single|Tech: Research/Design|28273|0|9|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|503186577|31|0|1|503555261|31|0|1|500725969|2||-2||2|1|||-2|500000294|-2|34|2|||46|2|||1|697483||4|3|45
503664796|BBBS of Greater Charlotte|Main Office|C|Completed|2014-01-31|2014-05-23|Baseline|2014-01-15|2014-01-31|Complete|Done|4|2|3|1|3|4|2.83|||||||||3|3|3|3|1|3|2.67|||||||||3|4|4|3.67||||||4|3|3|4|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|2|2.67||||||2|2|2|||||1|1||||4|4||||Green||Volunteer: Feels incompatible with child/family|3.7||1|1|1|1|M|Black||17|No|Mother|28227|One Parent: Female|$45,000 to $49,999|Y|Yes||Self|General Community||Match Support|M|White||51|28210|Bachelors Degree|Domestic Partner|Arts, Entertainment, Sports|28210|0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500002334|503666756|31|0|1|503674336|1|0|1|500744967|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|697540|-1|4|3|44
502247579|BBBS of Greater Charlotte|Main Office|C|Completed|2011-12-02|2016-05-10|Followup|2014-12-02|2014-12-29|Complete|Done|2|4|4|4|4|4|3.67|4|3|3|2|3|4|3.17|15.77|4|4|4|4|4|4|4|2|3|2|2|2|3|2.33|71.67|4|4|4|4|4|4|4|4|0|5|3|3|4|3.75|3|3|3|3|3|25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|4|4|-3.5|4|4|3|3.67|4|4|4|4|-8.25|3|2|2.5|3|3|3|-16.67|2|2|2|2|0|4|4||||Green|Amachi, Project Big, Project Big AND Amachi|Child/Family: Lost contact with volunteer/agency|53.3||2|2|1|1|F|Black||15|Yes|Mother|28217|One Parent: Female|Unknown||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||47|28226|Bachelors Degree|Single|Education: Teacher||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500017732|502248010|31|0|2|502681447|31|0|2|500575685|2||500003586||4|1|500000294, 500004640, 500004901|500000294, 500004640, 500004901|-2||-2|0|10|||2238|7|||1|698069|194970|4|3|45
502278991|BBBS of Greater Charlotte|Main Office|C|Active|2010-12-03|NaT|Followup|2014-12-03|2015-01-16|Complete|Done|4|3|3|2|4|4|3.33|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|||75.4||1|1|1|1|F|Black||12|No|Mother|28213|One Parent: Female|Unknown||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||40|28269|Bachelors Degree|Married|Tech: Management|28255|1|9|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502279417|31|0|2|502263116|31|0|2|500494784|2||-2||2|1|||-2|500000294|-2|6854|8|||6247|12|||1|698313||4|3|45
502589869|BBBS of Greater Charlotte|Main Office|C|Completed|2011-11-30|2015-10-29|Followup|2014-11-30|2015-01-13|Declined|Done||||||||4|2|2|3|1|1|2.17|||||||||2|4|4|4|4|4|3.67||||||4|4|4|4|||||||4|5|4|5|4.5||||||||||4|3|4|4|4|4|3|3.71||||||4|3|4|3.67|||||2|3|2.5||||2|2||||4|4||Green|Project Big|Child/Family: Lost contact with volunteer/agency|46.9||2|2|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28205|Bachelors Degree|Married|Business|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017777|502590381|31|0|2|502701252|1|0|2|500582617|2||500004641||4|1|500004640|500004640, 500005291|-2|500000294|-2|0|4|459|3|7496|10|||1|699253|290937|4|1|45
501069450|BBBS of Greater Charlotte|Main Office|C|Completed|2007-11-07|2017-02-28|Followup|2014-11-07|2014-11-13|Complete|Done|3|4|4|3|4|4|3.67|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|Amachi|Volunteer: Lost contact with child/agency|111.7||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||66|28075||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|501048131|31|0|1|500887364|31|0|1|500212043|2||-2||4|1|500000294|500000294|-2||-2|5635|9|||7464|9|||1|699534||4|3|45
503395663|BBBS of Greater Charlotte|Main Office|C|Completed|2014-02-21|2015-10-08|Baseline|2014-01-22|2014-02-21|Complete|Done|4|3|4|4|4|4|3.83|||||||||2|4|4|4|2|3|3.17|||||||||4|3|4|3.67||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||2|2||||4|4||||Green||Volunteer: Moved|19.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|$10,000 to $14,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28204|Masters Degree|Single|Finance: Accountant|28202|4|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503397520|31|0|1|503735537|1|0|1|500744097|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|699578|-1|4|3|44
500733695|BBBS of Greater Charlotte|Main Office|C|Completed|2006-12-26|2015-03-03|Followup|2014-12-26|2015-02-08|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red|Amachi|Child/Family: Lost contact with volunteer/agency|98.2||1|1|1|1|F|Black||19|Yes|GrandMother|28217|Grandparents|Less than $10,000|Y|No|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||34|28210|Bachelors Degree|Married|Finance: Accountant|28202|0|2|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|277|60|598|500000170|500013781|500733962|31|0|2|500307108|1|0|2|500150172|2||500003586||4|3|500000294|500000294|-2||-2|7294|13|||2238|7|||1|702572||4|1|45
501863951|BBBS of Greater Charlotte|Main Office|C|Completed|2009-12-18|2015-05-29|Followup|2014-12-18|2015-01-30|Complete|Done|3|2|4|2|4|4|3.17|||||||||2|3|3|4|4|4|3.33|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Red||Child: Lost interest|65.3||1|1|2|2|F|Black||14|No|Mother|28216|One Parent: Female|Unknown|Y|Yes||Self|General Community||Match Support|F|Black||37|28078|Bachelors Degree|Single|Business: Human Resources|28226|0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|501864324|31|0|2|501601161|31|0|2|500421259|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|703694||4|3|45
503634718|BBBS of Greater Charlotte|Main Office|C|Active|2014-02-27|NaT|Baseline|2014-02-04|2014-02-22|Complete|Done|2|1|1|1|1|2|1.33|||||||||4|4|2|1|2|3|2.67|||||||||3|2|2|2.33||||||3|2|4|2|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|2|2.5|||||1|1||||4|4||||Green|Cabarrus County||36.6||1|1|1|1|F|White||14|No|Father|28081|One Parent: Male|$15,000 to $19,999||Yes||Self|General Community|Cabarrus County|Match Support|F|White||28|28209|Bachelors Degree|Single|Finance|28217|3|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500013781|503636659|1|0|2|503595858|1|0|2|500746721|2||-2||2|1|500016374|500016374|-2|500016374|-2|0|10|||7458|9|||1|704398|-1|4|3|44
502308593|BBBS of Greater Charlotte|Main Office|C|Completed|2010-11-23|2015-05-28|Followup|2014-11-23|2015-01-20|Declined|Late||||||||4|2|3|1|3|4|2.83|||||||||3|3|4|4|3|3|3.33||||||3|2|3|2.67|||||||3|4|5|2|3.5||||||||||4|4|4|4|4|4|4|4||||||3|4|3|3.33|||||2|3|2.5||||1|1|||||||Red||Child/Family: Moved|54.1||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||40|28278|Bachelors Degree|Married|Tech: Computer/Programmer||3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|277|60|598|500000170|500008321|502309025|31|0|1|502262702|31|0|1|500492994|2||-2||4|3|||-2||-2|0|10|||12183|14|1209|1|1|705608|206463|4|1|45
503268271|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-27|2015-08-19|Followup|2014-12-27|2015-02-10|Complete|Done|3|3|3|2|4|4|3.17|3|4|4|1|4|4|3.33|-4.8|2|4|4|4|3|3|3.33|2|4|3|4|4|4|3.5|-4.86|4|3|3|3.33|4|4|4|4|-16.75|3|3|4|2|3|5|4|5|4|4.5|-33.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|4|4|4|4|-25|3|3|3|4|2|3|0|1|1|2|2|-50|4|4|4|4|0|Red||Volunteer: Lost contact with child/agency|31.7||1|1|1|1|F|Black||13|No|Mother|28226|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||40|28273|Some College|Married|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500008321|503270085|31|0|2|502993922|1|0|2|500669147|2||-2||4|3|||-2||-2|6854|8|||7496|10|3|3|1|706051|533978|4|3|45
502760967|BBBS of Greater Charlotte|Main Office|C|Active|2011-12-08|NaT|Followup|2014-12-08|2014-12-16|Complete|Done|3|3|2|3|3|4|3|1|2|4|1|3|3|2.33|28.76|3|4|4|4|4|4|3.83|4|4|4|4|3|4|3.83|0|4|4|4|4|4|2|2|2.67|49.81|3|3|3|3|3|5|5|5|5|5|-40|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|2|2|4|3|3.5|-42.86|2|2|2|2|0|4|4|4|4|0|Green|||63.2||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|$25,000 to $29,999|Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||29|28120|Bachelors Degree|Single|Govt: Clerical||0|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500021785|502761879|31|0|2|502666332|31|0|2|500579826|2||-2||2|1||500005291|-2||-2|2203|12|||7464|9|||1|707359|351583|4|3|45
500261295|BBBS of Greater Charlotte|Main Office|C|Completed|2005-12-21|2017-03-09|Followup|2014-12-21|2015-03-07|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child: Graduated|134.6||1|1|1|1|M|White||20||Mother|28104|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|White||60|28270|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500017732|500261310|1|0|1|500188435|1|0|1|500073081|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|707365||4|0|45
502335675|BBBS of Greater Charlotte|Main Office|C|Completed|2010-12-30|2016-10-31|Followup|2014-12-30|2015-02-13|Complete|Done|4|4|4|3|3|4|3.67|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red|Amachi, Project Big, Project Big AND Amachi|Child: Lost interest|70||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||Yes||School|General Community|Project Big AND Amachi|Match Support|M|White||27|28262||Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|277|60|598|500000170|500008321|502336110|31|0|1|502305990|1|0|1|500495220|2||500004772||4|3|500000294, 500004640, 500004901|500004901|-2|500000294, 500004640|-2|0|4|||7496|10|||1|708158||4|3|45
503638969|BBBS of Greater Charlotte|Main Office|C|Active|2013-12-20|NaT|Followup|2014-12-20|2014-12-29|Complete|Done|3|3|1|1|3|4|2.5|||||||||2|3|3|1|4|3|2.67|||||||||4|4|4|4||||||2|3||||||||||4|4|4|4|4|3|3|3.71||||||||||4|4|3|3.67||||||2|3|2.5|||||2|2||||4|4||||Green|||38.8||1|1|1|1|F|Black||12|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||23|28227||Single|Student: College|28202|2|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020910|503640929|31|0|2|503503174|31|0|2|500736646|2||-2||2|1|||-2||-2|0|10|||46|2|||1|708294||4|3|45
502431040|BBBS of Greater Charlotte|Main Office|C|Completed|2011-08-31|2016-08-26|Followup|2014-08-31|2014-10-14|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Moved|59.9||1|1|1|1|M|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||35|28207|Masters Degree|Married|Law: Lawyer|28202|8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|277|60|598|500000170|500020910|502431483|31|0|1|502609637|1|0|1|500550314|2||-2||4|1|||-2|500004640|-2|0|10|||7496|10|||1|710183||4|1|45
501347056|BBBS of Greater Charlotte|Main Office|C|Completed|2008-12-12|2015-10-12|Followup|2014-12-12|2015-01-27|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Graduated|82||1|1|1|1|M|Black||20|No|Mother|28217|One Parent: Female|Unknown||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28226|Bachelors Degree|Married|Tech: Engineer|28202|2|8|Recruitment Event|Workplace Partner|Big|General Community||Match Support|277|60|598|500000170|500017777|501347335|31|0|1|501217000|1|0|1|500322327|2||-2||4|2|||-2||-2|34|2|||7446|3|||1|712379||4|1|45
502983808|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-15|2016-02-10|Followup|2014-12-15|2015-01-30|Declined|Late||||||||1|1|2|1|1|3|1.5|||||||||1|4|4|1|1|3|2.33||||||4|4|4|4|||||||1|5|3|5|3.5||||||||||4|4|4|4|4|4|4|4||||||3|1|1|1.67|||||3|4|3.5||||1|1||||4|4||Yellow|Amachi|Volunteer: Time constraint|37.8||1|1|1|1|M|Black||15|Yes|Mother|28205|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Amachi|Match Support|M|White||27|28203|Bachelors Degree|Single|Business||0|2|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502985262|31|0|1|503140432|1|0|1|500668771|2||-2||4|2|500000294|500000294|-2|500000294|-2|0|4|||7464|9|||1|714410|538016|4|1|45
503433257|BBBS of Greater Charlotte|Main Office|C|Completed|2013-05-07|2014-09-04|Followup|2014-05-07|2014-06-26|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Child/Family: Lost contact with volunteer/agency|15.9||1|1|1|1|F|Black||12|No|Father|28213|One Parent: Male|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||55|28269|Associate Degree|Single|Business||28|0|Self|Self|Big|General Community||RTBM|277|60|598|500000170|500017777|503435122|31|0|2|503384599|31|0|2|500695071|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|714498||4|1|45
503703048|BBBS of Greater Charlotte|Main Office|C|Active|2014-03-12|NaT|Baseline|2014-03-04|2014-03-12|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|4|4|2|4|4|3.33|||||||||4|4|3|3.67||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|3|3|||||1|1||||4|4||||Green|||36.1||1|1|1|1|M|White||12|No|Mother|28226|One Parent: Female|$200,000 or more||No||Self|General Community||Match Support|M|White||59|28104|Bachelors Degree|Married|Finance||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|503705013|1|0|1|503354824|1|0|1|500753007|2||500009594||2|1|||-2||-2|0|10|1562|2|7671|13|1561|2|1|715206|-1|4|3|44
503401214|BBBS of Greater Charlotte|Main Office|C|Active|2014-03-26|NaT|Baseline|2014-03-04|2014-03-26|Complete|Done|4|4|2|4|4|3|3.5|||||||||2|4|4|4|2|4|3.33|||||||||4|4|3|3.67||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Yellow|||35.7||1|1|1|1|M|Black||12|No|Mother|28105|One Parent: Female|$50,000 to $59,999||No||Self|General Community||Match Support|M|White||31|28226|Bachelors Degree|Single|Finance: Accountant|28217|4|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020910|503403071|31|0|1|503758808|1|0|1|500752693|2||-2||2|2|||-2||-2|0|10|||7496|10|||1|715251|-1|4|3|44
503565637|BBBS of Greater Charlotte|Main Office|C|Active|2014-03-15|NaT|Baseline|2014-03-05|2014-03-12|Complete|Done|4|1|1|1|4|4|2.5|||||||||1|4|4|1|1|4|2.5|||||||||3|4|4|3.67||||||5|1|1|4|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||36||1|1|1|1|M|Black||12|Yes|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||49|28204|Bachelors Degree|Married|Finance: Accountant|28255|8|0|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|277|60|598|500000170|500020910|503567522|31|0|1|503604089|1|0|1|500752839|2||-2||2|1||500000294|-2|500000294, 500014681|-2|34|2|||7464|9|||1|715551|-1|4|3|44
503532014|BBBS of Greater Charlotte|Main Office|C|Completed|2014-03-21|2015-07-08|Baseline|2014-03-10|2014-03-21|Complete|Done|4|2|4|1|4|2|2.83|||||||||4|4|3|1|4|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|2|4|3.33||||||4|4|4|||||1|1||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|15.6||2|2|2|2|M|White||12|No|Mother|28025|One Parent: Female|$15,000 to $19,999||Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||58|28075|Masters Degree|Married|Business|32824|0|6|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500012459|503533889|1|0|1|503694720|1|0|1|500753716|2||-2||4|2||500000294, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7464|9|||1|717073|-1|4|3|44
503756716|BBBS of Greater Charlotte|Main Office|C|Completed|2014-03-31|2016-01-14|Baseline|2014-03-12|2014-03-31|Complete|Done|1|4|4|3|4|4|3.33|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green||Child: Lost interest|21.5||1|1|1|1|F|Black||14|No|Mother|28215|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||29|28270||Single|Unemployed||0|0|Self|Self|Big|General Community|Amachi|Enrollment|277|60|598|500000170|500020990|503758688|31|0|2|503596238|31|0|2|500754325|2||-2||4|1|||-2|500000294|-2|0|10|||7464|9|||1|718009|-1|4|3|44
503124706|BBBS of Greater Charlotte|Main Office|C|Completed|2014-03-31|2016-01-26|Baseline|2014-03-18|2014-03-31|Complete|Done|3|4|4|4|4|4|3.83|||||||||4|2|4|4|4|4|3.67|||||||||4|3|3|3.33||||||5|5|5|5|5|||||||3|4|3|3|3|3|3|3.14||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Green||Volunteer: Moved|21.9||1|1|1|1|M|Black||17|No|Mother|28226|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|Multi-race (Black & White)||29|28215|Some College|Married|Student: College|28223|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020752|503126373|31|0|1|503609606|36|0|1|500755317|2||-2||4|1|||-2||-2|0|10|||46|2|||1|719710|-1|4|3|44
502527969|BBBS of Greater Charlotte|Main Office|C|Completed|2012-12-01|2015-08-18|Followup|2014-12-01|2015-01-20|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Red||Child/Family: Lost contact with volunteer/agency|32.5||1|1|1|1|M|Black||11|No|Mother|28278|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|White||34|29708|High School Graduate|Single|Business: Mgt, Admin|29730|11|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502528422|31|0|1|503169378|1|0|1|500662254|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|720006||4|1|45
503479095|BBBS of Greater Charlotte|Main Office|C|Completed|2014-07-17|2016-03-29|Baseline|2014-03-21|2014-07-17|Complete|Done|4|1|2|1|4|4|2.67|||||||||2|3|4|2|3|4|3|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|2|2||||||||||4|4||||Green||Volunteer: Moved|20.4||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Enrollment|M|White||28|28270|Bachelors Degree|Married|Real Estate: Realtor|28203|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500021785|503480961|31|0|1|503915425|1|0|1|500768983|2||-2||4|1|||-2||-2|0|10|||46|2|||1|720937|-1|4|3|44
503758675|BBBS of Greater Charlotte|Main Office|C|Active|2014-03-27|NaT|Baseline|2014-03-24|2014-03-27|Complete|Done|3|4|4|2|1|3|2.83|||||||||2|4|4|1|2|4|2.83|||||||||4|3|3|3.33||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|3|3.5|||||1|1||||4|4||||Green|||35.6||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|M|Black||30|28202|Bachelors Degree|Single|Consultant|28281|2|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020910|503760648|31|0|1|503792275|31|0|1|500756323|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|721599|-1|4|3|44
503830048|BBBS of Greater Charlotte|Main Office|C|Completed|2014-04-08|2014-09-04|Baseline|2014-03-27|2014-04-08|Complete|Done|4|4|4|4|3|3|3.67|||||||||1|2|1|1|3|2|1.67|||||||||4|3|4|3.67||||||1|4|3|4|3|||||||4|3|4|4|3|4|3|3.57||||||||||2|2|1|1.67||||||1|2|1.5|||||2|2||||4|4||||Red||Volunteer: Feels incompatible with child/family|4.9||1|1|1|1|F|Hispanic||16|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||47|28205|Associate Degree|Single|Medical: Nurse||1|0|BBBS National Site|Web Link|Big|General Community||Enrollment|277|60|598|500000170|500017777|503832027|3|0|2|503559585|1|0|2|500757050|2||-2||4|3|||-2||-2|34|2|||46|2|||1|722998|-1|4|3|44
503429736|BBBS of Greater Charlotte|Main Office|C|Active|2014-04-29|NaT|Baseline|2014-03-28|2014-04-29|Complete|Done|3|1|3|4|4|3|3|||||||||1|3|2|4|2|3|2.5|||||||||3|2|2|2.33||||||5|3|4|5|4.25|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Green|||34.6||1|1|1|1|M|Black||14|No|Mother|28216|One Parent: Female|$60,000 to $74,999||No|AARTF|Neighbor/Friend|General Community||Match Support|M|White||27|28217|Masters Degree|Single|Finance|28202|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020753|503431601|31|0|1|503850437|1|0|1|500760086|2||-2||2|1|||-2||-2|6855|8|||17159|12|||1|723550|-1|4|3|44
503565188|BBBS of Greater Charlotte|Main Office|C|Completed|2014-04-22|2015-05-28|Baseline|2014-04-04|2014-04-22|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|4|4|1|4|4|3.17|||||||||3|2|3|2.67||||||4|5|3|4|4|||||||4|4|4|4|4|3|3|3.71||||||||||4|3|4|3.67||||||1|2|1.5|||||1|1||||4|4||||Yellow||Volunteer: Lost contact with child/agency|13.2||2|2|1|1|M|Black||12|No|Mother|28212|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Black||48|28269|Masters Degree|Married|Finance: Banking|28262|9|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|503567063|31|0|1|503814392|31|0|1|500758306|2||-2||4|2|||-2||-2|0|10|||46|2|||1|725936|-1|4|3|44
503524036|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-19|2017-02-28|Baseline|2014-04-06|2014-09-19|Complete|Done|2|4|4|2|1|1|2.33|||||||||3|1|2|2|2|3|2.17|||||||||3|4|3|3.33||||||1|2|4|4|2.75|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|PERL 2014-2016|Child/Family: Lost contact with volunteer/agency|29.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||39|28262|Bachelors Degree|Single|Finance|28262|3|2|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503525911|31|0|1|503913408|31|0|1|500774440|2||-2||4|1|500014681|500014681|-2|500014681|-2|0|10|||17159|12|||1|726336|-1|4|3|44
503710095|BBBS of Greater Charlotte|Main Office|C|Active|2014-06-19|NaT|Baseline|2014-04-08|2014-06-19|Complete|Done|4|4|3|2|3|4|3.33|||||||||1|2|3|3|1|3|2.17|||||||||3|4|3|3.33||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green|||32.9||1|1|1|1|M|Black||13|No|Mother|28202|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Finance: Accountant|28226|0|0|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500020910|503712061|31|0|1|503872736|1|0|1|500766579|2||-2||2|1|||-2||-2|0|10|||17101|1|||1|726855|-1|4|3|44
503722616|BBBS of Greater Charlotte|Main Office|C|Completed|2014-04-24|2015-10-19|Baseline|2014-04-08|2014-04-24|Complete|Done|3|3|2|3|1|3|2.5|||||||||3|3|2|2|3|3|2.67|||||||||4|3|2|3||||||3|3|2|3|2.75|||||||4|4|4|3|3|3|3|3.43||||||||||4|1|1|2||||||1|1|1|||||2|2||||4|4||||Green||Volunteer: Moved|17.8||2|2|1|1|F|Multi-race (Black & White)||15|No|Mother|28134|One Parent: Female|Unknown||Yes||Self|General Community||Match Support|F|White||55|28217|Some College|Married|Retail: Mgt|28217|14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503724588|36|0|2|503707316|1|0|2|500759403|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|726896|-1|4|3|44
503632799|BBBS of Greater Charlotte|Main Office|C|Active|2014-05-31|NaT|Baseline|2014-04-08|2014-05-31|Complete|Done|4|4|4|3|4|4|3.83|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||33.5||1|1|1|1|F|Black||13|No|Mother|28269|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||59|28209|Bachelors Degree|Divorced|Medical|28209|1|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503634738|31|0|2|503567146|1|0|2|500763613|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|726899|-1|4|3|44
503745830|BBBS of Greater Charlotte|Main Office|C|Completed|2014-04-23|2014-09-15|Baseline|2014-04-10|2014-04-23|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|4|3|4|3.67|||||||||4|2|2|2.67||||||4|2|4|2|3|||||||3|3|4|3|4|3|3|3.29||||||||||3|3|3|3||||||2|2|2|||||1|1||||4|4||||Yellow||Volunteer: Moved|4.8||1|1|1|1|M|Black||17|No|Mother|28206|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|M|Black||52|28212|Associate Degree|Divorced|Business: Mgt, Admin|60131|1|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503747802|31|0|1|503760503|31|0|1|500759184|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|727688|-1|4|3|44
503707241|BBBS of Greater Charlotte|Main Office|C|Completed|2014-04-30|2015-03-26|Baseline|2014-04-11|2014-04-30|Complete|Done|3|1|2|2|4|4|2.67|||||||||1|4|1|2|4|4|2.67|||||||||4|4|4|4||||||5|4|2|1|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Time constraint|10.8||1|1|1|1|F|Black||15|Yes|Mother|28214|One Parent: Female|$35,000 to $39,999|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Some Other Race||34|28216|Masters Degree|Living w/ Significant Other|Finance: Banking|28216|0|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018850|503709207|31|0|2|503767700|41|0|2|500759405|2||-2||4|1||500000294|-2||-2|34|2|||7464|9|||1|728131|-1|4|3|44
502146600|BBBS of Greater Charlotte|Main Office|C|Active|2014-04-30|NaT|Baseline|2014-04-14|2014-04-30|Complete|Done|3|3|4|3|3|3|3.17|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||3|1|1|1|1.5|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||1|3|2|||||2|2||||4|4||||Green|||34.5||1|1|2|2|F|Black||15|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||45|28227|Bachelors Degree|Married|Customer Service|28262|18|0|Big For A Day|Special Event|Big|General Community|Amachi|Match Support|277|60|598|500000170|500013781|502932575|31|0|2|503483337|31|0|2|500760757|2||-2||2|1|||-2|500000294|-2|6854|8|||16422|8|||1|728732|-1|4|3|44
503143377|BBBS of Greater Charlotte|Main Office|C|Active|2012-11-16|NaT|Followup|2014-11-16|2014-12-31|Complete|Done|2|2|3|2|2|3|2.33|||||||||2||2|3|3|3||||||||||3|2|2|2.33||||||2|2|3|3|2.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||3|3|3|||||2|2||||4|4||||Green|||51.9||1|1|1|1|F|Black||11|No|Mother|28210|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||28|28226|Bachelors Degree|Single|Education: Teacher|28173|2|6|TV|Media|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|503145049|31|0|2|503109316|1|0|2|500649731|2||-2||2|1|||-2|500000294|-2|0|10|||130|1|||1|732007||4|3|45
503770826|BBBS of Greater Charlotte|Main Office|C|Completed|2014-04-29|2015-04-30|Baseline|2014-04-25|2014-04-29|Complete|Done|3|2|3|2|2|3|2.5|||||||||4|2|3|4|4|4|3.5|||||||||4|4|4|4||||||2|4|5|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|12||1|1|1|1|M|White||15|No|Mother|28211|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||63|28105|Bachelors Degree|Married|Self-Employed, Entrepreneur|28105|7|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503772799|1|0|1|503820142|1|0|1|500761166|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|732698|-1|4|3|44
503706992|BBBS of Greater Charlotte|Main Office|C|Active|2014-04-30|NaT|Baseline|2014-04-28|2014-04-30|Complete|Done|3|2|2|2|3|4|2.67|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|4|3.5|||||1|1||||4|4||||Green|VOL - Mentoring Hispanic Youth||34.5||1|1|1|1|F|Hispanic|Mexican|13|No|Mother|28205|One Parent: Female|Unknown|Y|Yes|BBBS National Site|Web Link|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||44|28213|Bachelors Degree|Married|Medical|28216|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503708958|3|10|2|503709061|1|0|2|500761338|2||-2||2|1|500011312|500011312|-2||-2|34|2|||7464|9|||1|733329|-1|4|3|44
503584428|BBBS of Greater Charlotte|Main Office|C|Active|2014-05-14|NaT|Baseline|2014-04-30|2014-05-14|Complete|Done|1|4|4|3|3|4|3.17|||||||||4|2|4|3|2|4|3.17|||||||||4|4|4|4||||||4|3|4|2|3.25|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||2|1|1.5|||||1|1||||4|4||||Green|||34.1||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|Black||27|28216|Some College|Single|Retail: Sales||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503586305|31|0|1|503839843|31|0|1|500761714|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|734527|-1|4|3|44
503833956|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-12|2016-01-27|Baseline|2014-04-30|2014-05-12|Complete|Done|3|3|4|4|4|4|3.67|||||||||2|3|2|2|1|2|2|||||||||4|4|4|4||||||3|4|2|2|2.75|||||||4|4|4|4|2|3|2|3.29||||||||||4|3|3|3.33||||||3|2|2.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|20.5||1|1|1|1|F|Black||17|No|Mother|28208|Two Parent|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||38|28262|Masters Degree|Single|Finance|28262|0|6|Agency Sponsored|Special Event|Big|General Community|Amachi|Match Support|277|60|598|500000170|500018851|503835911|31|0|2|503635291|31|0|2|500761770|2||-2||4|1|||-2|500000294|-2|34|2|||16426|8|||1|734750|-1|4|3|44
503636487|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-27|NaT|Baseline|2014-05-02|2014-10-27|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|4|3|1|4|3.17|||||||||4|4|4|4||||||3|4|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||1|1||||4|4||||Green|PERL 2014-2016||28.6||1|1|1|1|M|Black||12|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28205|Bachelors Degree|Single|Finance: Accountant|28202|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503665377|31|0|1|503899296|1|0|1|500778337|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||17159|12|||1|735741|-1|4|3|44
502934728|BBBS of Greater Charlotte|Main Office|C|Active|2013-08-14|NaT|Followup|2014-08-14|2014-09-23|Complete|Done|3|2|3|2|3|3|2.67|||||||||2|4|3|3|3|3|3|||||||||3|4|4|3.67||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||43||1|1|1|1|M|Black||11|No|Mother|28215|One Parent: Female|$35,000 to $39,999||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||41|28211|Bachelors Degree|Single|Finance: Banking|28209|5|0|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|502936151|31|0|1|503516330|31|0|1|500705674|2||-2||2|1|||-2|500000294|-2|6854|8|||7464|9|||1|735825||4|3|45
503663975|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-22|2015-05-14|Baseline|2014-05-06|2014-05-22|Complete|Done|4|1|3|1|4|4|2.83|||||||||1|4|4|4|4|4|3.5|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|1|1|||||2|2||||4|4||||Red||Child/Family: Feels incompatible with volunteer|11.7||2|2|1|1|M|Black||13|Yes|Mother|28204|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community|Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Insurance|28277|5|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017777|503665933|31|0|1|503854225|31|0|1|500762272|2||-2||4|3||500000294|-2||-2|0|10|||17159|12|||1|736588|-1|4|3|44
503770823|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-15|2017-01-24|Baseline|2014-05-06|2014-05-15|Complete|Done|4|2|4|1|4|4|3.17|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||3|5|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green||Child/Family: Lost contact with volunteer/agency|32.4||1|1|1|1|M|White||13|No|Mother|28211|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||27|28270|Bachelors Degree|Single|Education: Teacher Asst/Aid|28202|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500021785|503772799|1|0|1|503850589|1|0|1|500762293|2||-2||4|1|||-2||-2|34|2|||46|2|||1|736644|-1|4|3|44
503381531|BBBS of Greater Charlotte|Main Office|C|Active|2014-06-05|NaT|Baseline|2014-05-08|2014-06-05|Complete|Done|4|4|4|3|4|4|3.83|||||||||3|4|4|2|2|4|3.17|||||||||4|4|4|4||||||4|3|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|||33.3||1|1|2|2|M|Black||14|No|Mother|28206|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||66|28269||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503383388|31|0|1|500540549|31|0|1|500762593|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|737860|-1|4|3|44
503717073|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-16|2016-10-14|Baseline|2014-05-09|2014-05-16|Complete|Done|4|3|2|1|4|4|3|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||3|1|1|5|2.5|||||||4|3|4|3|4|1|1|2.86||||||||||3|4|4|3.67||||||2|2|2|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|29||1|1|1|2|M|Black||14|Yes|Mother|28216|One Parent: Female|Unknown|Y|Yes||School|General Community||Match Support|M|Black||54|28277|Bachelors Degree|Single|Consultant|28202|7|6|Man Up Campaign|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Pending Match|277|60|598|500000170|500020910|503719040|31|0|1|503853194|31|0|1|500762798|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17101|1|||1|738691|-1|4|3|44
503813952|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-29|2015-05-14|Baseline|2014-05-09|2014-05-29|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||4|4|3|3|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|4|3|||||2|2||||4|4||||Green||Volunteer: Time constraint|11.5||1|1|1|1|F|Black||14|No|Mother|28262|One Parent: Female|$20,000 to $24,999|Y|No|BBBS National Site|Web Link|General Community||Enrollment|F|White||28|28202|Masters Degree|Single|Finance: Banking|28205|0|1|Other|Service Organization|Big|General Community||Match Support|277|60|598|500000170|500017732|503969639|31|0|2|503829786|1|0|2|500763221|2||-2||4|1|||-2||-2|34|2|||7452|6|||1|738695|-1|4|3|44
502299232|BBBS of Greater Charlotte|Main Office|C|Completed|2013-07-30|2015-08-17|Followup|2014-07-30|2014-10-14|Expired|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Yellow||Child: Family structure changed|24.6||1|1|1|1|M|Black||11|Yes|GrandMother|28273|Foster Home|$25,000 to $29,999|Y|Yes||Self|General Community|Amachi|Enrollment|M|White||32|28209|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|5|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500015820|501806520|31|0|1|503510609|1|0|1|500703319|2||-2||4|2||500000294|-2|500000294|-2|0|10|||7464|9|||1|738897||4|0|45
502653228|BBBS of Greater Charlotte|Main Office|C|Active|2011-09-11|NaT|Followup|2014-09-11|2014-10-22|Complete|Done|3|2|2|2|3|3|2.5|||||||||2|3|3|4|3|3|3|||||||||3|3|3|3||||||3|3|4|2|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|3|2.5|||||2|2||||4|4||||Green|||66.1||1|1|2|2|F|Black||11|No|Mother|28205|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|F|White||32|28134|Bachelors Degree|Single|Finance: Banking|28288|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502653964|31|0|2|502192090|1|0|2|500552244|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|738968||4|3|45
503774057|BBBS of Greater Charlotte|Main Office|C|Active|2014-05-23|NaT|Baseline|2014-05-12|2014-05-21|Complete|Done|2|2|4|1|1|3|2.17|||||||||3|1|2|2|2|2|2|||||||||3|4|4|3.67||||||2|3|1|1|1.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|||33.8||1|1|1|1|F|Multi-race (Black & Hispanic)||13|No|Mother|28215|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|White||61|28211|Bachelors Degree|Divorced|Tech: Management|28202|2|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503776034|38|0|2|503665969|1|0|2|500762915|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|739281|-1|4|3|44
503728057|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-22|2015-12-21|Baseline|2014-05-14|2014-05-22|Complete|Done|2|3|4|3|2|2|2.67|||||||||3|4|3|3|2|3|3|||||||||4|4|4|4||||||3|3|2|4|3|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|3|3.67||||||2|1|1.5|||||1|1||||4|4||||Yellow|Amachi|Volunteer: Feels incompatible with child/family|19||1|1|2|2|M|Black||15|Yes|Mother|28227|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|M|Black||30|28213|Masters Degree|Single|Education|28217|0|7|Recruitment Event|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|503730029|31|0|1|503788318|31|0|1|500763247|2||-2||4|2|500000294||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7458|9|||1|740487|-1|4|3|44
503755565|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-29|2015-08-06|Baseline|2014-05-21|2014-05-29|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|4|4|4|2|4|3.67|||||||||4|3|3|3.33||||||4|4|4|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow||Volunteer: Time constraint|14.3||1|1|1|1|M|Black||13|No|Mother|28227|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Enrollment|M|White||55|28031|Bachelors Degree|Separated|Business: Sales|53964|3|3|Local Print|Media|Big|General Community||Match Support|277|60|598|500000170|500015820|503757537|31|0|1|503814505|1|0|1|500763994|2||-2||4|2|||-2||-2|0|10|||7439|1|||1|745222|-1|4|3|44
503782875|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-30|2014-11-06|Baseline|2014-05-21|2014-05-30|Complete|Done|2|2|2|2|2|3|2.17|||||||||2|3|3|3|3|3|2.83|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||3|3||||Green||Agency: Challenges with program/partnership|5.3||1|1|1|1|F|Black||12|No|Mother|28227|Two Parent|$40,000 to $44,999||No|BBBS National Site|Web Link|General Community||Match Support|F|White||22|28206|Some College|Single|Child/Day Care Worker||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|503784852|31|0|2|503732680|1|0|2|500763995|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|745226|-1|4|3|44
503767186|BBBS of Greater Charlotte|Main Office|C|Active|2014-06-23|NaT|Baseline|2014-05-21|2014-06-23|Complete|Done|4|4|1|1|1|3|2.33|||||||||1|1|4|1|1|4|2|||||||||4|4|4|4||||||4|3|5|4|4|||||||4|4|4|4|4|4|2|3.71||||||||||3|4|4|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|||32.8||1|1|1|1|F|Black||16|No|Mother|28227|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Black||30|28205|Bachelors Degree|Single|Business|28262|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500020910|503769162|31|0|2|503788125|31|0|2|500766047|2||-2||2|1|||-2||-2|0|10|||46|2|||1|745252|-1|4|3|44
503816186|BBBS of Greater Charlotte|Main Office|C|Completed|2014-05-29|2014-10-20|Baseline|2014-05-21|2014-05-29|Complete|Done|3|4|2|2|3|4|3|||||||||2|3|3|4|3|4|3.17|||||||||3|3|3|3||||||3|4|3|3|3.25|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|3|3.33||||||1|4|2.5|||||2|2||||4|4||||Yellow||Volunteer: Feels incompatible with child/family|4.7||2|2|1|1|F|Black||14|No|Mother|28206|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||30|28226|Bachelors Degree|Single|Business: Human Resources|28203|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|501097065|31|0|2|501675299|31|0|2|500764043|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|745502|-1|4|3|44
502324604|BBBS of Greater Charlotte|Main Office|C|Completed|2013-10-30|2014-11-06|Followup|2014-10-30|2014-10-30|Complete|Done|4|4|2|1|3|4|3|||||||||1|4|4|1|3|4|2.83|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||3|3|4|3.33||||||3|2|2.5|||||1|1||||4|4||||Yellow||Child/Family: Feels incompatible with volunteer|12.2||3|3|1|1|F|Black||11|No|Mother|28216|One Parent: Female|Unknown||Yes|TV|Media|General Community||Match Support|F|White||26|28262||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|502325039|31|0|2|503589790|1|0|2|500720750|2||-2||4|2|||-2||-2|56|1|||7464|9|||1|753584||4|3|45
503803127|BBBS of Greater Charlotte|Main Office|C|Active|2014-06-27|NaT|Baseline|2014-06-03|2014-06-27|Complete|Done|4|3|4|2|3|4|3.33|||||||||2|4|3|2|4|3|3|||||||||3|4|4|3.67||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|2|2|||||2|2||||4|4||||Green|||32.6||1|1|1|1|M|Black||14|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|Black||42|28270|Bachelors Degree|Married|Unknown||0|0|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500020910|503798593|31|0|1|503866013|31|0|1|500766041|2||-2||2|1|||-2||-2|0|4|||17101|1|||1|755946|-1|4|3|44
502582366|BBBS of Greater Charlotte|Main Office|C|Active|2014-06-30|NaT|Baseline|2014-06-12|2014-06-30|Complete|Done|1|2|2|1|2|4|2|||||||||1|1|3|2|2|3|2|||||||||4|4|4|4||||||4|3|5|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|||32.5||1|1|1|1|M|Black||13|No|Mother|28215|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community||Match Support|M|Black||31|28215|Some College|Single|Transport: Driver|28269|2|4|Local Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|502582874|31|0|1|503858870|31|0|1|500766366|2||-2||2|1|||-2||-2|0|10|||7437|1|||1|762956|-1|4|3|44
503879123|BBBS of Greater Charlotte|Main Office|C|Active|2014-06-21|NaT|Baseline|2014-06-12|2014-06-21|Complete|Done|2|1|4|4|2|4|2.83|||||||||4|3|4|4|4|4|3.83|||||||||4|4|4|4||||||4|4|4|3|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|3|2.5|||||2|2||||4|4||||Green|||32.8||1|1|1|1|M|Black||13|No|Mother|28212|One Parent: Female|$25,000 to $29,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28202|Masters Degree|Single|Finance: Banking|28244|0|3|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|503881119|31|0|1|503889097|1|0|1|500766443|2||-2||2|1|||-2||-2|34|2|||7464|9|||1|763180|-1|4|3|44
503492511|BBBS of Greater Charlotte|Main Office|C|Completed|2014-06-13|2015-02-05|Baseline|2014-06-13|2014-06-13|Complete|Done|4|1|2|1|4|4|2.67|||||||||1|4|3|3|1|4|2.67|||||||||4|4|4|4||||||5|2|4|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||1|1|1|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|7.8||1|1|1|1|M|Black||11|No|Mother|28216|One Parent: Female|$15,000 to $19,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||62|28210|Bachelors Degree|Divorced|Business: Engineer|28202|35|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503494379|31|0|1|503852376|1|0|1|500764721|2||-2||4|3|||-2||-2|34|2|||7464|9|||1|763762|-1|4|3|44
503686272|BBBS of Greater Charlotte|Main Office|C|Completed|2014-06-30|2016-04-18|Baseline|2014-06-18|2014-06-30|Complete|Done|4|2|1|1|1|4|2.17|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||3|1|5|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||4|1|2.5|||||2|2||||4|4||||Green||Volunteer: Lost contact with child/agency|21.6||1|1|1|1|M|Black||11|No|Mother|28216|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Enrollment|M|White||32|28210|Masters Degree|Single|Finance|28211|8|1|Recruitment Event|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|503688237|31|0|1|503817633|1|0|1|500766948|2||-2||4|1|||-2||-2|0|10|||7460|12|||1|765471|-1|4|3|44
503866348|BBBS of Greater Charlotte|Main Office|C|Active|2014-06-30|NaT|Baseline|2014-06-20|2014-06-30|Complete|Done|2|4|2|1|1|2|2|||||||||3|1|2|3|2|3|2.33|||||||||4|4|4|4||||||3|2|3|2|2.5|||||||4|4|4|3|4|4|4|3.86||||||||||3|2|3|2.67||||||4|4|4|||||1|1||||4|4||||Green|||32.5||1|1|1|1|M|Black||12|No|GrandMother|28216|Grandparents|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|M|White||45|28269|Bachelors Degree|Married|Finance: Banking|28273|1|0|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500008321|503838583|31|0|1|503862591|1|0|1|500767276|2||-2||2|1|||-2||-2|0|10|||17101|1|||1|766724|-1|4|3|44
503913977|BBBS of Greater Charlotte|Main Office|C|Completed|2014-06-24|2016-05-04|Baseline|2014-06-24|2014-06-24|Complete|Done|4|4|4|1|4|4|3.5|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||2|5|4|3|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||3|3||||Yellow||Child: Family structure changed|22.3||2|2|2|2|M|White||14|No|GrandMother|28031|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|M|White||61|28202|Masters Degree|Married|Retired||0|0|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|503915984|1|0|1|503898216|1|0|1|500767515|2||-2||4|2|||-2||-2|0|4|||17101|1|||1|767824|-1|4|3|44
503739899|BBBS of Greater Charlotte|Main Office|C|Active|2014-07-03|NaT|Baseline|2014-06-25|2014-07-03|Complete|Done|3|1|1|1|3|4|2.17|||||||||1|4|3|1|1|4|2.33|||||||||4|4|4|4||||||4|4|5|4|4.25|||||||4|4|4|3|4|4|3|3.71||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||32.4||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Insurance|28277|0|10|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020753|503702247|31|0|2|503802084|1|0|2|500767689|2||-2||2|1|||-2||-2|0|10|||7464|9|||1|768358|-1|4|3|44
503895740|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-28|2015-09-15|Baseline|2014-07-02|2014-08-27|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|3|4|3.83|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Yellow||Volunteer: Feels incompatible with child/family|12.6||2|2|1|1|F|Black||12|No|Mother|28273|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||34|28214|Some College|Single|Transport: Driver|28273|9|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500012459|503897736|31|0|2|503765053|31|0|2|500768490|2||-2||4|2|||-2||-2|0|10|||7464|9|||1|771599|-1|4|3|44
503880559|BBBS of Greater Charlotte|Main Office|C|Completed|2014-07-23|2014-09-04|Baseline|2014-07-03|2014-07-23|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green||Volunteer: Feels incompatible with child/family|1.4||1|1|2|2|F|Black||13|Yes|Father|28027|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Enrollment|F|Black||38|28269|Masters Degree|Single|Business|28262|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|277|60|598|500000170|500002335|503882555|31|0|2|503860995|31|0|2|500768591|2||-2||4|1|||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|771896|-1|4|1|44
503281015|BBBS of Greater Charlotte|Main Office|C|Completed|2013-11-25|2014-12-18|Followup|2014-11-25|2014-12-16|Complete|Done|3|3|3|3|3|3|3|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|3|2.5|||||2|2||||4|4||||Green||Child: Family structure changed|12.7||1|1|1|1|M|Black||11|No|Mother|28105|One Parent: Female|$30,000 to $34,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||45|28173|Bachelors Degree|Married|Finance|28277|13|5|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018987|503282834|31|0|1|503585313|1|0|1|500731009|2||-2||4|1|||-2||-2|34|2|||7464|9|||1|773040||4|3|45
503885975|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-01|2015-10-19|Baseline|2014-07-10|2014-08-01|Complete|Done|3|3|4|1|4|4|3.17|||||||||3|4|3|3|1|3|2.83|||||||||4|3|4|3.67||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||1|1|1|||||2|2||||4|4||||Red||Volunteer: Moved|14.6||2|2|1|1|M|Black||12|No|Mother|28216|One Parent: Female|$45,000 to $49,999||No||Relative|General Community||Match Support|M|White||28|28262|Associate Degree|Single|Finance: Banking|28081|1|1|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500017777|503887971|31|0|1|503885544|1|0|1|500769090|2||-2||4|3|||-2||-2|0|3|||17101|1|||1|773442|-1|4|3|44
503810996|BBBS of Greater Charlotte|Main Office|C|Active|2014-07-31|NaT|Baseline|2014-07-11|2014-07-31|Complete|Done|3|3|4|1|3|4|3|||||||||2|2|4|2|1|4|2.5|||||||||4|4|4|4||||||5|2|3|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||2|2||||4|4||||Green|||31.5||1|1|1|1|M|Black||12|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|Black||63|28078|Bachelors Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|503812973|31|0|1|503799211|31|0|1|500769226|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||7671|13|||1|773759|-1|4|3|44
503743876|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-10|2016-08-01|Baseline|2014-07-11|2014-09-10|Complete|Done|4|1|2|1|2|4|2.33|||||||||1|2|3|3|2|4|2.5|||||||||4|2|3|3||||||4|5|3|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green||Child/Family: Moved|22.7||1|1|1|1|M|Black||13|No|Mother|28212|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Enrollment|M|White||44|28203|Masters Degree|Single|Finance|29715|10|0|Igniting Breakfast|Special Event|Big|General Community||Match Support|277|60|598|500000170|500020752|503261158|31|0|1|503908096|1|0|1|500769242|2||-2||4|1|||-2||-2|0|10|||17266|8|||1|773786|-1|4|3|44
502602926|BBBS of Greater Charlotte|Main Office|C|Active|2014-08-05|NaT|Baseline|2014-07-14|2014-08-05|Complete|Done|3|3|4|3|4|4|3.5|||||||||3|4|3|4|4|4|3.67|||||||||4|4|3|3.67||||||3|5|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||2|1|1.5|||||2|2||||4|4||||Green|||31.3||1|1|1|1|F|Black||11|No|Mother|28216|One Parent: Female|$25,000 to $29,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Some Other Race||30|28214|Bachelors Degree|Married|Business|28214|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500013781|502603443|31|0|2|503808719|41|0|2|500769460|2||-2||2|1|||-2||-2|6854|8|||7462|13|||1|774377|-1|4|3|44
503331975|BBBS of Greater Charlotte|Main Office|C|Completed|2014-07-25|2014-11-06|Baseline|2014-07-14|2014-07-23|Complete|Done|1|4|4|4|3|2|3|||||||||4|3|3|4|4|4|3.67|||||||||4|2|4|3.33||||||3|4|4|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||3|3|3|||||1|1||||4|4||||Red||Child: Lost interest|3.4||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||34|28269|Bachelors Degree|Married|Medical: Healthcare Worker|28209|0|4|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500012459|503333815|31|0|2|503796877|31|0|2|500769464|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|774384|-1|4|3|44
503899239|BBBS of Greater Charlotte|Main Office|C|Completed|2014-07-30|2017-01-26|Baseline|2014-07-21|2014-07-30|Complete|Done|4|3|4|3|3|4|3.5|||||||||2|3|4|3|3|3|3|||||||||3|3|3|3||||||3|4|4|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||4|4||||Green||Child/Family: Feels incompatible with volunteer|29.9||1|1|1|1|M|Black||15|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||38|28269|Some College|Married|Tech: Management|28273|3|1|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500021785|503901239|31|0|1|503871007|1|0|1|500770094|2||-2||4|1|||-2||-2|0|10|||17101|1|||1|776024|-1|4|3|44
503834613|BBBS of Greater Charlotte|Main Office|C|Completed|2014-07-29|2015-03-05|Baseline|2014-07-22|2014-07-29|Complete|Done|3|4|2|3|3|3|3|||||||||2|4|3|4|2|3|3|||||||||4|4|4|4||||||3|4|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|3|3|3.33||||||3|2|2.5|||||1|1||||4|4||||Yellow||Volunteer: Time constraint|7.2||1|1|1|1|M|White||15|No|Mother|28226|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community||RTBM|M|White||73|28277|High School Graduate|Married|Arts, Entertainment, Sports||0|0|Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500012459|503836592|1|0|1|503790527|1|0|1|500770182|2||-2||4|2|||-2||-2|0|10|||131|1|||1|776269|-1|4|3|44
503746685|BBBS of Greater Charlotte|Main Office|C|Completed|2014-11-17|2016-07-29|Baseline|2014-07-24|2014-11-17|Complete|Done|4|3|4|2|4|4|3.5|||||||||3|3|4|1|4|4|3.17|||||||||4|3|3|3.33||||||4|4|4|4|4|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Lost contact with child/agency|20.4||1|1|1|1|F|Black||16|No|Mother|28277|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||31|28209|Juris Doctorate (JD)|Single|Law|28210|1|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|503755760|31|0|2|503961087|1|0|2|500790718|2||-2||4|3|500014681|500014681|-2|500014681|-2|34|2|||17159|12|||1|776943|-1|4|3|44
502943644|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-25|2015-10-30|Baseline|2014-08-06|2014-08-25|Complete|Done|2|4|4|4|2|4|3.33|||||||||2|4|3|1|2|2|2.33|||||||||4|4|4|4||||||3|4|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|14.2||2|2|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999||Yes||Self|General Community||Match Support|F|Black||23|28213||Single|Arts, Entertainment, Sports||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|502945070|31|0|2|503899413|31|0|2|500771637|2||-2||4|3|||-2||-2|0|10|||7464|9|||1|783186|-1|4|3|44
502068488|BBBS of Greater Charlotte|Main Office|C|Active|2014-08-26|NaT|Baseline|2014-08-11|2014-08-26|Complete|Done|2|1|1|1|4|1|1.67|||||||||3|2|4|1|1|2|2.17|||||||||4|3|4|3.67||||||4|2|5|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|Cabarrus County||30.7||1|1|1|1|M|White||12|No|Mother|28269|One Parent: Female|$60,000 to $74,999||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|White||35|28075|Masters Degree|Single|Finance: Accountant|28202|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|502068912|1|0|1|503953186|1|0|1|500771917|2||500016307||2|1|500016374|500016374|-2|500016374|-2|6854|8|||7464|9|||1|784072|-1|4|3|44
503569115|BBBS of Greater Charlotte|Main Office|C|Completed|2013-12-19|2015-03-19|Followup|2014-12-19|2015-01-15|Complete|Done|3|2|1|4|1|3|2.33|||||||||2|4|4|1|2|3|2.67|||||||||3|4|4|3.67||||||1|3|1|1|1.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|3|3.5|||||2|2||||4|4||||Green||Child/Family: Moved|14.9||1|1|1|1|F|Black||11|No|Mother|2649|One Parent: Female|Unknown||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Education: Teacher|28012|3|0|Self|Self|Big|General Community||Enrollment|277|60|598|500000170|500015820|503570990|31|0|2|503619714|1|0|2|500735248|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|784233||4|3|45
503941222|BBBS of Greater Charlotte|Main Office|C|Active|2014-08-29|NaT|Baseline|2014-08-12|2014-08-29|Complete|Done|4|4|4|1|2|4|3.17|||||||||3|4|4|4|3|4|3.67|||||||||4|4|4|4||||||2|5|2|2|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|3|4|3.67||||||3|3|3|||||2|2||||4|4||||Yellow|||30.6||1|1|1|1|F|Black||12|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|White||28|28205|Masters Degree|Single|Business: Mgt, Admin|28262|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|503931754|31|0|2|503889588|1|0|2|500772492|2||-2||2|2|||-2||-2|0|4|||17159|12|||1|784292|-1|4|3|44
503700282|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-27|2014-12-23|Baseline|2014-08-12|2014-08-27|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|2|4|3.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green||Volunteer: Time constraint|3.9||1|1|1|1|M|Black||13|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|M|Black||42|28214|Some College|Domestic Partner|Service: Restaurant|28208|8|6|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500018987|503702247|31|0|1|503874948|31|0|1|500771987|2||-2||4|1|||-2||-2|0|10|||17101|1|||1|784298|-1|4|3|44
503929747|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-29|2016-07-29|Baseline|2014-08-12|2014-08-29|Complete|Done|3|4|4|4|2|4|3.5|||||||||1|4|3|3|2|3|2.67|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|23||1|1|1|1|F|Black||12|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Multi-race (Asian & White)||28|28203|Bachelors Degree|Single|Finance|28211|0|4|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|503931754|31|0|2|503910740|37|0|2|500772491|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|784301|-1|4|3|44
503796616|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-25|2015-10-20|Baseline|2014-08-12|2014-08-25|Complete|Done|3|1|1|1|3|4|2.17|||||||||2|3|4|2|2|4|2.83|||||||||3|4|3|3.33||||||3|2|4|3|3|||||||3|4|3|4|4|4|4|3.71||||||||||3|2|3|2.67||||||3|4|3.5|||||1|1||||4|4||||Green||Volunteer: Time constraint|13.8||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||30|28273|Bachelors Degree|Single|Business: Human Resources|28203|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500018987|503798593|31|0|2|503828896|1|0|2|500772098|2||-2||4|1|||-2||-2|0|10|||7496|10|||1|784433|-1|4|3|44
503937201|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-22|2015-12-09|Baseline|2014-08-13|2014-08-22|Complete|Done|4|1|4|1|4|4|3|||||||||3|4|4|2|1|4|3|||||||||4|4|4|4||||||3|4|3|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|4|3.67||||||3|3|3|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|15.6||1|1|1|1|F|Black||14|No|Mother|28031|Two Parent|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||49|28115|High School Graduate|Single|Customer Service|28115|13|1|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503939209|31|0|2|503582646|1|0|2|500772180|2||-2||4|3|||-2||-2|0|4|||7464|9|||1|784654|-1|4|3|44
503831166|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-21|2016-01-26|Baseline|2014-08-13|2014-08-21|Complete|Done|2|3|2|3|1|2|2.17|||||||||3|4|4|3|3|3|3.33|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Green||Volunteer: Time constraint|17.2||1|1|1|1|M|Black||15|No|Mother|28227|One Parent: Female|$60,000 to $74,999||No|AARTF|BBBS Board/Staff|General Community||Match Support|M|Black||23|28227|Some College|Single|Student: College|28078|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|277|60|598|500000170|500020752|503833145|31|0|1|503861120|31|0|1|500772203|2||-2||4|1|||-2||-2|7294|13|||7496|10|||1|784689|-1|4|3|44
503952645|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-22|NaT|Baseline|2014-08-18|2014-10-22|Complete|Done|3|4|3|4|3|4|3.5|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||5|5|4|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||28.8||1|1|1|1|F|White||14|No|Father|28025|One Parent: Male|$40,000 to $44,999|Y|No|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||31|28025|Bachelors Degree|Married|Business: Mgt, Admin|28027|4|7|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|503954653|1|0|2|503942996|31|0|2|500772607|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|34|2|||7464|9|||1|785703|-1|4|3|44
503532788|BBBS of Greater Charlotte|Main Office|C|Active|2014-08-23|NaT|Baseline|2014-08-18|2014-08-22|Complete|Done|3|4|4|1|4|3|3.17|||||||||2|3|2|3|2|3|2.5|||||||||4|4|4|4||||||3|4|2|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Green|Cabarrus County||30.8||1|1|1|1|F|Black||15|Yes|GrandMother|28075|Grandparents|$10,000 to $14,999|Y|Yes||Relative|General Community|Amachi, Cabarrus County|Match Support|F|Black||33|28269|PHD|Single|Education: Admin|28081|4|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|277|60|598|500000170|500022817|503534663|31|0|2|503939365|31|0|2|500772617|2||500016307||2|1|500016374|500000294, 500016374|-2|500016374|-2|0|3|||17159|12|||1|785713|-1|4|3|44
503838769|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-30|2015-09-16|Baseline|2014-08-20|2014-08-30|Complete|Done|3|3|4|2|4|3|3.17|||||||||3|3|3|3|3|3|3|||||||||4|3|3|3.33||||||3|4|2|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|1|2|||||2|2||||4|4||||Red||Child/Family: Moved|12.6||1|1|1|1|M|Black||14|No|Mother|28269|One Parent: Female|$25,000 to $29,999||No||Self|General Community||Match Support|M|Black||62|28210|Bachelors Degree|Divorced|Business|28202|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|277|60|598|500000170|500008321|503840748|31|0|1|503948333|31|0|1|500772925|2||-2||4|3|||-2||-2|0|10|||7671|13|||1|786363|-1|4|3|44
503898651|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-17|2016-02-29|Baseline|2014-08-21|2014-09-17|Complete|Done|3|4|2|1|3|4|2.83|||||||||2|3|3|4|3|3|3|||||||||4|4|4|4||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Child/Family: Lost contact with volunteer/agency|17.4||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||40|28056|Some College|Single|Real Estate: Realtor|28202|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|503891857|31|0|2|503494199|31|0|2|500773073|2||-2||4|3|||-2||-2|0|10|||46|2|||1|786597|-1|4|3|44
503930457|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-30|2014-12-23|Baseline|2014-08-21|2014-08-30|Complete|Done|4|1|2|1|4|4|2.67|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||1|1||||4|4||||Green||Child/Family: Moved|3.8||1|1|1|1|F|Black||12|No|Mother|28217|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Match Support|F|White||46|28226|Masters Degree|Married|Self-Employed, Entrepreneur|28277|16|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|503932464|31|0|2|503544824|1|0|2|500773041|2||-2||4|1|||-2||-2|0|10|||46|2|||1|786603|-1|4|3|44
503813942|BBBS of Greater Charlotte|Main Office|C|Completed|2014-08-30|2017-02-28|Baseline|2014-08-21|2014-08-30|Complete|Done|3|3|4|1|3|4|3|||||||||4|1|4|4|4|4|3.5|||||||||4|3|4|3.67||||||4|3|5|5|4.25|||||||4|4|4|4|4|3|3|3.71||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|30||1|1|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community||Match Support|M|Black||38|28269||Single|Unemployed||0|0|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500020752|503815919|31|0|1|503873603|31|0|1|500773055|2||-2||4|1|||-2||-2|0|3|||17101|1|||1|786621|-1|4|3|44
503804225|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-15|2016-01-29|Baseline|2014-08-21|2014-09-15|Complete|Done|3|3|3|2|3|3|2.83|||||||||2|3|3|3|1|3|2.5|||||||||4|4|4|4||||||2|5|4|4|3.75|||||||4|4|4|4|3|3|3|3.57||||||||||2|3|1|2||||||4|2|3|||||1|1||||4|4||||Red||Volunteer: Lost contact with child/agency|16.5||1|1|1|1|F|Black||17|No|Mother|28208|One Parent: Female|$25,000 to $29,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Multi-race (Black & Hispanic)||59|28216|Some College|Divorced|Law: Legal Secretary|28202|14|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500013781|503805695|31|0|2|503881040|38|0|2|500773105|2||-2||4|3|||-2||-2|34|2|||7464|9|||1|786691|-1|4|3|44
503959684|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-15|2015-10-29|Baseline|2014-08-26|2014-09-15|Complete|Done|3|1|4|1|3|4|2.67|||||||||4|4|3|3|4|3|3.5|||||||||4|4|4|4||||||4|5|4|2|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green||Child/Family: Moved|13.4||1|1|1|1|F|Black||13|No|Mother|28227|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||26|28207|Masters Degree||Finance: Accountant|28202|0|11|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017777|503961693|31|0|2|503985328|1|0|2|500775400|2||-2||4|1|||-2||-2|0|10|||7464|9|||1|787764|-1|4|3|44
502612404|BBBS of Greater Charlotte|Main Office|C|Completed|2014-10-06|2015-05-27|Baseline|2014-08-28|2014-10-06|Complete|Done|3|1|4|4|3|4|3.17|||||||||4|3|4|2|1|4|3|||||||||4|3|3|3.33||||||5|4|4|4|4.25|||||||4|4|4|4|3|4|2|3.57||||||||||3|4|1|2.67||||||1|1|1|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Moved|7.7||2|2|1|1|F|Some Other Race||15|No|Aunt|28217|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||26|28217|Bachelors Degree|Single|Business|28277|0|8|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|500188044|41|0|2|503790988|31|0|2|500773744|2||-2||4|3|500014681||-2|500014681|-2|0|10|||46|2|||1|788378|-1|4|3|44
503535102|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-17|2015-05-14|Baseline|2014-09-02|2014-09-17|Complete|Done|4|2|2|1|3|4|2.67|||||||||2|3|3|2|2|4|2.67|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Yellow||Volunteer: Lost contact with child/agency|7.9||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28217|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Enrollment|F|Black||26|28214|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|503536977|36|0|2|503882165|31|0|2|500774003|2||-2||4|2|||-2||-2|0|10|||46|2|||1|789389|-1|4|3|44
503851354|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-29|2015-10-30|Baseline|2014-09-04|2014-09-29|Complete|Done|3|3|4|4|4|4|3.67|||||||||3|1|4|2|3|3|2.67|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||2|4|4|3.33||||||2|1|1.5|||||1|1||||4|4||||Red||Volunteer: Moved|13||1|1|1|1|M|Black||13|Yes|Mother|28227|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||34|28209|Masters Degree|Single|Finance: Accountant|28210|2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|503853343|31|0|1|503962684|1|0|1|500774775|2||-2||4|3|||-2|500000294|-2|0|10|||46|2|||1|790002|-1|4|3|44
503546374|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-29|2015-03-26|Baseline|2014-09-04|2014-09-29|Complete|Done|3|4|4|4|4|2|3.5|||||||||4|3|4|3|2|3|3.17|||||||||4|2|2|2.67||||||3|3|2|5|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|2|2.67||||||3|3|3|||||1|1||||4|4||||Yellow|PERL 2014-2016|Child: Severity of challenges|5.8||1|1|2|2|M|Black||17|No|Mother|28216|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Asian||33|28204|Bachelors Degree|Married|Business: Engineer|28007|3|9|Man Up Campaign|Media|Big|General Community|Amachi, PERL 2014-2016|Match Support|277|60|598|500000170|500015820|503548249|31|0|1|503890372|4|0|1|500774577|2||-2||4|2|500014681|500014681|-2|500000294, 500014681|-2|0|4|||17101|1|||1|790147|-1|4|3|44
503544893|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-26|2015-10-06|Baseline|2014-09-08|2014-09-26|Complete|Done|4|1|2|2|2|4|2.5|||||||||2|2|4|3|2|4|2.83|||||||||4|4|4|4||||||3|2|4|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|12.3||1|1|2|2|F|Black||14|No|Mother|28227|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community||Match Support|F|Black||46|28216|Bachelors Degree|Single|Business: Marketing|28036|0|3|Self|Self|Big|General Community|VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500012459|503546768|31|0|2|503844843|31|0|2|500777054|2||-2||4|2|||-2|500007920, 500011312, 500011315, 500011316|-2|0|10|||7464|9|||1|790639|-1|4|3|44
503628199|BBBS of Greater Charlotte|Main Office|C|Completed|2014-09-18|2015-03-06|Baseline|2014-09-09|2014-09-18|Complete|Done|4|2|4|1|3|4|3|||||||||3|4|4|4|4|4|3.83|||||||||1|1|1|1||||||5|5|5|4|4.75|||||||4|4|4|4|3|4|1|3.43||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|5.6||1|1|1|1|M|Black||13|No|Mother|28273|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||54|28226|Masters Degree|Single|Tech: Computer/Programmer|28202|0|3|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503630137|31|0|1|503966130|1|0|1|500775002|2||-2||4|1||500014681|-2|500000294|-2|0|10|||17159|12|||1|790992|-1|4|3|44
503953654|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-10|NaT|Baseline|2014-09-11|2014-10-10|Complete|Done|3|1|4|1|3|3|2.5|||||||||1|4|3|2|3|3|2.67|||||||||3|4|3|3.33||||||3|4|5|2|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|4|3.33||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016||29.2||1|1|1|1|M|Black||14|Yes|Mother|28208|One Parent: Female|Less than $10,000|Y|No||Therapist/Counselor|General Community|Amachi, PERL 2014-2016|Match Support|M|White||28|28209|Bachelors Degree|Single|Tech: Engineer||0|5|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503955662|31|0|1|503976139|1|0|1|500775808|2||-2||2|1|500014681|500000294, 500014681|-2|500014681|-2|0|5|||46|2|||1|791743|-1|4|3|44
503704573|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-08|NaT|Baseline|2014-09-18|2014-10-08|Complete|Done|3|2|3|1|3|2|2.33|||||||||3|3|3|2|3|3|2.83|||||||||4|4|4|4||||||3|5|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016||29.2||1|1|1|1|M|Black||15|No|Mother|28273|One Parent: Female|$20,000 to $24,999||No||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28277|Bachelors Degree|Single|Business: Marketing|29067|0|3|Man Up Campaign|Media|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|503706538|31|0|1|503883049|1|0|1|500776636|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||17101|1|||1|793510|-1|4|3|44
503833936|BBBS of Greater Charlotte|Main Office|C|Active|2014-09-28|NaT|Baseline|2014-09-18|2014-09-28|Complete|Done|2|3|3|2|3|2|2.5|||||||||4|3|3|4|4|4|3.67|||||||||4|4|4|4||||||2|3|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|||29.6||1|1|1|1|M|Multi-race (Asian & White)||13|No|Mother|28078|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Married|Unemployed|28031|6|2|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018851|503835915|37|0|1|502489398|1|0|1|500776719|2||-2||2|1|||-2||-2|0|10|||46|2|||1|793575|-1|4|3|44
503723888|BBBS of Greater Charlotte|Main Office|C|Completed|2014-10-13|2015-12-02|Baseline|2014-09-18|2014-10-13|Complete|Done|1|2|4|1|4|4|2.67|||||||||3|4|3|3|2|4|3.17|||||||||4|4|4|4||||||5|2|2|5|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Time constraint|13.6||1|1|1|1|M|Black||11|Yes|Mother|28215|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community||Enrollment|M|Black||26|28227|Bachelors Degree|Single|Customer Service||1|3|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|503725860|31|0|1|503858682|31|0|1|500779634|2||-2||4|3|||-2||-2|0|10|||17101|1|||1|793585|-1|4|3|44
503849038|BBBS of Greater Charlotte|Main Office|C|Completed|2014-10-15|2015-12-28|Baseline|2014-09-29|2014-10-15|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|3|4|2|3|3|||||||||4|4|4|4||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|2|3|||||1|1||||4|4||||Green||Volunteer: Lost contact with child/agency|14.4||1|1|1|1|M|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999||No||Self|General Community||Match Support|M|Black||32|28202|Bachelors Degree|Single|Consultant|28202|0|9|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|503851023|31|0|1|503930671|31|0|1|500778856|2||-2||4|1|||-2||-2|0|10|||17101|1|||1|796933|-1|4|3|44
503923102|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-13|NaT|Baseline|2014-10-01|2014-10-13|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|2|3|4|3.33|||||||||4|4|4|4||||||4|5|5|5|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||29.1||1|1|1|1|M|Black||17|No|Mother|28213|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|M|Black||48|28262||Single|Retired||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|503925109|31|0|1|503996589|31|0|1|500781196|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|798208|-1|4|3|44
503723868|BBBS of Greater Charlotte|Main Office|C|Completed|2014-10-13|2015-10-15|Baseline|2014-10-01|2014-10-13|Complete|Done|4|4|4|3|4|4|3.83|||||||||4|4|4|2|4|4|3.67|||||||||4|4|4|4||||||5|3|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red||Volunteer: Moved|12.1||1|1|1|1|M|Black||13|Yes|Mother|28215|One Parent: Female|$10,000 to $14,999||Yes||Self|General Community||Enrollment|M|Black||25|28205|Bachelors Degree|Single|Tech: Research/Design|28202|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|503725860|31|0|1|503940354|31|0|1|500779635|2||-2||4|3|||-2||-2|0|10|||17159|12|||1|798237|-1|4|3|44
503972507|BBBS of Greater Charlotte|Main Office|C|Completed|2014-10-13|2017-02-27|Baseline|2014-10-03|2014-10-13|Complete|Done|2|4|4|1|3|4|3|||||||||2|4|4|4|2|4|3.33|||||||||4|4|4|4||||||4|3|5|3|3.75|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||2|4|3|||||1|1||||4|4||||Green||Volunteer: Time constraint|28.5||1|1|2|2|F|Black||14|Yes|Mother|28278|One Parent: Female|$50,000 to $59,999|Y|No||Self|General Community||Match Support|M|Black||46|28214|Bachelors Degree|Single|Finance: Economist|28217|14|0|Brochure|Media|Big|General Community||Match Support|277|60|598|500000170|500013781|503974518|31|0|2|500189600|31|0|1|500780309|2||500003586||4|1|||-2||-2|0|10|||127|1|||1|799000|-1|4|3|44
503869451|BBBS of Greater Charlotte|Main Office|C|Completed|2014-10-27|2014-12-30|Baseline|2014-10-13|2014-10-27|Complete|Done|2|2|1|3|1|2|1.83|||||||||2|1|2|1|3|2|1.83|||||||||3|4|4|3.67||||||3|3|5|2|3.25||||||||3|4|4|3|3|3|||||||||||3|3|3|3||||||1|4|2.5|||||2|2||||4|4||||Green||Volunteer: Moved|2.1||2|2|1|1|F|White||13|No|Mother|28212|Two Parent|Less than $10,000|Y|Yes||Therapist/Counselor|General Community||Enrollment|F|White||30|28205|Masters Degree|Single|Business|28201|2|3|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500017777|503871445|1|0|2|503940385|1|0|2|500783066|2||-2||4|1|||-2||-2|0|5|||46|2|||1|802598|-1|4|3|44
504004117|BBBS of Greater Charlotte|Main Office|C|Active|2014-11-10|NaT|Baseline|2014-10-13|2014-11-10|Complete|Done|3|4|4|3|3|3|3.33|||||||||4|4|4|4|1|4|3.5|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||28.2||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||26|28269|Masters Degree|Single|Human Services: Social Worker|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504006132|31|0|2|503929259|31|0|2|500783097|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|802635|-1|4|3|44
503803718|BBBS of Greater Charlotte|Main Office|C|Active|2014-11-13|NaT|Baseline|2014-10-13|2014-11-13|Complete|Done|4|4|4|1|4|4|3.5|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|5|5|4|4.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2|||||||||Green|||28.1||1|1|1|1|M|Black||15|No|Mother|28208|One Parent: Female|$20,000 to $24,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Some Other Race||33|28056|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28204|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|503805695|31|0|1|503930530|41|0|1|500783205|2||-2||2|1|||-2||-2|34|2|||46|2|||1|802744|-1|4|3|44
503895506|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-21|NaT|Baseline|2014-10-15|2014-10-21|Complete|Done|2|4|4|3|4|4|3.5|||||||||3|4|4|3|3|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016||28.8||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28212|Two Parent|Unknown|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||30|28226||Single|Unemployed||0|0|Relative|Relative|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|503897502|3|10|2|504026849|3|0|2|500784082|2||-2||2|1|500011312, 500014681|500014681|-2|500014681|-2|0|4|||17161|11|||1|803884|-1|4|3|44
504031334|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-29|NaT|Baseline|2014-10-23|2014-10-29|Complete|Done|3|3|3|2|3|3|2.83|||||||||3|3|4|3|3|4|3.33|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|3|2.5|||||1|1||||4|4||||Green|||28.6||1|1|1|1|F|Black||15|No|Mother|28262|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||37|28208|Bachelors Degree|Single|Tech: Research/Design|28202|3|8|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500018851|503917391|31|0|2|503882331|1|0|2|500787330|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|808164|-1|4|3|44
503915384|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-26|NaT|Baseline|2014-10-23|2014-10-26|Complete|Done|3|3|3|3|3|3|3|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|2|2|3|2.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|3|3|||||1|1||||4|4||||Green|PERL 2014-2016||28.6||1|1|1|1|M|Black||13|No|Mother|28262|One Parent: Female|$20,000 to $24,999||Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|Multi-race (Asian & White)||36|28203|Masters Degree|Married|Finance: Banking|20815|11|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500018851|503917391|31|0|1|503995835|37|0|1|500787470|2||-2||2|1|500014681|500014681|-2|500014681|-2|34|2|||7464|9|||1|808387|-1|4|3|44
503831971|BBBS of Greater Charlotte|Main Office|C|Completed|2014-11-17|2015-06-30|Baseline|2014-10-27|2014-11-17|Complete|Done|3|3|3|4|3|4|3.33|||||||||2|3|3|2|3|3|2.67|||||||||4|3|3|3.33||||||3|3|3|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||2|4|3|||||2|2||||4|4||||Yellow||Child/Family: Lost contact with volunteer/agency|7.4||1|1|2|2|M|Black||15|Yes|Mother|28269|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Amachi|Match Support|M|Hispanic||31|28209|High School Graduate|Single|Finance|28262|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500012459|503833950|31|0|1|504011759|3|0|1|500788190|2||-2||4|2||500000294|-2||-2|0|10|||46|2|||1|809554|-1|4|3|44
503961917|BBBS of Greater Charlotte|Main Office|C|Active|2014-10-31|NaT|Baseline|2014-10-27|2014-10-31|Complete|Done|1|2|2|2|2|2|1.83|||||||||4|2|4|2|3|3|3|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||28.5||1|1|1|1|M|White||14|No|Father|28081|One Parent: Male|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||28|28277|Bachelors Degree||Finance|28255|0|4|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503636659|1|0|1|504052039|1|0|1|500788399|2||-2||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|5|||17159|12|||1|809764|-1|4|3|44
503995803|BBBS of Greater Charlotte|Main Office|C|Completed|2014-11-24|2015-10-01|Baseline|2014-10-30|2014-11-24|Complete|Done|1|2|2||1|1||||||||||2|2|3|2|4|3|2.67|||||||||4|4|4|4||||||4|2|4|4|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Time constraint|10.2||1|1|1|1|F|Black||12|No|Mother|28206|Two Parent|$10,000 to $14,999|Y|Yes||Relative|General Community|PERL 2014-2016|Match Support|F|Black||44|28269||Single|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|503997818|31|0|2|503963125|31|0|2|500790223|2||-2||4|3|500014681|500014681|-2|500014681|-2|0|3|||17159|12|||1|812296|-1|4|3|44
503983132|BBBS of Greater Charlotte|Main Office|C|Active|2014-11-17|NaT|Baseline|2014-11-03|2014-11-17|Complete|Done|4|4|4|1|4|4|3.5|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|2|4|3|3.57||||||||||4|4|4|4||||||1|4|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||27.9||1|1|1|1|M|Black||16|Yes|GrandMother|28270|One Parent: Female|$15,000 to $19,999|Y|No||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||49|28226|Juris Doctorate (JD)|Married|Law: Lawyer|28202|4|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|503985143|31|0|1|503995895|1|0|1|500791249|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|5|||46|2|||1|814090|-1|4|3|44
503552606|BBBS of Greater Charlotte|Main Office|C|Active|2014-11-21|NaT|Baseline|2014-11-12|2014-11-21|Complete|Done|4|4|4|4|4|4|4|||||||||3|3|4|4|4|4|3.67|||||||||4|4|4|4||||||5|4|3|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|4|3|||||1|1||||4|4||||Green|||27.8||1|1|2|2|M|Black||14|No|Mother|28079|One Parent: Female|Unknown||No||Self|General Community||Match Support|M|Black||45|28079|Bachelors Degree|Married|Business||13|6|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|277|60|598|500000170|500017732|503554481|31|0|1|501052547|31|0|1|500794702|2||-2||2|1|||-2|500000294|-2|0|10|||7671|13|||1|818843|-1|4|3|44
504085882|BBBS of Greater Charlotte|Main Office|C|Completed|2014-11-21|2017-02-28|Baseline|2014-11-12|2014-11-21|Complete|Done|3|1|4|2|4|4|3|||||||||3|4|4|4|2|3|3.33|||||||||4|4|4|4||||||5|4|4|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||3|3|2|2.67||||||2|4|3|||||2|2||||4|4||||Red|PERL 2014-2016|Child/Family: Time constraints|27.3||1|1|1|1|F|Black||16|No|GrandMother|28269|One Parent: Female|Unknown|Y|Yes||Foster Home|General Community|PERL 2014-2016|Match Support|F|Black||24|28217|Bachelors Degree|Single|Finance||0|2|AA Task Force|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|503144847|31|0|2|503977000|31|0|2|500794719|2||-2||4|3|500014681|500014681|-2|500014681|-2|0|7|||9229|13|||1|818859|-1|4|3|44
504059280|BBBS of Greater Charlotte|Main Office|C|Completed|2014-12-16|2016-08-29|Baseline|2014-11-15|2014-12-16|Complete|Done|3|4|4|1|3|4|3.17|||||||||2|3|4|4|2|4|3.17|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|3|3.33||||||4|3|3.5|||||1|1||||4|4||||Red|VOL - Mentoring Hispanic Youth|Child: Family structure changed|20.4||1|1|1|1|M|Hispanic|Other Central American|13|No|Mother|28214|One Parent: Female|Unknown|Y|Yes||Therapist/Counselor|General Community|VOL - Mentoring Hispanic Youth|Match Support|M|Hispanic||37|28078|Associate Degree|Single|Finance|28217|0|3|Coworker|Workplace Partner|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|277|60|598|500000170|500017777|504061304|3|14|1|503998203|3|0|1|500796014|2||-2||4|3|500011312|500011312|-2|500011312|-2|0|5|||7447|3|||1|820730|-1|4|3|44
504081573|BBBS of Greater Charlotte|Main Office|C|Completed|2014-11-25|2015-09-17|Baseline|2014-11-15|2014-11-25|Complete|Done|4|4|4|4|4|4|4|||||||||4|4|4|4|4|4|4|||||||||4|4|4|4||||||5|2|5|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green||Volunteer: Moved|9.7||2|2|1|1|F|Black||14|No|Mother|28206|One Parent: Female|Unknown|Y|No||Relative|General Community||Enrollment|F|White||27|28278|Bachelors Degree|Single|Education: Teacher|28056|1|9|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017777|501091694|31|0|2|503880925|1|0|2|500796131|2||-2||4|1|||-2||-2|0|3|||17159|12|||1|820734|-1|4|3|44
503873575|BBBS of Greater Charlotte|Main Office|C|Completed|2014-11-24|2015-10-22|Baseline|2014-11-17|2014-11-24|Complete|Done|4|3|3|3|2|4|3.17|||||||||2|4|3|2|2|4|2.83|||||||||4|4|4|4||||||2|4|5|5|4|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|2|2.67||||||3|2|2.5|||||2|2||||4|4||||Green||Child/Family: Moved|10.9||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||39|28078|Bachelors Degree|Single|Business: Sales|28117|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500018987|503875571|31|0|2|504004351|1|0|2|500796129|2||-2||4|1|||-2||-2|0|10|||46|2|||1|821002|-1|4|3|44
503934189|BBBS of Greater Charlotte|Main Office|C|Active|2014-11-25|NaT|Baseline|2014-11-17|2014-11-25|Complete|Done|2|4|2|4|3|2|2.83|||||||||2|3||3|3|3||||||||||4|3|4|3.67||||||4|3|4|3|3.5|||||||4|4|4|4|4|3|3|3.71||||||||||3|4|3|3.33||||||2|3|2.5|||||2|2||||4|4||||Green|||27.7||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|M|White||35|28211|Masters Degree|Single|Finance: Accountant|28202|2|0|Man Up Campaign|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|503936197|31|0|1|503918487|1|0|1|500796401|2||-2||2|1|||-2||-2|0|4|||17101|1|||1|821302|-1|4|3|44
503978153|BBBS of Greater Charlotte|Main Office|C|Active|2014-12-15|NaT|Baseline|2014-11-21|2014-12-15|Complete|Done|4|1|1|1|3|4|2.33|||||||||1|2|3|2|3|3|2.33|||||||||4|4|4|4||||||2|3|4|4|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Green|PERL 2014-2016||27||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||37|28227|Associate Degree|Single|Student: College|28223|1|0|Web in a Box, v1|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|503980164|31|0|2|504039547|31|0|2|500798168|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||15467|2|||1|823862|-1|4|3|44
503989203|BBBS of Greater Charlotte|Main Office|C|Active|2014-12-15|NaT|Baseline|2014-11-26|2014-12-15|Complete|Done|3|3|4|3|2|2|2.83|||||||||2|3|3|2|4|3|2.83|||||||||4|4|4|4||||||2|4|4|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|PERL 2014-2016||27||1|1|1|1|M|White||13|No|Mother|28216|One Parent: Female|$35,000 to $39,999|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28203|Bachelors Degree|Single|Finance: Banking|28203|7|8|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|503991217|1|0|1|504066226|1|0|1|500799476|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|5|||17159|12|||1|826224|-1|4|3|44
504038458|BBBS of Greater Charlotte|Main Office|C|Active|2014-12-16|NaT|Baseline|2014-12-02|2014-12-16|Complete|Done|3|1|4|1|1|2|2|||||||||2|4|3|3|2|3|2.83|||||||||4|4|4|4||||||3|5|5|1|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|||27||1|1|1|1|F|Black||12|No|Mother|28216|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|White||25|28209|Bachelors Degree|Single|Finance|28202|1|3|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|277|60|598|500000170|500020752|504040320|31|0|2|503971368|1|0|2|500800323|2||-2||2|1|||-2|500000294|-2|0|10|||17159|12|||1|827870|-1|4|3|44
503977573|BBBS of Greater Charlotte|Main Office|C|Completed|2014-12-29|2015-11-30|Baseline|2014-12-04|2014-12-29|Complete|Done|4|2|1|1|3|3|2.33|||||||||4|2|4|4|1|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||2|2||||4|4||||Red|PERL 2014-2016|Volunteer: Moved|11||2|2|1|1|F|Black||13|No|Mother|28208|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||29|28277|Bachelors Degree|Single|Business: Clerical|28202|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500008321|503980164|31|0|2|504047655|31|0|2|500801295|2||-2||4|3|500014681||-2|500014681|-2|0|10|||17159|12|||1|828943|-1|4|3|44
503666549|BBBS of Greater Charlotte|Main Office|C|Active|2014-12-11|NaT|Baseline|2014-12-05|2014-12-11|Complete|Done|4|1|4|1|3|4|2.83|||||||||3|4|4|4|4|4|3.83|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016, Cabarrus County||27.1||1|1|1|1|M|Black||13|No|Mother|28025|One Parent: Female|$75,000 to $99,999||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|Black||35|28027|Bachelors Degree|Married|Finance|28217|1|9|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|277|60|598|500000170|500022817|503668509|31|0|1|504106972|31|0|1|500801599|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||46|2|||1|829407|-1|4|3|44
504139056|BBBS of Greater Charlotte|Main Office|C|Active|2014-12-09|NaT|Baseline|2014-12-05|2014-12-09|Complete|Done|4|4|4|4|4|4|4|||||||||2|4|4|2|4|4|3.33|||||||||4|4|4|4||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|||27.2||1|1|1|1|F|Black||13|No|Mother|28217|One Parent: Female|Unknown|Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||28|28105|Masters Degree|Married|Business: Mgt, Admin|28211|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|504094626|31|0|2|503991266|1|0|2|500801765|2||-2||2|1|||-2||-2|0|5|||17159|12|||1|829533|-1|4|3|44
503893808|BBBS of Greater Charlotte|Main Office|C|Completed|2014-12-20|2015-10-28|Baseline|2014-12-11|2014-12-20|Complete|Done|4|4|4|2|4|4|3.67|||||||||4|1|4|4|4|4|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Red||Volunteer: Moved|10.3||2|2|1|1|M|Black||13|No|GrandMother|28208|One Parent: Female|Unknown||No||School|General Community||Match Support|M|Asian||27|28203|Bachelors Degree|Single|Finance: Accountant|28202|1|10|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|277|60|598|500000170|500013745|503227914|31|0|1|503976460|4|0|1|500803592|2||-2||4|3|||-2|500014506|-2|0|4|||7462|13|||1|832093|-1|4|3|44
504083467|BBBS of Greater Charlotte|Main Office|C|Active|2014-12-22|NaT|Baseline|2014-12-19|2014-12-22|Complete|Done|4|4|4|4|4|3|3.83|||||||||2|4|3|3|3|3|3|||||||||4|4|4|4||||||3|2|3|3|2.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016||26.8||1|1|1|1|M|Black||11|No|Mother|28226|One Parent: Female|$30,000 to $34,999||No||School|General Community|PERL 2014-2016|Match Support|M|White||34|28214|Bachelors Degree||Transport: Flight Attendant|21804|7|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500018851|504085496|31|0|1|504003996|1|0|1|500805363|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||17159|12|||1|835500|-1|4|3|44
