InterviewNum|AgencyName|AgencyGroup|OfficeName|TeamName|Hybrid|MatchType|MatchStatus|QueueDescription|TimeInQueue|MatchSupportLevel|MatchReportSources|PendingMatchDate|MatchOpenDate|MatchCloseDate|MatchClosureReasons|MatchClosurePrimaryReason|MatchClosureSecondaryReason|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildGrade|ChildLivingSituation|ChildIncomeLevel|MilitaryParent|ParentDeployed|ChildFamilyAssistance|ChildFreeReducedlunch|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|Beg|Open|Close|End|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|ChildPartKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolPartKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|MatchKey|QueueKey|MatchTypeKey|MatchActivityKey|MatchSiteKey|StatusKey|MatchSupportLevelKey|ChildReportSourcesKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|MatchReportSourcesKey|CustodialAdultEmployerHash
21|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|733|Green||2015-02-24|2015-02-26|NaT||||24.1||1|1|1|1|M|Black||14|No|Mother|28278|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|Black||29|28209|Bachelors Degree|Single|Finance|20877|0|8|TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504160892|504162947|31|0|1|504171934|31|0|1|500815454|10|2|-2||2|1||-2||-2|0|4|||130|1|||1||2876415545463317777
27|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|715|Green||2015-03-08|2015-03-16|NaT||||23.5||1|1|1|1|M|Black||10|No|Mother|28211|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||31|28209|Bachelors Degree|Married|Medical|70112|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503314773|503314167|31|0|1|504176084|1|0|1|500817494|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||4253272603994307857
30|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|705|Yellow||2015-03-10|2015-03-26|NaT||||23.2||1|1|1|1|F|Black||11|No|Mother|28227|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||29|28226|Bachelors Degree|Single|Finance: Accountant|28202|0|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504194601|504184323|31|0|2|504032490|1|0|2|500817776|10|2|-2||2|2||-2||-2|0|4|||7464|9|||1||5822555200185981373
33|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|700|Green||2015-03-14|2015-03-31|NaT||||23||1|1|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Business: Sales|28277|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501843066|501843435|31|0|2|504152982|1|0|2|500818696|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||0
37|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|686|Green||2015-04-13|2015-04-14|NaT||||22.5||1|1|1|1|F|Black||13|No|Mother|28205|5|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|Black||27|28262|Some College|Single|Medical: Healthcare Worker|28210|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504242976|504245092|31|0|2|504198992|31|0|2|500823043|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||3988279022378749151
38|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|680|Green|Cabarrus County|2015-04-13|2015-04-20|NaT||||22.3||1|1|1|1|F|Black||7|No|Mother|28083||One Parent: Female|$25,000 to $29,999|||Y|No||Self|General Community|Cabarrus County|Match Support|F|White||54|28081|Some College|Married|Finance: Banking|28026|13|5|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504075474|502762654|31|0|2|503792949|1|0|2|500822904|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|4058276550489173605
42|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|670|Green|Cabarrus County|2015-04-16|2015-04-30|NaT||||22||1|1|1|1|F|Black||9|No|Mother|28083|1|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|F|Multi-race (Asian & White)||33|28025|Associate Degree|Married|Business: Marketing|28269|10|0|Self|Self|Big|General Community|Amachi, Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504241299|504243414|31|0|2|504194344|37|0|2|500823537|10|2|500016307||2|1|500016374|-2|500000294, 500016374|-2|34|2|||7464|9|||1|500016374|1579263579908564057
43|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|665|Green||2015-04-28|2015-05-05|NaT||||21.8||1|1|1|1|F|White||15|No|Mother|28227|8|One Parent: Female|$35,000 to $39,999||||Yes||School|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Law: Paralegal|28211|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504235352|504237484|1|0|2|504200139|1|0|2|500825073|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||8961132295198487522
44|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|665|Green||2015-04-22|2015-05-05|NaT||||21.8||1|1|1|1|M|White||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999||||Yes||School|General Community||Match Support|M|White||51|28173|Masters Degree|Married|Self-Employed, Entrepreneur|28173|19|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504235369|504237484|1|0|1|503937954|1|0|1|500824366|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||8961132295198487522
45|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|658|Green||2015-04-15|2015-05-12|NaT||||21.6||1|1|1|1|F|White||10|No|Mother|28277|4|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|F|White||29|29708|Bachelors Degree|Married|Medical|28105|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503889301|503891297|1|0|2|504021478|1|0|2|500823483|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||6156547733130613405
46|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|657|Green||2015-05-08|2015-05-13|NaT||||21.6||1|1|1|1|F|White||10|No|Mother|28214|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|F|White||28|28206|Bachelors Degree|Single|Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504231269|504233379|1|0|2|503927707|1|0|2|500826291|10|2|-2||2|1||-2||-2|0|3|||46|2|||1||0
49|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|651|Green|PERL 2014-2016|2015-04-29|2015-05-19|NaT||||21.4||1|1|1|1|F|White||10|No|GrandMother|28210|3|Other Relative|Unknown||||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||28|28205|Some College|Single|Transport: Driver|28277|8|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504234369|503470938|1|0|2|504116244|35|0|2|500825294|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||46|2|||1|500014681|7044657180546140448
50|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|648|Green||2015-05-22|2015-05-22|NaT||||21.3||1|1|2|2|F|Black||13|No|Mother|28212|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502930499|502931919|31|0|2|502564910|31|0|2|500828045|10|2|-2||2|1||-2||-2|0|10|||17161|11|||1||3402014428779854546
54|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|623|Green|PERL 2014-2016|2015-06-09|2015-06-16|NaT||||20.5||1|1|1|1|M|Black||15|No|GrandMother|28208|7|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|3|10|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|503944459|503946467|31|0|1|504260502|1|0|1|500829606|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||7462|13|||1|500014681|7044657180546140448
55|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|623|Green||2015-05-29|2015-06-16|NaT||||20.5||1|1|1|1|M|Black||13|No|Mother|28216|6|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|M|White||26|28202|Bachelors Degree|Single|Business|28217|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504247189|504249305|31|0|1|504228103|1|0|1|500828700|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||3402014428779854546
62|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|608|Green||2015-07-01|2015-07-01|NaT||||20||1|1|1|1|M|Black||9|No|Mother|28269|1|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|M|Black||28|28205|Bachelors Degree|Single|Finance|28202|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504219209|504221323|31|0|1|504301519|31|0|1|500831883|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||0
66|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|582|Green||2015-07-16|2015-07-27|NaT||||19.1||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|||Y|Yes||Relative|General Community||Match Support|F|White||29|28209|Bachelors Degree|Single|Retail: Mgt|28217|3|3|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504312629|504314787|31|0|2|504262612|1|0|2|500833665|10|2|-2||2|1||-2||-2|0|3|||17159|12|||1||237874676114443178
67|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|582|Green|PERL 2014-2016|2015-07-20|2015-07-27|NaT||||19.1||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Asian||28|28203|Bachelors Degree|Single|Consultant|28202|1|1|Current/Previous Big|Other Big|Big|General Community|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500008321|504312569|504314787|31|0|2|504208036|4|0|2|500833808|10|2|-2||2|1|500014681|-2|500014505, 500015184|-2|0|4|||17159|12|||1|500014681|237874676114443178
68|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|581|Green||2015-07-23|2015-07-28|NaT||||19.1||1|1|1|1|M|Black||10||GrandMother|28213|2|Grandparents|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||28|28204||Single|Finance: Accountant|28277|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503022461|501332937|31|0|1|504323998|1|0|1|500834322|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||0
70|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|565|Green||2015-08-13|2015-08-13|NaT||||18.6||1|1|1|1|F|Black||13|No|Mother|28214|6|One Parent: Female|$50,000 to $59,999||||Yes||Self|General Community||Match Support|F|White||29|28273|Masters Degree|Married|Finance: Accountant|28210|3|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504328960|504331182|31|0|2|504215323|1|0|2|500836079|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||8503368421346667831
71|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|565|Green||2015-07-23|2015-08-13|NaT||||18.6||1|1|1|1|F|Black||10|No|Mother|28216|2|One Parent: Female|$30,000 to $34,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||34|28031||Single|Self-Employed, Entrepreneur||9|8|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504186133|504188242|31|0|2|504122609|1|0|2|500834256|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1||8136849793711030748
72|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|564|Green||2015-07-22|2015-08-14|NaT||||18.5||1|1|1|1|M|Black||13|No|Mother|28273|6|One Parent: Female|$35,000 to $39,999||||No||Self|General Community||Match Support|M|Black||56|28273|Some College|Married|Govt|28228|0|7|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|504284556|504286757|31|0|1|504260574|31|0|1|500834204|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||2392572474128905139
75|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|547|Green|PERL 2014-2016, Cabarrus County|2015-08-14|2015-08-31|NaT||||18||1|1|1|1|F|Black||9|No|Mother|28075|1|Two Parent|$10,000 to $14,999||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||26|28027|Bachelors Degree|Single|Medical|28025|0|8|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504298787|504301001|31|0|2|504325174|31|0|2|500836212|10|2|500016307||2|1|500014681, 500016374|-2|500016374|-2|0|4|||46|2|||1|500014681, 500016374|7044657180546140448
79|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|532|Green||2015-09-01|2015-09-15|NaT||||17.5||1|1|1|1|M|Black||9|Yes|GrandMother|28269|1|Grandparents|Less than $10,000|||Y|Yes||School|General Community|Amachi|Match Support|M|White||32|28205|Bachelors Degree|Married|Real Estate: Realtor|28202|6|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504185266|503032503|31|0|1|504213307|1|0|1|500838024|10|2|-2||2|1|500000294|-2||-2|0|4|||17159|12|||1||7044657180546140448
80|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|531|Green|PERL 2014-2016|2015-09-10|2015-09-16|NaT||||17.4||1|1|1|1|M|Some Other Race||13|No|Mother|28217|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||38|28205|Masters Degree|Married|Human Services: Social Worker|28204|5|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504155180|501093096|41|0|1|502462446|1|0|1|500839295|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||7464|9|||1|500014681|358434295995756137
81|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|525|Green|PERL 2014-2016|2015-09-13|2015-09-22|NaT||||17.2||2|2|1|1|F|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Community|PERL 2014-2016|Match Support|F|White||26|28202|Bachelors Degree|Single|Finance: Banking|28262|1|7|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|504013056|504015071|31|0|2|504219921|1|0|2|500839610|10|2|-2||2|1|500014681|-2||-2|0|4|||17159|12|||1|500014681|0
82|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|524|Green|PERL 2014-2016|2015-09-10|2015-09-23|NaT||||17.2||2|2|1|1|M|Black||10|No|Mother|28214|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||25|28227|Bachelors Degree|Single|Insurance|28277|1|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503779386|503781363|31|0|1|504333970|31|0|1|500839160|10|2|-2||2|1|500014681|-2||-2|0|4|||7464|9|||1|500014681|1546374315672654438
83|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|519|Green||2015-08-22|2015-09-28|NaT||||17.1||3|3|1|1|F|Black||14|No|Mother|28216|7|Two Parent|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||43|28269|Masters Degree|Single|Business: Mgt, Admin||0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502186245|501610196|31|0|2|504248899|1|0|2|500836970|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||7044657180546140448
84|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|518|Green|PERL 2014-2016|2015-09-23|2015-09-29|NaT||||17||1|1|1|1|M|Black||11|No|Mother|28214|4|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28273|Bachelors Degree|Single|Insurance|28226|7|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|504153965|504156015|31|0|1|504372591|1|0|1|500841770|10|2|-2||2|1|500014681|-2||-2|0|4|||7464|9|||1|500014681|0
85|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|512|Green||2015-09-24|2015-10-05|NaT||||16.8||1|1|1|1|F|Black||12|No|Mother|28215|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Multi-Race (None of the above)||27|28269|Bachelors Degree|Single|Transport: Flight Attendant|28208|1|5|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504358312|504320644|31|0|2|504048355|7|0|2|500842174|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||2141487034287122220
86|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|512|Green||2015-09-28|2015-10-05|NaT||||16.8||1|1|1|1|M|Black||10|No|Mother|28213|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Consultant|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504179804|504181918|31|0|1|504337207|1|0|1|500842586|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||7044657180546140448
89|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|498|Green||2015-10-06|2015-10-19|NaT||||16.4||1|1|1|1|F|Black||8|No|Mother|28203|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||24|28202|Masters Degree|Single|Education: Teacher|28208|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504388144|504390375|31|0|2|504365599|1|0|2|500844802|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||2876415545463317777
93|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|487|Green||2015-10-08|2015-10-30|NaT||||16||1|1|1|1|F|Black||10|No|Mother|28216|4|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|F|Black||31|28216|Bachelors Degree|Single|Arts, Entertainment, Sports|28202|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504345626|504347850|31|0|2|504373316|31|0|2|500845709|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||1712849328738258411
94|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|487|Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2015-10-08|2015-10-30|NaT||||16|Y|1|1|1|1|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28204|Masters Degree|Married|Consultant||0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|504254978|504257111|3|0|1|504379733|1|0|1|500845639|10|2|-2||2|1|500014681|-2|500014681|-2|0|5|||46|2|||1|500011312, 500014681|0
96|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|481|Green||2015-10-20|2015-11-05|NaT||||15.8||1|1|1|1|M|Black||8|No|Mother|28269|K|One Parent: Female|$30,000 to $34,999||||Yes||School|General Community||Match Support|M|White||27|28204|Bachelors Degree|Married|Business: Mgt, Admin|28117|0|6|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504275417|504277617|31|0|1|504249590|1|0|1|500849815|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||4148565630505427365
97|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|475|Green||2015-10-21|2015-11-11|NaT||||15.6||1|1|1|1|M|Black||10|Yes|Mother|28216|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community|Amachi|Match Support|M|Black||41|28214|Some College|Married|Business|28287|0|3|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504207638|504209750|31|0|1|504357457|31|0|1|500850393|10|2|-2||2|1|500000294|-2||-2|0|4|||17159|12|||1||7674215580094440446
98|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|475|Green|PERL 2014-2016|2015-10-29|2015-11-11|NaT||||15.6||1|1|1|1|F|Black||10|No|Mother|28216|3|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Hispanic||26|28031|Bachelors Degree|Single|Tech: Research/Design|28117|0|8|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504390954|504393193|31|0|2|504231700|3|0|2|500853984|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1|500014681|3650724132819756420
99|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|474|Green|Cabarrus County|2015-11-10|2015-11-12|NaT||||15.6||1|1|1|1|M|Black||6|No|Mother|28081|K|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28025|Bachelors Degree|Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504366634|502790820|31|0|1|504346767|1|0|1|500858202|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||17159|12|||1|500016374|7044657180546140448
102|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|470|Green|PERL 2014-2016|2015-11-05|2015-11-16|NaT||||15.4||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28216|Bachelors Degree|Married|Business|28202|0|10|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504378557|1|0|1|500856483|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|500014681|3402014428779854546
104|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|469|Green|PERL 2014-2016, Cabarrus County|2015-11-10|2015-11-17|NaT||||15.4||1|1|1|1|M|White||15|Yes|Mother|28025|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28025|High School Graduate|Single|Business: Sales|28025|5|0|Local TV|Media|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|503821678|503823656|1|0|1|504468148|1|0|1|500858177|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7438|1|||1|500014681, 500016374|7044657180546140448
105|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|469|Green|PERL 2014-2016, Cabarrus County|2015-11-10|2015-11-17|NaT||||15.4||1|1|1|1|M|White||12|Yes|Mother|28025|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||32|28025|Bachelors Degree||Business: Sales||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|503821686|503823656|1|0|1|504460050|1|0|1|500858397|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7496|10|||1|500014681, 500016374|7044657180546140448
108|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|463|Green|PERL 2014-2016|2015-11-06|2015-11-23|NaT||||15.2||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28208|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||30|28204|Some College|Single|Medical|28208|3|3|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504278828|504281028|38|0|2|504354967|35|0|2|500857068|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500014681|2378213070582218846
109|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|462|Green||2015-11-13|2015-11-24|NaT||||15.2||1|1|1|1|M|Black||12|No|Mother|28211|5|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||48|28105||Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504227502|504229617|31|0|1|504460839|31|0|1|500859784|10|2|-2||2|1|500000294|-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1||2077565980961547475
110|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|456|Yellow|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2015-11-17|2015-11-30|NaT||||15||1|1|2|2|F|Hispanic||13|No|Mother|28205|6|Two Parent|Unknown||||Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504331538|504333760|3|0|2|503843020|3|0|2|500860738|10|2|-2||2|2|500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500011312, 500014681|0
114|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|442|Green|Amachi, PERL 2014-2016|2015-11-20|2015-12-14|NaT||||14.5||1|1|1|1|F|Black||15|Yes|Mother|28215|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi, PERL 2014-2016|Match Support|F|White||30|28203|Bachelors Degree|Single|Business|60611|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|503611732|503613600|31|0|2|504421910|1|0|2|500862006|10|2|-2||2|1|500000294, 500014681|-2|500014681|-2|0|10|||17159|12|||1|500000294, 500014681|0
115|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|441|Green|PERL 2014-2016|2015-11-30|2015-12-15|NaT||||14.5||1|1|1|1|F|Black||15|No|Mother|28215|9|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||26|28213|Bachelors Degree|Single|Business: Mgt, Admin|28105|2|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500021785|504393421|504395660|31|0|2|504395484|31|0|2|500863556|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||46|2|||1|500014681|5081726734274569781
120|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|411|Green|PERL 2014-2016|2016-01-04|2016-01-14|NaT||||13.5||1|1|1|1|F|Black||10|No|Mother|28203|3|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||25|28209|Bachelors Degree|Single|Business|28277|1|0|Bowl For Kids Sake|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504388295|504390534|31|0|2|504404378|1|0|2|500870013|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||132|8|||1|500014681|2141487034287122220
124|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|395|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-01-20|2016-01-30|NaT||||13||1|1|1|1|F|Black||7|No|Mother|28075|K|Two Parent|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||36|28036|Bachelors Degree|Married|Self-Employed, Entrepreneur|28036|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504453477|504455735|31|0|2|503803589|1|0|2|500873679|10|2|-2||2|1||-2||-2|0|5|||7464|9|||1|500007920, 500011315, 500011316|2141487034287122220
125|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|394|Green||2016-01-12|2016-01-31|NaT||||12.9||1|1|1|1|M|Black||8|Yes|Mother|28215|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|M|White||30|28205|Bachelors Degree||Arts, Entertainment, Sports|28206|0|3|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504231851|504233090|31|0|1|503291779|1|0|1|500871254|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||7327400833679234452
126|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|394|Green||2016-01-08|2016-01-31|NaT||||12.9||1|1|2|2|F|Black||8|Yes|Mother|28262|2|One Parent: Female|$25,000 to $29,999|||Y|Yes||Relative|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504538972|504402454|31|0|2|502171015|31|0|2|500870863|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|3|||7496|10|||1||6156547733130613405
127|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|393|Green|Cabarrus County|2016-01-25|2016-02-01|NaT||||12.9||1|1|1|1|F|Multi-race (Hispanic & White)||8|No|Mother|28025||One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|Multi-race (Black & White)||24|28027|Bachelors Degree|Single|Law: Police Officer|28078|1|3|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504533508|504535058|35|0|2|504443510|36|0|2|500875127|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|2141487034287122220
128|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|390|Green|Cabarrus County|2016-01-25|2016-02-04|NaT||||12.8||1|1|1|1|F|Multi-race (Black & White)||6|No|Mother|28025|K|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Cabarrus County|Match Support|F|White||36|28025|Some College|Divorced|Finance: Banking|28262|0|5|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504533461|504535058|36|0|2|504565015|1|0|2|500875147|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||17159|12|||1|500016374|2141487034287122220
130|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|382|Green|PERL 2014-2016|2016-01-29|2016-02-12|NaT||||12.6||1|1|1|1|M|Black||11|Yes|Mother|28215|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||29|28262|Some College|Single|Business|28204|0|4|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT, VOL - Thrive - Intro|Match Support|0|1|0|1|277|60|598|500000170|500020753|504230975|504233090|31|0|1|504284612|31|0|1|500876290|10|2|-2||2|1|500000294, 500014681|-2|500008492, 500011315, 500011316, 500014681|-2|0|4|||7462|13|||1|500014681|7327400833679234452
131|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|381|Green|Cabarrus County|2016-02-01|2016-02-13|NaT||||12.5||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28025|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||28|28027|Masters Degree|Single|Govt|28273|3|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504468562|504470835|36|0|1|504556956|31|0|1|500876668|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|500016374|7044657180546140448
135|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|372|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-09|2016-02-22|NaT||||12.2||1|1|1|1|F|Multi-race (Black & White)||10|Yes|Foster Parent|28216|4|One Parent: Female|$40,000 to $44,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||45|28208|Bachelors Degree|Single|Education: Teacher|28208|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504498650|504500981|36|0|2|504131389|31|0|2|500878445|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1|500007920, 500011315, 500011316|0
136|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|371|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-10|2016-02-23|NaT||||12.2||1|1|1|1|M|Black||11|No|Mother|28262|3|One Parent: Female|$30,000 to $34,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504295805|504298006|31|0|1|504337975|1|0|1|500878715|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1|500007920, 500011315, 500011316|5923747279518652886
138|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|367|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-22|2016-02-27|NaT||||12.1||1|1|1|1|F|Black||9|Yes|Mother|28208|2|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|F|Black||35|28216|Masters Degree|Married|Medical||0|3|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504404998|504403590|31|0|2|504481744|31|0|2|500880569|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|500007920, 500011315, 500011316|4309014537710246316
140|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|365|Yellow||2016-02-23|2016-02-29|NaT||||12||2|2|1|1|M|White||9|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||22|28215|Some College|Single|Finance|28215|0|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|503661137|503646117|1|0|1|504531427|1|0|1|500881061|10|2|-2||2|2||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||0
141|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|365|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-17|2016-02-29|NaT||||12||1|1|1|1|M|Black||9|No|Mother|28214|2|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|White||23|28202|Bachelors Degree|Single|Consultant|28202|0|5|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500021785|504153377|504155427|31|0|1|504487777|1|0|1|500879869|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|500007920, 500011315, 500011316|1335047838269305508
142|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|365|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-19|2016-02-29|NaT||||12||1|1|1|1|F|Black||7|No|Mother|28211|K|One Parent: Female|$25,000 to $29,999|Yes: Active|No|Y|Yes||Self|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Business|28270|10|8|AA Task Force|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504345301|504347523|31|0|2|504373845|1|0|2|500880266|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||6247|12|||1|500007920, 500011315, 500011316|1981915209225039472
143|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|358|Green|PERL 2014-2016, Cabarrus County|2016-02-29|2016-03-07|NaT||||11.8||1|1|1|1|M|Hispanic||8|No|Foster Parent|28078|1|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||50|28036||Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504433829|504436084|3|0|1|504470539|1|0|1|500882069|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|5|||46|2|||1|500014681, 500016374|7470110347975227693
144|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|355|Green|PERL 2014-2016|2016-02-26|2016-03-10|NaT||||11.7||1|1|1|1|M|Black||13|No|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28202|Bachelors Degree|Single|Law|28202|0|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504237243|504239358|31|0|1|504456306|1|0|1|500881682|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|500014681|7044657180546140448
145|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|355|Green||2016-03-04|2016-03-10|NaT||||11.7||1|1|1|1|M|Black||9|No|Mother|28213|3|One Parent: Female|$35,000 to $39,999||||Yes||School|General Community||Match Support|M|White||41|28078|Bachelors Degree|Married|Self-Employed, Entrepreneur|28031|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504262369|504264514|31|0|1|504538390|1|0|1|500883013|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||2806833304218536184
146|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|351|Green||2016-02-29|2016-03-14|NaT||||11.5||1|1|1|1|F|Black||13|No|Mother|28278|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||39|28134|Bachelors Degree|Single|Business: Marketing|28204|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504161470|504162947|31|0|2|504396335|1|0|2|500882097|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||2876415545463317777
148|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|342|Yellow|Cabarrus County|2016-03-09|2016-03-23|NaT||||11.2||1|1|1|1|M|Black||10|No|Mother|28027|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||35|28083|High School Graduate|Married|Medical||8|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504563369|504565703|31|0|1|504600175|1|0|1|500883737|10|2|500016307||2|2|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|500016374|6200244613298520712
150|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|336|Green|Amachi|2016-03-15|2016-03-29|NaT||||11||1|1|2|2|M|Black||7|Yes|Mother|28208|K|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|Black||35|28273|Some College|Married|Business: Marketing|28203|1|1|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504405002|504403590|31|0|1|504241664|31|0|1|500884837|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|500000294|4309014537710246316
151|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|329|Green||2016-03-01|2016-04-05|NaT||||10.8||1|1|1|1|M|Black||7|No|Mother|28273|K|One Parent: Female|$45,000 to $49,999|||Y|Yes||School|General Community||Match Support|M|White||25|28210|Bachelors Degree|Single|Finance|28211|10|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504276350|504278550|31|0|1|504273397|1|0|1|500882201|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||1176389127668227778
152|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|328|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-03-30|2016-04-06|NaT||||10.8||1|1|1|1|M|Black||12|No|Mother|28208|5|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Community||Match Support|M|White||32|28203|Juris Doctorate (JD)|Single|Law: Lawyer|28277|1|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|503952082|503954090|31|0|1|504546069|1|0|1|500887070|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|3|||46|2|||1|500007920, 500011315, 500011316|0
153|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|315|Green||2016-04-08|2016-04-19|NaT||||10.3||1|1|1|1|M|White||11|No|Mother|28277|4|One Parent: Female|$75,000 to $99,999||||No||School|General Community||Match Support|M|White||53|28270|Masters Degree|Married|Self-Employed, Entrepreneur||15|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504581060|504583394|1|0|1|504503934|1|0|1|500888341|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||5081726734274569781
154|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|315|Green||2016-03-14|2016-04-19|NaT||||10.3||1|1|1|1|F|Black||8|No|Mother|28217|1|One Parent: Female|$25,000 to $29,999|||Y|No||Self|General Community||Match Support|F|White||28|28210|Masters Degree|Single|Finance: Accountant|28210|0|3|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504532539|504534872|31|0|2|504467958|1|0|2|500884487|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||1136572582102976964
157|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|310|Green|Cabarrus County, mentor2.0 2016|2016-03-28|2016-04-24|NaT||||10.2||1|1|1|1|F|Black||13|No|Mother|28027|7|Two Parent|$60,000 to $74,999||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||30|28269|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|2|Recruitment Event|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504602680|504605091|31|0|2|504579649|1|0|2|500886605|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7462|13|||1|500016374, 500016394|993637920138474088
158|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|309|Green||2016-04-08|2016-04-25|NaT||||10.2||1|1|1|1|M|White||11|No|Mother|28277|5|One Parent: Female|$60,000 to $74,999||||No||School|General Community||Match Support|M|White||40|28173|Bachelors Degree|Married|Business: Mgt, Admin|33637|9|4|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504240231|504242346|1|0|1|504523981|1|0|1|500888425|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||7406803744350640674
159|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|308|Green|Cabarrus County|2016-04-05|2016-04-26|NaT||||10.1||1|1|1|1|M|Black||8|No|Mother|28027|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||Therapist/Counselor|General Community|Cabarrus County|Match Support|M|White||28|28083|Some College|Married|Business||10|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504612286|504614697|31|0|1|504634827|1|0|1|500887835|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|5|||7464|9|||1|500016374|3409063327463232933
160|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|306|Green|PERL 2014-2016, Cabarrus County|2016-04-07|2016-04-28|NaT||||10.1||1|1|1|1|M|White||10|No|GrandMother|28124|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||35|28027|Bachelors Degree|Single|Tech: Computer/Programmer|28202|2|6|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, mentor2.0, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504640447|504638197|1|0|1|504266263|1|0|1|500888255|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014505, 500016374|-2|0|4|||17159|12|||1|500014681, 500016374|0
164|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|304|Green|VOL - PreMatch, VOL - Mentoring Hispanic Youth, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-04-21|2016-04-30|NaT||||10||1|1|1|1|M|Hispanic||7|No|Mother|28205|K|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|Hispanic||37|28205|Bachelors Degree|Single|Tech: Engineer|28255|7|10|Community Engagement|Special Event|Big|General Community|VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504636958|504639369|3|0|1|504549037|3|0|1|500889969|10|2|-2||2|1||-2|500007920, 500011312, 500011315, 500011316|-2|0|4|||18809|8|||1|500007920, 500011312, 500011315, 500011316|0
165|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|294|Green|PERL 2014-2016|2016-05-02|2016-05-10|NaT||||9.7||1|1|3|3|M|Multi-race (Black & White)||12|Yes|Mother|28215|6|One Parent: Female|$35,000 to $39,999||||No||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||57|28269|Bachelors Degree|Married|Finance: Accountant|28202|34|2|Omega Psi Phi|Fraternity/Sorority|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|502183411|502183840|36|0|1|500189229|31|0|1|500891295|10|2|-2||2|1|500000294, 500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||8694|14|||1|500014681|4203557099934965158
167|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|285|Green||2016-05-03|2016-05-19|NaT||||9.4||1|1|1|1|F|Black||7|No|Mother|28212||One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|Black||25|28277|Bachelors Degree|Single|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504260164|504262304|31|0|2|504523141|31|0|2|500891594|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||4802885652788112046
169|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|280|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-04-19|2016-05-24|NaT||||9.2||1|1|1|1|F|Black||10|No|Mother|28208|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||29|28210|Bachelors Degree|Single|Business: Sales|28269|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504556546|504558880|31|0|2|504283498|1|0|2|500889681|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1|500007920, 500011315, 500011316|6084148439133243542
170|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|279|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-11|2016-05-25|NaT||||9.2||2|2|1|1|M|Black||13||GrandMother|28213|3|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||25|28205|Bachelors Degree|Married|Real Estate: Realtor|28202|0|2|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|501332660|501332937|31|0|1|504556335|1|0|1|500892769|10|2|-2||2|1|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||17159|12|||1|500007920, 500011315, 500011316|0
171|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|273|Green||2016-05-16|2016-05-31|NaT||||9||1|1|1|1|F|Black||15|No|Mother|28212|8|One Parent: Female|$40,000 to $44,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||48|28212|Associate Degree|Single|Finance||11|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504473782|504476056|31|0|2|504550297|1|0|2|500893115|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1||2806833304218536184
172|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|273|Green||2016-05-13|2016-05-31|NaT||||9||1|1|1|1|M|Black||13|No|Mother|28227|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|Black||27|28205|Some College|Single|Retail: Sales|28210|2|6|Local Radio|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504425160|504427415|31|0|1|504509415|31|0|1|500893007|10|2|-2||2|1||-2||-2|0|4|||7437|1|||1||5544164653861671456
173|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|273|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-23|2016-05-31|NaT||||9||1|1|1|1|M|Black||8|No|Mother|28213|1|One Parent: Female|$40,000 to $44,999||||No||School|General Community||Match Support|M|White||27|28203|Bachelors Degree||Transport: Driver|28105|2|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504155409|504157461|31|0|1|504606544|1|0|1|500894080|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|500007920, 500011315, 500011316|5439372922340750169
174|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|263|Green|Cabarrus County|2016-05-24|2016-06-10|NaT||||8.6||4|4|1|1|F|Black||12|No|Mother|28081|5|One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|Black||25|28025|Bachelors Degree|Single|Insurance|28213|1|10|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|502789637|502790820|31|0|2|504703410|31|0|2|500894186|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|7044657180546140448
176|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|263|Green||2016-05-10|2016-06-10|NaT||||8.6||1|1|1|1|F|Black||9|No|Mother|28206|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||28|28203|Bachelors Degree|Living w/ Significant Other|Finance|28202|0|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504473041|504475315|31|0|2|504582115|1|0|2|500892533|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1||5228205320249384837
177|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|259|Green|Cabarrus County|2016-06-14|2016-06-14|NaT||||8.5||1|1|1|1|F|White||11|No|GrandMother|28124|5|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community|Cabarrus County|Match Support|F|White||45|28025|Some College||Business|28262|1|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504635786|504638197|1|0|2|504662207|1|0|2|500896660|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|0
178|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|257|Green|PERL 2014-2016|2016-05-27|2016-06-16|NaT||||8.4||1|1|1|1|F|Multi-Race (None of the above)||13|No|Mother|28215|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Black||26|28262|Bachelors Degree|Single|Journalist/Media|28206|2|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504507791|504510086|7|0|2|504650231|31|0|2|500895078|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500014681|7044657180546140448
179|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|257|Green||2016-05-24|2016-06-16|NaT||||8.4||1|1|1|1|F|Black||11|No|Mother|28216|4|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||27|28209|Bachelors Degree|Single|Medical|28054|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504628520|504630931|31|0|2|504409458|1|0|2|500894207|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||7044657180546140448
180|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|253|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-23|2016-06-20|NaT||||8.3||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28213|7|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|Asian||25|28204|Bachelors Degree|Single|Finance|28215|0|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504691840|504694268|36|0|1|504535890|4|0|1|500894068|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1|500007920, 500011315, 500011316|8773162532572605235
181|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|250|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-06-16|2016-06-23|NaT||||8.2||1|1|1|1|F|Black||9|No|Mother|28215|3|One Parent: Female|$75,000 to $99,999||||Yes||School|General Community||Match Support|F|White||35|28215|Associate Degree|Divorced|Business|28215|0|8|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504507824|504510119|31|0|2|504575855|1|0|2|500896954|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|500007920, 500011315, 500011316|4318803846885526429
182|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|245|Green||2016-06-10|2016-06-28|NaT||||8||1|1|1|1|M|Black||9|No|Mother|28203|3|Two Parent|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||26|28202|Masters Degree|Single|Finance: Economist||0|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504601244|504603655|31|0|1|504577016|1|0|1|500896409|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|5|||7464|9|||1||904091744937704216
183|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|243|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-06-16|2016-06-30|NaT||||8||1|1|1|1|F|Black||12|No|Mother|28211|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||27|28205|Some College||Medical|28269|0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504471617|504473895|31|0|2|504458762|31|0|2|500897003|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1|500007920, 500011315, 500011316|1545381051186164660
184|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|243|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-06-16|2016-06-30|NaT||||8||2|2|1|1|F|Black||12|No|Mother|28214|5|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||26|28203|Bachelors Degree|Married|Business: Mgt, Admin|29707|0|4|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|503976557|503978568|31|0|2|504538747|1|0|2|500896984|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||18809|8|||1|500007920, 500011315, 500011316|3198188609986797983
259|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|98|Green||2016-10-21|2016-11-22|NaT||||3.2||2|2|1|1|F|Black||10|No|Mother|28215|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||27|28204|Masters Degree||Business: Human Resources|28202|0|3|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|503602769|503604646|31|0|2|504787610|31|0|2|500918350|10|2|-2||2|1|500007920, 500011315, 500011316, 500014681|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||1786514887916898235
260|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|92|Green||2016-11-11|2016-11-28|NaT||||3||1|1|1|1|M|White||13|No|Mother|28277|8|One Parent: Female|$60,000 to $74,999||||No||Self|General Community|PERL 2014-2016|Match Support|M|White||26|28207|Masters Degree|Living w/ Significant Other|Tech: Engineer|28203|1|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504808434|504810913|1|0|1|504557160|1|0|1|500926948|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||5571803589598086587
261|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|91|Green||2016-11-08|2016-11-29|NaT||||3||1|1|1|1|F|Black||15|No|Mother|28211|9|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||47|28215|Masters Degree|Married|Education|28202|5|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504471621|504473895|31|0|2|504580592|31|0|2|500925801|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||1545381051186164660
262|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|91|Green||2016-10-24|2016-11-29|NaT||||3||1|1|1|1|F|Black||11|No|Mother|28209|5|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||23|28203|Bachelors Degree||Finance: Accountant|28031|0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504662612|504665039|31|0|2|504595097|1|0|2|500918825|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||2719955880210213907
263|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|90|Green||2016-11-09|2016-11-30|NaT||||3||1|1|1|1|F|White||12|Yes|Non-Relative: Other|28205|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||28|28202|Bachelors Degree|Single|Finance|28202|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504539986|504538455|1|0|2|504793129|1|0|2|500926111|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||2082620892288628337
264|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|86|Green|Cabarrus County|2016-11-22|2016-12-04|NaT||||2.8||1|1|1|1|F|Black||12|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||24|28262|Masters Degree|Single|Human Services: Social Worker|28027|0|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504937152|504939686|31|0|2|504797758|31|0|2|500930335|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|0
267|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|84|Green||2016-11-11|2016-12-06|NaT||||2.8||1|1|1|1|M|Black||12|No|Mother|28213|5|One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||33|28203|Bachelors Degree|Married|Business|32207|9|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|502383218|502383656|31|0|1|504867282|1|0|1|500926962|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|6854|8|||46|2|||1||20998188998147742
268|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|78|Green|Cabarrus County|2016-11-22|2016-12-12|NaT||||2.6||1|1|1|1|F|Black||8|No|Mother|28027|3|One Parent: Female|$15,000 to $19,999||||Yes||School|General Community|Cabarrus County|Match Support|F|White||51|28027|Masters Degree|Married|Business|28213|1|10|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504937124|504939686|31|0|2|504828127|1|0|2|500930334|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||17159|12|||1|500016374|0
271|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|69|Green||2016-12-05|2016-12-21|NaT||||2.3||1|1|1|1|M|Black||15|No|Mother|28227|8|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||25|28277|Bachelors Degree|Single|Business|28208|1|8|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504662357|504664784|31|0|1|504791469|31|0|1|500933117|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1||3557919386369667257
272|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|69|Green||2016-12-01|2016-12-21|NaT||||2.3||1|1|1|1|M|Black||12|No|Mother|28210|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|M|Black||30|28210|Bachelors Degree|Married|Military||1|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504565095|504567429|31|0|1|504860995|31|0|1|500932205|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||6156547733130613405
274|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|69|Green||2016-12-01|2016-12-21|NaT||||2.3||1|1|1|1|M|Black||7|No|Mother|28208|1|One Parent: Female|$40,000 to $44,999||||Yes||School|General Community||Match Support|M|White||25|28203|Bachelors Degree|Single|Medical|85286|1|1|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504532089|504534422|31|0|1|504631918|1|0|1|500932298|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||786532283575222488
