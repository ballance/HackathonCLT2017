MatchNum|AgencyName|AgencyGroup|OfficeName|TeamName|Hybrid|MatchType|MatchStatus|QueueDescription|TimeInQueue|MatchSupportLevel|MatchReportSources|PendingMatchDate|MatchOpenDate|MatchCloseDate|MatchClosureReasons|MatchClosurePrimaryReason|MatchClosureSecondaryReason|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildGrade|ChildLivingSituation|ChildIncomeLevel|MilitaryParent|ParentDeployed|ChildFamilyAssistance|ChildFreeReducedlunch|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|Beg|Open|Close|End|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|ChildPartKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolPartKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|MatchKey|QueueKey|MatchTypeKey|MatchActivityKey|MatchSiteKey|StatusKey|MatchSupportLevelKey|ChildReportSourcesKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|MatchReportSourcesKey|ChildSchoolHash|CustodialAdultEmployerHash
M2|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2938|Green||2007-11-13|2007-11-30|2015-12-16|Child: Graduated|Child: Graduated||96.5||1|1|2|2|F|Black||20|No|Relative: Other|28269||Grandparents|$20,000 to $24,999||||Yes||BBBS Board/Staff|General Community||Match Support|F|Black||35|28213|Masters Degree|Single|Business||4|0|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|1|0|1|0|277|60|598|500000170|500002335|501045214|501045484|31|0|2|500953330|31|0|2|500217682|10|2|-2||4|1||-2|500014505, 500016394|-1|0|13|||46|2|||1||0|0
M3|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|4094|Green||2006-01-03|2005-12-21|NaT||||134.5||1|1|1|1|M|White||20||Mother|28104|11|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||60|28270|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500261295|500261310|1|0|1|500188435|1|0|1|500073081|10|2|-2||3|1||-2||-2|0|10|||7464|9|||1||0|0
M4|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2567|Green||2009-09-04|2009-10-08|2016-10-18|Child: Graduated|Child: Graduated||84.3||3|3|1|1|F|Black||20|No|Mother|28226|11|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|F|White||33|28277|Bachelors Degree|Living w/ Significant Other|Unknown|28209|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|500826592|500826861|31|0|2|501314246|1|0|2|500382768|10|2|-2||4|1||-2||-2|0|5|||7464|9|||1||7501346876523517480|0
M5|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2924|Green|Amachi|2007-07-13|2007-07-20|2015-07-22|Child: Graduated|Child: Graduated||96.1||3|4|1|1|M|Black||20|Yes|Mother|28227|12|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|Amachi|Match Support|M|Black||57|28262||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500186682|500188056|31|0|1|500887363|31|0|1|500184396|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|0|0
M6|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2733|Green||2008-01-09|2008-01-28|2015-07-23|Child: Graduated|Child: Graduated||89.8||2|2|1|1|M|Black||20||Mother|28210|12|Other/Unknown|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28078|High School Graduate|Single|Finance: Accountant|28202|0|4|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500185601|500187235|31|0|1|501082220|1|0|1|500236473|10|2|-2||4|1||-2||-2|6854|8|||7458|9|||1||5493390640808358320|0
M7|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3128|Green||2007-02-13|2007-02-21|2015-09-15|Child: Graduated|Child: Graduated||102.8||1|1|3|3|M|Black||20|No|Mother|28083|12|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||52|28025||Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500012459|500546821|500547073|31|0|1|500790181|31|0|1|500159910|10|2|-2||4|1||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1||0|0
M8|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|833|Green||2013-04-11|2013-04-11|2015-07-23|Child: Graduated|Child: Graduated||27.4||4|4|2|2|F|Black||20|No|GrandMother|28269|12|One Parent: Female|$35,000 to $39,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|500874765|501755813|31|0|2|502038804|31|0|2|500692473|10|2|-2||4|1||-2||-2|34|2|||7496|10|||1||4565518866290635873|0
M9|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1861|Green||2010-06-07|2010-06-18|2015-07-23|Child: Graduated|Child: Graduated||61.1||1|1|2|2|F|Black||20|No|Mother|28217|12|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|502142541|502142970|31|0|2|501905673|31|0|2|500455759|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1||253338316288302752|0
M10|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3282|Red||2006-08-16|2006-08-23|2015-08-18|Child: Graduated|Child: Graduated||107.8||1|1|1|1|M|Black||20||Mother|28214||One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||38|28209|Bachelors Degree|Single|Construction|28247|0|2|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500474486|500474735|31|0|1|500491064|31|0|1|500118168|10|2|-2||4|3||-2||-2|34|2|||7447|3|||1||0|0
M11|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3908|Green|Amachi|2004-06-21|2004-06-21|2015-03-04|Child: Graduated|Child: Graduated||128.4||1|1|1|1|M|Black||20||Mother|28213|12|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||54|28203|Bachelors Degree|Married|Law: Lawyer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500186956|500188141|31|0|1|500189727|1|0|1|500037841|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|0|0
M12|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2856|Green||2007-10-11|2007-10-18|2015-08-13|Child: Graduated|Child: Graduated||93.8||2|2|1|1|F|Black||20||Mother|28217|11|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||35|28211|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|500186106|500187698|31|0|2|500778380|1|0|2|500202993|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||1010189231295710785|0
M13|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4411|Green||2003-07-23|2003-07-23|2015-08-20|Child: Graduated|Child: Graduated||144.9||1|1|1|1|M|Black||20||Mother|28216|11|One Parent: Female|Unknown||||No|Brochure|Media|General Community||Match Support|M|White||45|28226|Bachelors Degree|Married|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|500186435|500187988|31|0|1|500189358|1|0|1|500037395|10|2|-2||4|1||-2||-2|51|1|||7496|10|||1||253338316288302752|0
M14|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1410|Green||2011-08-08|2011-09-02|2015-07-13|Child: Graduated|Child: Graduated||46.3||1|1|1|1|M|Black||20|No|Mother|28212|11|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||31|28203|Masters Degree|Single|Finance: Banking||0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502436202|502436645|31|0|1|502642999|1|0|1|500549046|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1||1010189231295710785|6156547733130613405
M15|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3125|Green||2006-07-06|2006-08-01|2015-02-20|Child: Graduated|Child: Graduated||102.7||1|1|1|1|M|White||20||Mother|28226|11|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||39|28211|Masters Degree|Married|Law: Lawyer|28204|2|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|500395038|500395288|1|0|1|500392006|1|0|1|500104016|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1||7501346876523517480|0
M16|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2495|Yellow||2008-12-03|2008-12-12|2015-10-12|Child: Graduated|Child: Graduated||82||1|1|1|1|M|Black||20|No|Mother|28217|5|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28226|Bachelors Degree|Married|Tech: Engineer|28202|2|8|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|501347056|501347335|31|0|1|501217000|1|0|1|500322327|10|2|-2||4|2||-2||-2|34|2|||7446|3|||1||0|0
M17|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1949|Yellow||2010-05-28|2010-06-08|2015-10-09|Child: Graduated|Child: Graduated||64||1|1|2|2|F|Black||19|No|Mother|28269|7|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500017777|502045254|502045664|31|0|2|502171015|31|0|2|500454926|10|2|-2||4|2||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1||0|0
M18|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1807|Green|2010-2012 OJJDP JJI|2011-08-18|2011-08-31|2016-08-11|Child: Graduated|Child: Graduated||59.4||1|1|1|1|F|Black||19||Mother|28216|11|Two Parent|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||51|28277|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|502601023|502601540|31|0|2|502546883|1|0|2|500550809|10|2|-2||4|1|500005291|-2||-2|6854|8|||7464|9|||1|500005291|2374609189072499123|3351268171347533976
M19|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1247|Green||2012-02-06|2012-02-21|2015-07-22|Child: Graduated|Child: Graduated||41||1|1|1|1|F|Black||19|No|Mother|28226|11|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community||Match Support|F|White||34|28226|Bachelors Degree|Married|Unknown|29715|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502824908|502826191|31|0|2|502891382|1|0|2|500596373|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||5493390640808358320|0
M20|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3034|Red|Amachi|2006-10-29|2006-10-29|2015-02-18|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||99.7||2|3|1|1|F|Black||19|Yes|Mother|28262|10|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||48|28212||Single|Medical: Healthcare Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500185907|500187470|31|0|2|500697782|31|0|2|500134557|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|702163000107564368|0
M21|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1159|Green||2012-02-23|2012-03-08|2015-05-11|Child: Graduated|Child: Graduated||38.1||1|1|1|1|F|Black||19|No|Mother|28213|11|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||32|28262|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502893765|502895172|31|0|2|502874079|31|0|2|500599963|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||253338316288302752|0
M22|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1291|Green||2012-03-27|2012-03-30|2015-10-12|Child: Graduated|Child: Graduated||42.4||1|1|1|1|M|Black||19|No|GrandMother|28208|8|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community||Match Support|M|White||59|28277|Masters Degree|Single|Tech: Computer/Programmer|28203|3|4|Local Print|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502431164|502431607|31|0|1|502850528|1|0|1|500606503|10|2|-2||4|1||-2||-2|0|5|||7439|1|||1||0|0
M23|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3172|Green|Amachi|2006-05-25|2006-05-25|2015-01-30|Child: Graduated|Child: Graduated||104.2||1|1|4|4|F|Black||19|Yes|Mother|28083||One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500008321|500408135|500408385|31|0|2|500189709|31|0|2|500099932|10|2|500003586||4|1|500000294|-2|500000294, 500016374|-2|6854|8|||2230|7|||1|500000294|0|0
M24|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4066|Yellow||2004-10-29|2004-10-29|2015-12-17|Child: Graduated|Child: Graduated||133.6||3|3|1|1|M|Black||19|No|Mother|28025||One Parent: Female|Unknown||||No||Self|General Site||Match Support|M|Black||42|28025|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500186260|500187857|31|0|1|500189139|31|0|1|500037139|10|2|-2||4|2||-1||-2|0|10|||7464|9|||1||0|0
M25|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2402|Green||2009-01-13|2009-01-28|2015-08-27|Child: Graduated|Child: Graduated||78.9||1|1|1|1|F|Black||19|No|Mother|28027|6|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||39|28212|Bachelors Degree|Single|Medical: Healthcare Worker|28210|1|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|501516900|501517192|31|0|2|501438601|31|0|2|500332399|10|2|-2||4|1||-2||-2|6854|8|||7462|13|||1||0|2968153613205640519
M26|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1048|Yellow||2012-04-12|2012-05-04|2015-03-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.4||1|1|1|1|F|Black||19|No|Mother|28216|11|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|F|Black||48|28217|Bachelors Degree|Divorced|Medical: Admin|28232|11|5|Local TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502966254|500784955|31|0|2|502895517|31|0|2|500609631|10|2|-2||4|2||-2||-2|0|10|||7438|1|||1||3292090474897428830|1786514887916898235
M27|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1337|Green||2011-11-11|2011-12-08|2015-08-06|Child: Graduated|Child: Graduated||43.9||1|1|1|1|M|Black||19|No|Mother|28206|9|One Parent: Female|Less than $10,000|||Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||33|28213|Associate Degree|Single|Transport: Driver|28205|5|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500017732|502714405|502715293|31|0|1|502764673|31|0|1|500577475|10|2|-2||4|1|500005291|-2||-2|56|1|||7446|3|||1||1766165378108010922|0
M28|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2665|Red||2008-04-16|2008-05-01|2015-08-18|Child: Graduated|Child: Graduated||87.6||1|1|1|1|M|Black||19||Mother|28226||One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|White||37|28210|Some College|Single|Business: Mgt, Admin||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501092911|501064244|31|0|1|501176101|1|0|1|500261235|10|2|-2||4|3||-2||-2|0|4|||46|2|||1||0|0
M29|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3433|Red||2007-03-15|2007-03-27|2016-08-19|Child: Graduated|Child: Graduated||112.8||1|1|1|1|M|White||19|No|Mother|28081|9|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||46|28202||Single|Business: Sales||0|4|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500020753|500799303|500799571|1|0|1|500798390|1|0|1|500167062|10|2|-2||4|3|500016374|-2|500016374|-2|34|2|||7464|9|||1||0|0
M30|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3919|Red|Amachi|2005-02-10|2005-02-10|2015-11-04|Child: Graduated|Child: Graduated||128.8||1|1|1|1|F|Black||19|Yes|Mother|28205|12|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Match Support|F|Black||50|28215|Some College|Single|Finance: Banking||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500186905|500188151|31|0|2|500189677|31|0|2|500037790|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||7453|7|||1|500000294|0|0
M31|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2461|Yellow|Amachi|2008-08-11|2008-08-14|2015-05-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||80.9||1|1|4|4|F|Black||19|Yes|GrandMother|28273|10|Grandparents|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501300101|501300379|31|0|2|500346193|31|0|2|500281421|10|2|500003586||4|2|500000294|-2||-2|7294|13|||46|2|||1|500000294|0|0
M32|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2989|Red|Amachi|2006-12-26|2006-12-26|2015-03-03|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||98.2||1|1|1|1|F|Black||19|Yes|GrandMother|28217|12|Grandparents|Less than $10,000|||Y|No|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||34|28210|Bachelors Degree|Married|Finance: Accountant|28202|0|2|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500733695|500733962|31|0|2|500307108|1|0|2|500150172|10|2|500003586||4|3|500000294|-2||-2|7294|13|||2238|7|||1|500000294|253338316288302752|0
M33|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2484|Red||2008-08-27|2008-09-05|2015-06-25|Child: Graduated|Child: Graduated||81.6||2|2|1|1|M|Black||19||Mother|28214||One Parent: Female|Unknown||||No|AARTF|Neighbor/Friend|General Community||Match Support|M|Black||36|28214|Bachelors Degree|Single|Tech: Computer/Programmer|28147|0|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500185723|500187335|31|0|1|501310677|31|0|1|500284133|10|2|-2||4|3||-2||-2|6855|8|||7464|9|||1||0|0
M34|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2807|Green||2007-11-26|2007-11-26|2015-08-03|Child/Family: Moved|Child/Family: Moved||92.2||1|1|1|1|M|Black||19|No|Mother|28205|4|One Parent: Female|$15,000 to $19,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28226|Masters Degree|Single|Finance: Accountant||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|501060196|501060469|31|0|1|501036081|1|0|1|500223215|10|2|-2||4|1||-2||-2|34|2|||46|2|||1||0|0
M35|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2557|Green||2008-03-11|2008-04-29|2015-04-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||84||1|1|1|1|M|Black||19|No|Aunt|28269||One Parent: Female|$10,000 to $14,999|||Y|No||Therapist/Counselor|General Community||Match Support|M|Black||35|28213|Bachelors Degree|Single|Business: Sales||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500968246|500968516|31|0|1|501179573|31|0|1|500251681|10|2|-2||4|1||-2||-2|0|5|||46|2|||1||0|0
M36|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3360|Red||2006-04-25|2006-05-02|2015-07-14|Child: Graduated|Child: Graduated||110.4||1|1|1|1|M|Black||19||Mother|28215||Other/Unknown|Unknown||||No|Other|Faith Organization|General Community||Match Support|M|Black||49|28213|Bachelors Degree|Married|Finance: Banking|28288|4|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500185571|500187198|31|0|1|500188438|31|0|1|500089543|10|2|-2||4|3||-2||-2|5635|9|||7464|9|||1||0|0
M37|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2044|Green||2009-07-14|2009-08-07|2015-03-13|Volunteer: Moved|Volunteer: Moved||67.2||1|1|2|2|F|Black||19|No|Mother|28269|11|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||31|28269|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500011349|501641337|501641648|31|0|2|500835981|31|0|2|500373972|10|2|-2||4|1|500000294|-2|500000294|-2|0|10|||46|2|||1||4565518866290635873|7124320636013019662
M38|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2644|Green||2009-03-23|2009-03-28|2016-06-23|Child: Graduated|Child: Graduated||86.9||1|1|1|1|M|Black||19|No|Mother|28105|10|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||55|28173|||Unknown|28203|0|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|501506214|501506506|31|0|1|501588885|31|0|1|500351462|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||8735132144641863371|710802550313155478
M39|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2586|Red||2009-07-21|2009-07-21|2016-08-19|Child: Graduated|Child: Graduated||85||1|1|2|2|M|Hispanic||19|No|Mother|28025|12|One Parent: Female|Unknown||||Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500020753|501645192|501645515|3|0|1|501519306|1|0|1|500374818|10|2|-2||4|3|500016374|-2|500016374|-2|0|10|||7464|9|||1||6236652402957148873|0
M40|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2028|Green|2010-2012 OJJDP JJI|2011-08-10|2011-08-18|NaT||||66.6||1|1|1|1|M|Black||19|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Juris Doctorate (JD)|Single|Student: College|28208|0|0||Law Student Association|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|502205848|502206277|31|0|1|502624702|1|0|1|500549350|10|2|-2||2|1|500005291|-2||-2|0|10|||0|15|||1|500005291|702163000107564368|0
M41|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1947|Green|2010-2012 OJJDP JJI|2011-03-09|2011-03-31|2016-07-29|Child/Family: Moved|Child/Family: Moved||64||2|2|2|2|F|Black||19|No|Mother|28211|11|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28211||Married|Finance: Banking|28255|0|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501868921|501869291|31|0|2|501382633|1|0|2|500524206|10|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|500005291|7501346876523517480|0
M42|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1890|Green|Project Big, 2010-2012 OJJDP JJI|2011-05-09|2011-05-12|2016-07-14|Child: Graduated|Child: Graduated||62.1||1|1|3|4|F|Black||19||Mother|28208|7|Two Parent|$15,000 to $19,999||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||48|28214|Bachelors Degree|Single|Tech: Management|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Project Big|Enrollment|1|0|1|0|277|60|598|500000170|500017732|502537477|502537922|31|0|2|500189507|31|0|2|500535475|10|2|-2||4|1|500004640, 500005291|-2|500000294, 500004640|-2|0|4|||2238|7|||1|500004640, 500005291|0|0
M43|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|140|Green||2014-10-14|2014-10-16|2015-03-05|Child/Family: Moved|Child/Family: Moved||4.6||2|2|2|3|M|Black||19|No|GrandMother|28208|9|Grandparents|Unknown|||Y|Yes||School|General Site|mentor2.0 2014|Match Support|M|White||33|28202|Bachelors Degree|Married|Finance|28202|0|2|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|503236068|503237859|31|0|1|503976384|1|0|1|500783505|10|1|500014504||4|1|500014506|-1|500014505, 500014506|-2|0|4|||7462|13|||1||702163000107564368|0
M44|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1947|Green|Project Big, 2010-2012 OJJDP JJI|2011-03-30|2011-03-31|2016-07-29|Child: Graduated|Child: Graduated||64||2|2|1|1|M|Black||19|No|Mother|28216|11|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||38|28277|Bachelors Degree|Single|Arts, Entertainment, Sports|28203|3|6|UnitedMethodistChrch|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501631547|501631870|31|0|1|502170945|1|0|1|500528464|10|2|500004641||4|1|500004640, 500005291|-2||-2|0|10|||8529|7|||1|500004640, 500005291|253338316288302752|0
M45|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3066|Green|Amachi|2007-10-01|2007-10-01|2016-02-22|Child: Graduated|Child: Graduated||100.7||1|1|1|1|M|Black||19|Yes|Aunt|28208|11|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Match Support|M|White||46|28209|Masters Degree|Single|Self-Employed, Entrepreneur|28209|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500871683|500871952|31|0|1|500933829|1|0|1|500199601|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|2374609189072499123|0
M46|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1976|Red|2010-2012 OJJDP JJI, Cabarrus County|2011-03-11|2011-03-23|2016-08-19|Child: Graduated|Child: Graduated||64.9||2|2|1|1|F|Black||19|No|Mother|28027|9|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||43|28075|Bachelors Degree|Married|Business: Mgt, Admin||7|0|Recruitment Event|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500020753|501811385|501811730|31|0|2|502460013|31|0|2|500524684|10|2|-2||4|3|500016374|-2|500016374|-2|6854|8|||7459|10|||1|500005291, 500016374|5826822768343582573|0
M47|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2031|Green|Amachi|2010-12-02|2010-12-08|2016-06-30|Child: Graduated|Child: Graduated||66.7||4|4|1|1|M|Black||19|Yes|Mother|28227|11|One Parent: Female|Unknown|||Y|No||School|General Community|Amachi|Match Support|M|Black||52|28227|Masters Degree|Married|Education: Teacher|28227|2|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi, Project Big|Match Support|1|0|1|0|277|60|598|500000170|500013781|500186742|500188056|31|0|1|502397541|31|0|1|500501282|10|2|500003586||4|1|500000294|-2|500000294, 500004640|-2|0|4|||12183|14|635|1|1|500000294|1766165378108010922|0
M48|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3029|Green||2008-02-28|2008-02-29|2016-06-15|Child: Graduated|Child: Graduated||99.5||1|1|1|1|M|Multi-race (Black & White)||19|No|Mother|28227|10|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Consultant|28226|0|8|Other|Service Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|501185594|501185866|36|0|1|501153366|1|0|1|500248756|10|2|-2||4|1||-2||-2|0|4|||7452|6|||1||0|0
M49|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4275|Green||2004-10-14|2004-10-14|2016-06-28|Child: Graduated|Child: Graduated||140.5||1|1|1|1|M|White||18||Mother|28273||One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||51|28262|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500186133|500187724|1|0|1|500188930|1|0|1|500036930|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||0|0
M50|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2442|Green||2010-06-22|2010-06-30|NaT||||80.2||2|2|1|1|F|Black||18|No|Mother|28205|9|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||33|28203|High School Graduate|Single|Retail: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|501626226|501622822|31|0|2|502036832|1|0|2|500457771|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||0|0
M51|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3083|Green||2008-01-14|2008-02-19|2016-07-29|Child: Graduated|Child: Graduated||101.3||1|1|1|1|M|Black||18|No|Mother|28204|10|Two Parent|$40,000 to $44,999||||Yes||Self|General Community||Match Support|M|White||33|28202|Bachelors Degree|Married|Business: Marketing||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500997880|500998153|31|0|1|500990660|1|0|1|500237316|10|2|-2||4|1||-2||-2|0|10|||46|2|||1||7501346876523517480|6334475452707074991
M52|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1743|Red|2010-2012 OJJDP JJI|2011-07-19|2011-07-22|2016-04-29|Child: Graduated|Child: Graduated||57.3||1|1|1|1|M|Black||18|No|Mother|28208|7|One Parent: Female|$10,000 to $14,999||||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||46|28278|Bachelors Degree|Separated|Transport: Pilot|28208|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502588461|502588977|31|0|1|502636478|31|0|1|500546741|10|2|-2||4|3|500005291|-2||-2|6854|8|||46|2|||1|500005291|6745751685887553036|0
M53|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1085|Green||2013-05-10|2013-05-10|2016-04-29|Volunteer: Moved|Volunteer: Moved||35.6||1|1|1|1|F|Black||18|No|Mother|28216|9|Two Parent|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||33|28269|Bachelors Degree|Single|Human Services: Non-Profit|28202|0|8|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|503469094|503470960|31|0|2|501717376|1|0|2|500696470|10|2|-2||4|1||-2|500000294|-2|6854|8|||7464|9|||1||2374609189072499123|0
M54|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2764|Red||2009-01-12|2009-01-31|2016-08-26|Child: Graduated|Child: Graduated||90.8||1|1|1|1|F|Hispanic||18|No|Mother|28212|4|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community||Match Support|F|Hispanic||65|28269|Masters Degree|Single|Medical: Admin|28262|8|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500017777|501201377|501201651|3|0|2|501497622|3|0|2|500331903|10|2|-2||4|3||-2||-2|7016|11|||7446|3|||1||0|0
M55|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4389|Green||2004-06-17|2004-06-17|2016-06-23|Child: Graduated|Child: Graduated||144.2||1|1|1|1|M|Black||18||Mother|28215|10|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||42|27514||Married|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|500185778|500187368|31|0|1|500188776|1|0|1|500036776|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||6875312010577189564|0
M56|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|913|Red||2012-06-22|2012-07-31|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||30||1|1|1|1|M|Black||18|No|Mother|28031|8|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|White||26|28031|High School Graduate|Single|Personal Trainer/Coach|28117|0|4|Relative|Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502863781|502865175|31|0|1|503002010|1|0|1|500621061|10|2|-2||4|3||-2||-2|0|10|||17161|11|||1||3974159976843499574|1286881276054717070
M57|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2189|Green||2009-06-15|2009-06-19|2015-06-17|Child/Family: Moved|Child/Family: Moved||71.9||1|1|1|1|M|Black||18|No|Mother|30058|10|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||34|28215||Married|Consultant|28285|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501402710|501402995|31|0|1|501728845|1|0|1|500368860|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||0|5987230989236352701
M58|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1503|Green||2012-11-15|2013-01-24|NaT||||49.4||1|1|1|1|F|Hispanic||18|No|Mother|28277|9|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||24|28104|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503052841|503027860|3|0|2|503122069|1|0|2|500660497|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||3966805366522644621|8598768071652363430
M59|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|880|Yellow||2013-01-24|2013-01-26|2015-06-25|Child: Lost interest|Child: Lost interest||28.9||1|1|1|1|M|Black||18|Yes|Mother|28226|9|One Parent: Female|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Asian||29|28277|Bachelors Degree|Single|Real Estate: Realtor|28277|2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503268324|503270085|31|0|1|503253968|4|0|1|500676990|10|2|-2||4|2|500000294|-2||-2|6854|8|||7464|9|||1||7501346876523517480|7044657180546140448
M60|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1647|Red||2010-11-10|2010-11-23|2015-05-28|Child/Family: Moved|Child/Family: Moved||54.1||1|1|1|1|M|Black||18|No|Mother|28210|7|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||40|28278|Bachelors Degree|Married|Tech: Computer/Programmer||3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502308593|502309025|31|0|1|502262702|31|0|1|500492994|10|2|-2||4|3||-2||-2|0|10|||12183|14|1209|1|1||0|0
M61|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1305|Green||2012-10-19|2012-10-29|2016-05-26|Child: Graduated|Child: Graduated||42.9||2|3|2|3|F|Black||18|Yes|Mother|28210|9|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community|Amachi|Match Support|F|White||40|28214|Bachelors Degree|Single|Human Services: Non-Profit||3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500185812|500187400|31|0|2|500188912|1|0|2|500648551|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1||7872663507285703533|2604443421896951982
M62|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2296|Green|Amachi|2010-03-01|2010-03-18|2016-06-30|Child: Graduated|Child: Graduated||75.4||2|2|1|1|F|Black||18|No|Mother|28217|12|One Parent: Female|$25,000 to $29,999|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||40|28203|Some College|Living w/ Significant Other|Finance: Banking|28281|1|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500948129|500948399|31|0|2|501891556|1|0|2|500438403|10|2|500003586||4|1|500000294|-2||-2|34|2|||7464|9|||1|500000294|7301546317881317703|0
M63|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1909|Green|2010-2012 OJJDP JJI|2011-04-28|2011-05-12|2016-08-02|Child: Graduated|Child: Graduated||62.7||2|2|1|1|F|Black||18|No|GrandMother|28208|9|Grandparents|Unknown||||Yes|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||68|28262|Bachelors Degree|Living w/ Significant Other|Business: Clerical||2|0|Relative|Relative|Big|General Community|Amachi, Project Big|Match Support|1|0|1|0|277|60|598|500000170|500017732|502185074|502185503|31|0|2|502490418|31|0|2|500533846|10|2|-2||4|1|500005291|-2|500000294, 500004640|-2|5635|9|||17161|11|||1|500005291|2374609189072499123|0
M64|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1348|Red||2013-05-29|2013-06-21|2017-02-28|Child/Family: Moved|Child/Family: Moved||44.3||1|1|1|1|F|Black||18|No|Mother|28262|9|Two Parent|$75,000 to $99,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||25|28269|Bachelors Degree|Single|Education: Teacher|28210|0|4|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008321|503216769|503218550|31|0|2|503344849|31|0|2|500698465|10|2|-2||4|3||-2||-2|34|2|||46|2|||1||7432163260389731024|9141786906325747498
M65|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1561|Green|2010-2012 OJJDP JJI|2011-06-01|2011-06-30|2015-10-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||51.3||1|1|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28215|11|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28078|Bachelors Degree|Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|502570396|502570850|38|0|2|502545897|31|0|2|500539251|10|2|-2||4|1|500005291|-2||-2|34|2|||46|2|||1|500005291|6875312010577189564|6250057851021950913
M66|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2257|Green||2010-06-23|2010-06-25|2016-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||74.2||1|1|1|1|F|Black||18|No|Mother|28269|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||33|28262|Bachelors Degree|Single|Medical: Nurse|28262|4|9|AA Task Force|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502045258|502045664|31|0|2|502190790|31|0|2|500457916|10|2|-2||4|1||-2||-2|0|10|||6247|12|||1||0|0
M67|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1765|Green|2010-2012 OJJDP JJI|2011-09-26|2011-10-31|2016-08-30|Child: Graduated|Child: Graduated||58||1|1|1|1|F|Black||18|No|Mother|28208|12|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28262|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|502510347|502510796|31|0|2|502677833|31|0|2|500557844|10|2|-2||4|1|500005291|-2||-2|0|5|||7464|9|||1|500005291|216500609169513656|0
M68|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2603|Green||2010-01-04|2010-01-20|NaT||||85.5||3|3|1|1|M|White||18|No|Mother|28031|10|One Parent: Male|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||60|28269|||Medical: Admin|28207|0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500796255|500796529|1|0|1|501846438|1|0|1|500424314|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1||3455806768141331471|0
M69|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2613|Red|Amachi|2008-11-18|2008-11-24|2016-01-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||85.8||3|3|1|1|M|Black||18|Yes|Mother|28215|10|One Parent: Female|Unknown||||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Tech: Computer/Programmer||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500252077|501750989|31|0|1|501365749|1|0|1|500317108|10|2|500003586||4|3|500000294|-2||-2|7295|11|||46|2|||1|500000294|1010189231295710785|0
M70|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1354|Green||2013-06-11|2013-06-22|NaT||||44.5||2|2|1|1|M|Black||18|No|Mother|28269|10|One Parent: Female|$40,000 to $44,999|||Y|Yes||Self|General Community||Match Support|M|White||57|28277|Some College|Married|Business: Sales||28|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502370669|502371107|31|0|1|503472866|1|0|1|500700192|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||7458247995093008174|0
M71|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1202|Green||2012-10-23|2012-11-17|2016-03-03|Volunteer: Moved|Volunteer: Moved||39.5||2|2|3|3|F|Black||18|Yes|Mother|28216|9|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||41|28269|||Business: Human Resources|28206|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|501237971|503287812|31|0|2|501598429|31|0|2|500649363|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1||7432163260389731024|0
M72|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|973|Green||2013-09-17|2013-10-16|2016-06-15|Child: Graduated|Child: Graduated||32||1|1|1|1|F|Black||18|No|GrandMother|28213|10|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|White||29|28211|Juris Doctorate (JD)|Married|Law|28202|0|9|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503425736|503427601|31|0|2|503519747|1|0|2|500711543|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||7432163260389731024|7044657180546140448
M73|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1254|Green||2013-09-12|2013-09-30|NaT||||41.2||2|2|1|1|F|Black||18|No|GrandMother|28214|9|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||26|28078|Masters Degree|Single|Education: Teacher|28212|0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502421176|502421614|31|0|2|503497451|31|0|2|500710577|10|2|-2||3|1||-2||-2|0|4|||7464|9|||1||702163000107564368|6054903719040220574
M74|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|495|Green|PERL 2014-2016, Cabarrus County|2015-10-06|2015-10-29|NaT||||16.3||4|4|1|1|F|White||18|No|Father|28025||One Parent: Male|Unknown||||No||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||68|28027|Associate Degree|Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|500341548|500341682|1|0|2|504323327|1|0|2|500844725|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|3|||17159|12|||1|500014681, 500016374|0|0
M75|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|349|Green||2014-10-07|2014-10-07|2015-09-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||11.5||1|1|2|2|F|Black||18|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||48|28079||Married|Finance|28255|4|2|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043491|504045509|31|0|2|503984584|31|0|2|500781133|10|1|500014504||4|1||-1|500014506|-1|0|4|||7462|13|||1||702163000107564368|0
M76|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|2913|Yellow|Project Big|2009-02-24|2009-03-16|NaT||||95.7||1|1|1|1|F|Black||18|No|Mother|28216|4|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||36|28269||Married|Self-Employed, Entrepreneur|28202|0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|501621811|501622131|31|0|2|501621016|31|0|2|500344465|10|2|500004641||3|2||-2||-2|0|10|||7464|9|||1|500004640|7869308672550505300|0
M77|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|518|Yellow||2014-04-28|2014-05-30|2015-10-30|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17||2|2|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28216|8|Two Parent|$35,000 to $39,999|||Y|Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||37|28031|Masters Degree|Single|Business: Mgt, Admin|94103|1|1|BBBS National Site|Web Link|Big|General Community|VOL - Mentoring Hispanic Youth|Enrollment|1|0|1|0|277|60|598|500000170|500008321|503026933|503028507|38|0|2|503758613|1|0|2|500761412|10|2|-2||4|2|500011312|-2|500011312|-2|0|10|||46|2|||1||9134125726462845918|7044657180546140448
M78|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4234|Green|Amachi|2004-06-03|2004-06-03|2016-01-06|Child: Graduated|Child: Graduated||139.1||1|1|1|1|M|Black||18|Yes|Mother|28208|8|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||51|28256|High School Graduate|Married|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500018987|500186645|500188043|31|0|1|500189545|31|0|2|500037636|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|0|0
M79|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2155|Green|Cabarrus County|2011-04-13|2011-04-13|NaT||||70.8||2|2|2|2|F|Black||18|Yes|Mother|28025|9|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|F|Black||43|28027||Divorced|Finance: Banking||0|7|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|500887862|500888132|31|0|2|500923430|31|0|2|500530980|10|2|500016307||2|1|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|500016374|5826822768343582573|0
M80|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1496|Green||2013-01-24|2013-01-31|NaT||||49.1||1|1|1|1|M|Black||18|No|Mother|28215|12|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|Black||41|28105|Bachelors Degree|Single|Tech: Management|28202|0|6|AA Task Force|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|502839827|502841119|31|0|1|503311280|31|0|1|500677083|10|2|-2||2|1||-2||-2|0|10|||6247|12|||1||6875312010577189564|3714886275549507192
M81|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|350|Green||2014-10-06|2014-10-06|2015-09-21|Child: Changed school/site|Child: Changed school/site||11.5||1|1|1|1|F|Hispanic||18|Yes|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||27|28202|Masters Degree|Single|Business||2|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504031009|504033027|3|0|2|503971990|1|0|2|500780903|10|1|500014504||4|1||-1|500014506|-1|0|4|||7462|13|||1||702163000107564368|0
M82|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2797|Green||2009-06-25|2009-07-10|NaT||||91.9||1|1|1|1|M|Black||18|No|Mother|28213|8|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||35|28209|Bachelors Degree|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|501604443|501604760|31|0|1|501729878|1|0|1|500371104|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||3677730851176818072|0
M83|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3221|Green||2007-07-23|2007-08-21|2016-06-15|Child: Graduated|Child: Graduated||105.8||1|1|1|1|M|Black||18|No|Mother|28226|6|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|M|Some Other Race||35|28209|||Business: Sales||0|0|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|500826594|500826861|31|0|1|500920342|41|0|1|500185735|10|2|-2||4|1||-2||-2|0|5|||6450|12|||1||0|0
M84|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2944|Green||2009-02-09|2009-02-13|NaT||||96.7||1|1|2|2|M|Multi-race (Black & White)||18|No|Mother|28213|9|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Mgt, Admin|28215|10|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501378357|501378636|36|0|1|501174997|31|0|1|500339619|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||253338316288302752|0
M85|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1688|Yellow|Cabarrus County|2012-05-22|2012-07-23|NaT||||55.5||1|1|1|1|M|Black||18|No|Mother|28025|10|One Parent: Female|$35,000 to $39,999|Yes: Active|No||Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||48|28269|Some College|Married|Tech: Management|28204|10|0|AA Task Force|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502578459|502578962|31|0|1|502869485|31|0|1|500615803|10|2|500016307||2|2|500016374|-2|500016374|-2|6854|8|||9229|13|||1|500016374|4170438818698997252|0
M86|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1276|Green||2011-11-14|2011-11-15|2015-05-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||41.9||1|1|1|1|M|White||18|No|Mother|28105|6|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||30|28211|Bachelors Degree|Single|Finance: Accountant|28204|0|5|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017777|502604900|502605417|1|0|1|502582742|1|0|1|500577855|10|2|-2||4|1||-2|500000294|-2|6854|8|||7464|9|||1||8545312001163392820|0
M87|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1309|Red||2013-02-19|2013-02-25|2016-09-26|Child/Family: Moved|Child/Family: Moved||43||1|1|1|1|M|Black||18|No|Mother|28216|8|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||33|28209|Bachelors Degree|Married|Business: Mgt, Admin|28202|6|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502974629|502976067|31|0|1|503188801|1|0|1|500682863|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||9134125726462845918|887254134148570071
M88|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3226|Green||2008-05-06|2008-05-07|NaT||||106||1|1|1|1|F|White||18|No|Father|28207|4|One Parent: Male|Unknown||||No||Self|General Community||Match Support|F|White||33|28226||Single|Human Services: Non-Profit|28205|0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501212047|501212321|1|0|2|501242250|1|0|2|500264889|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||0|0
M89|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1415|Green||2013-04-02|2013-04-22|NaT||||46.5||1|1|1|1|M|Black||18|Yes|Mother|28262|8|One Parent: Female|$45,000 to $49,999|||Y|No||Self|General Community||Match Support|M|White||31|28203|Masters Degree|Single|Consultant||0|9|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503110827|503112489|31|0|1|503278385|1|0|1|500691045|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||0|7674215580094440446
M90|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1334|Red||2011-10-07|2011-11-11|2015-07-07|Agency: Concern with Volunteer re: child safety|Agency: Concern with Volunteer re: child safety||43.8||1|1|1|1|M|White||18|No|Mother|28210|10|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||39|28210|Masters Degree|Single|Finance|28106|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|502499851|502500300|1|0|1|502690262|1|0|1|500562789|10|2|-2||4|3||-2||-2|0|10|||46|2|||1||5493390640808358320|0
M91|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-11-06|2015-11-06|NaT||||16||1|1|3|3|M|Black||18|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||45|28262|Bachelors Degree|Married|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504447856|504450112|31|0|1|502087592|31|0|1|500856992|10|1|500014504||2|1||-1|500014505, 500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M92|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|168|Green||2014-10-06|2014-11-03|2015-04-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||5.5||1|1|3|3|F|Black||18|No|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||36|28078|Masters Degree|Married|Business: Marketing|28273|1|1|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504042248|504044266|31|0|2|502056302|31|0|2|500780778|10|1|500014504||4|1||-1|500014505, 500014506|-1|0|4|||7671|13|||1||702163000107564368|0
M93|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|806|Green||2013-05-07|2013-05-22|2015-08-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||26.5||1|1|2|2|M|Black||17|No|Mother|28215|8|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||54|28262|Bachelors Degree|Married|Business||7|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500017732|502982301|502983753|31|0|1|503442370|31|0|1|500695892|10|2|-2||4|1||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1||0|0
M94|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1206|Yellow||2012-03-30|2012-04-30|2015-08-19|Volunteer: Moved|Volunteer: Moved||39.6||1|1|1|1|M|Black||17|No|Mother|28214|7|One Parent: Female|Less than $10,000||||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||32|28214|Bachelors Degree|Married|Self-Employed, Entrepreneur|29715|0|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502319972|502320407|31|0|1|502911091|1|0|1|500607368|10|2|-2||4|2|500005291|-2||-2|6854|8|||7464|9|||1||806697982905023857|3482130045776789614
M95|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3239|Green|Amachi|2008-02-27|2008-04-24|NaT||||106.4||1|1|1|1|M|Black||17|Yes|Mother|28212|11|One Parent: Female|Less than $10,000|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||46|28215|Bachelors Degree|Single|Business: Mgt, Admin|28226|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500814240|500814509|31|0|1|500981509|31|0|1|500248568|10|2|500003586||2|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294|1010189231295710785|0
M96|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|388|Green||2014-10-14|2014-10-20|2015-11-12|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||12.7||2|2|2|2|M|Black||17|No|Mother|28208|9|Two Parent|Unknown||||No||School|General Site|mentor2.0 2014|Match Support|M|Black||39|28269|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Site|mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500016847|500187081|500187961|31|0|1|500189197|31|0|1|500783502|10|1|500014504||4|1|500014506|-1|500014506|-1|0|4|||7464|9|||1||702163000107564368|0
M97|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|238|Green||2014-10-14|2014-10-16|2015-06-11|Volunteer: Moved|Volunteer: Moved||7.8||1|1|1|1|F|Hispanic||17|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site|mentor2.0 2014|RTBM|F|White||41|28277||Married|Finance: Banking|28202|0|0|Self|Self|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504070330|504072358|3|0|2|504032595|1|0|2|500783500|7|1|500014504||4|1|500014506|-1|500014506|-1|0|4|||7464|9|||1||702163000107564368|0
M98|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2405|Green||2010-01-21|2010-01-28|2016-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||79||1|1|1|1|M|Black||17||Mother|28215|11|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||54|28203|||Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017777|501936316|501936714|31|0|1|501872326|1|0|1|500428557|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||0|0
M99|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1487|Red||2013-01-15|2013-01-31|2017-02-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||48.9||1|1|1|1|M|Hispanic||17|No|Mother|28277|8|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Asian||30|28277|Bachelors Degree|Single|Finance||1|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020753|503026286|503027860|3|0|1|503259120|4|0|1|500674960|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||3966805366522644621|8598768071652363430
M100|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|86|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-11-02|2016-01-27|Child/Family: Time constraints|Child/Family: Time constraints||2.8||1|1|2|2|F|Hispanic||17|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|White||35|28205|Masters Degree|Married|Education: Teacher|28205|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504425940|504428195|3|0|2|502716664|1|0|2|500851872|10|1|500014504||4|1|500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M101|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1072|Red||2012-09-07|2012-10-17|2015-09-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||35.2||1|1|1|1|F|Black||17|No|Mother|28227|9|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||26|28269|Bachelors Degree|Single|Business|28262|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|501000843|501001116|31|0|2|503106526|31|0|2|500632934|10|2|-2||4|3||-2||-2|34|2|||7496|10|||1||8029775806705219538|7044657180546140448
M102|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|246|Green||2014-10-22|2014-10-22|2015-06-25|Child: Changed school/site|Child: Changed school/site||8.1||1|1|1|1|M|Black||17|No|Mother|28208|8|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Site|mentor2.0 2014|Match Support|M|White||42|28105|Masters Degree|Married|Librarian|28202|11|0|Neighbor/Friend|Neighbor/Friend|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500016847|502277840|502278010|31|0|1|503953636|1|0|1|500786451|10|1|500014504||4|1|500014506|-1|500014505, 500014506|-1|0|3|||7496|10|||1||702163000107564368|8325788680696113408
M103|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1140|Green||2014-01-06|2014-01-10|2017-02-23|Volunteer: Moved|Volunteer: Moved||37.5||1|1|1|1|M|White||17|No|GrandMother|28278|10|One Parent: Female|$20,000 to $24,999||||No||Self|General Community||Match Support|M|White||37|29708|Bachelors Degree|Single|Real Estate: Realtor|28273|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020910|503671116|503673077|1|0|1|503672609|1|0|1|500741347|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||7501346876523517480|0
M104|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Yellow||2014-03-06|2014-03-28|2016-08-26|Volunteer: Time constraint|Volunteer: Time constraint||29||2|2|1|1|F|Multi-race (Black & White)||17|No|Mother|28134|7|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|Black||48|28269|Masters Degree|Single|Education: Admin|28213|13|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017777|503013779|503724588|36|0|2|501311929|31|0|2|500753159|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1||5493390640808358320|3402014428779854546
M105|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2540|Green|Project Big|2010-03-18|2010-03-24|NaT||||83.4||1|1|1|1|M|Multi-race (Black & Hispanic)||17|No|Mother|28214|10|One Parent: Female|Unknown||||No|TV|Media|General Community|Project Big|Match Support|M|White||34|28164|Masters Degree||Finance|28210|3|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501919423|501919819|38|0|1|502034798|1|0|1|500442066|10|2|500004641||2|1|500004640|-2||-2|56|1|||7464|9|||1|500004640|216500609169513656|0
M106|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-09-23|2015-10-26|NaT||||16.4||2|2|2|2|M|Black||17|No|Mother|28217|9|One Parent: Female|Unknown||||No||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|White||52|28105|Bachelors Degree|Married|Business||2|6|Local Print|Media|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500022907|504031043|504033061|31|0|1|503776239|1|0|1|500841767|10|1|500014504||2|1|500014505, 500015184|-1|500014505, 500014506|-1|0|4|||7439|1|||1|500014505, 500015184|702163000107564368|0
M107|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|324|Green||2014-10-07|2014-10-07|2015-08-27|Volunteer: Time constraint|Volunteer: Time constraint||10.6||2|2|2|2|M|Black||17|No|Mother|28217|9|One Parent: Female|Unknown||||No||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Black||34|28269|Some College|Married|Business|28025|5|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504031043|504033061|31|0|1|503956879|31|0|1|500781238|10|1|||4|1|500014505, 500015184|-1|500014506, 500016374|-2|0|4|||7671|13|||1||702163000107564368|0
M108|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|4004|Green|Cabarrus County|2006-03-21|2006-03-21|NaT||||131.5||2|2|1|1|F|White||17|No|Mother|28027|8|Two Parent|Unknown||||No||Relative|General Community|Cabarrus County|Match Support|F|White||32|28146|Bachelors Degree|Single|Human Services: Social Worker||0|0|other|College Partner|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|500361200|500361450|1|0|2|500368628|1|0|2|500085591|10|2|500016307||2|1|500016374|-2|500016374|-2|0|3|||7670|5|||1|500016374|5273065343662533495|0
M109|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3232|Green||2008-05-01|2008-05-01|NaT||||106.2||1|1|1|1|M|Black||17|No|Mother|28277|9|One Parent: Female|$40,000 to $44,999||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||36|28270|Juris Doctorate (JD)|Married|Law: Lawyer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500378354|500378596|31|0|1|501181060|1|0|1|500264206|10|2|-2||2|1||-2||-2|6854|8|||46|2|||1||4102911263088044|0
M110|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1424|Yellow|2010-2012 OJJDP JJI|2011-03-29|2011-04-11|2015-03-05|Child: Lost interest|Child: Lost interest||46.8||3|3|1|1|F|Black||17||Mother|28215|8|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28215|High School Graduate|Married|Finance: Banking|28255|13|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500012459|501011735|500417756|31|0|2|502473442|31|0|2|500528270|10|2|-2||4|2|500005291|-2||-2|0|10|||7446|3|||1|500005291|6724463016047116758|0
M111|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1315|Red|Amachi|2012-01-11|2012-01-23|2015-08-30|Volunteer: Moved|Volunteer: Moved||43.2||1|1|1|1|F|Black||17|Yes|Mother|28273|7|One Parent: Female|$30,000 to $34,999||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||31|28217||Single|Customer Service||0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502725777|502726673|31|0|2|502710032|31|0|2|500590950|10|2|-2||4|3|500000294|-2||-2|34|2|||7464|9|||1|500000294|8567789404096574827|4376931673251632105
M112|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1425|Yellow||2012-06-25|2012-06-25|2016-05-20|Volunteer: Time constraint|Volunteer: Time constraint||46.8||2|2|3|3|M|Black||17||Mother|28210|5|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28277|Bachelors Degree|Married|Business||0|0|Michael Baisden|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502530688|502531141|31|0|1|502166996|31|0|1|500621632|10|2|-2||4|2|500005291|-2||-2|0|3|||11272|1|||1||5386346637278076349|0
M113|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3469|Green||2007-09-05|2007-09-07|NaT||||114||1|1|1|1|M|Black||17|No|Mother|28277||One Parent: Female|$60,000 to $74,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||58|28270|Bachelors Degree|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500931662|500931932|31|0|1|500894084|1|0|1|500193824|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1||0|0
M114|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|924|Yellow||2014-01-08|2014-01-17|2016-07-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||30.4||1|1|1|1|M|Black||17|No|Mother|28270|9|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||32|28226|Bachelors Degree|Married|Consultant|28202|4|4|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|503662199|503664159|31|0|1|503639494|1|0|1|500741727|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1||1010189231295710785|0
M115|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2213|Green|Amachi|2011-01-20|2011-02-14|NaT||||72.7||1|1|1|1|F|Black||17|Yes|Relative: Other|28227|5|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||34|28212|Masters Degree|Single|Education: Teacher|28216|6|3|Self|Self|Big|General Community|Amachi, Project Big|Match Support|1|0|0|1|277|60|598|500000170|500020752|502255150|502255582|31|0|2|502392989|1|0|2|500512287|10|2|500003586||2|1|500000294|-2|500000294, 500004640|-2|0|5|||7464|9|||1|500000294|0|0
M116|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2380|Red||2010-04-26|2010-05-07|2016-11-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||78.2||1|1|1|1|F|Black||17|No|Mother|28083||One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi, Cabarrus County|Match Support|F|Black||39|28269||Single|Self-Employed, Entrepreneur|28027|7|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500020753|501716763|501716992|31|0|2|502112513|31|0|2|500449029|10|2|-2||4|3|500000294, 500016374|-2|500016374|-2|6854|8|||7458|9|||1||0|0
M117|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|4618|Green|Amachi|2004-07-15|2004-07-15|NaT||||151.7||1|1|1|1|F|Black||17|Yes|Mother|28217|11|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||73|28203||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|500186952|500188132|31|0|2|500189723|1|0|2|500037836|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|702163000107564368|0
M118|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1099|Green||2013-01-11|2013-01-24|2016-01-28|Volunteer: Moved|Volunteer: Moved||36.1||1|1|1|1|M|Black||17|No|Mother|28210|7|One Parent: Female|$40,000 to $44,999|||Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||32|28203|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502839019|502840311|31|0|1|502432390|31|0|1|500674451|10|2|-2||4|1||-2||-2|6854|8|||7496|10|||1||6202343250032725030|5468286809853673926
M119|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1616|Red||2011-11-30|2011-12-21|2016-05-24|Child: Graduated|Child: Graduated||53.1||1|1|2|2|F|Black||17|No|Mother|28083|9|One Parent: Female|$60,000 to $74,999||||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500020753|502702145|502702991|31|0|2|502204211|31|0|2|500582836|10|2|-2||4|3||-2||-2|6854|8|||7464|9|||1||0|3402014428779854546
M120|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|623|Yellow||2014-06-02|2014-06-20|2016-03-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.5||1|1|1|1|M|Black||17|No|Mother|28216|8|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|White||31|28262|Bachelors Degree|Single|Tech: Engineer|28262|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|503360420|503362265|31|0|1|503831013|1|0|1|500765209|10|2|-2||4|2||-2||-2|0|10|||46|2|||1||540227296891876425|8983800016848597675
M121|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2126|Green|Amachi, Project Big, Project Big AND Amachi|2011-04-30|2011-04-30|2017-02-23|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||69.8||1|1|1|1|F|Black||17|Yes|Mother|28206|5|Other/Unknown|Unknown||||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||61|28134|Bachelors Degree|Married|Medical: Admin||33|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|1|0|1|0|277|60|598|500000170|500020910|502570183|502570637|31|0|2|502570153|31|0|2|500534090|10|2|500004772||4|1|500000294, 500004640, 500004901|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|500000294, 500004640, 500004901|7869308672550505300|0
M122|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1701|Green||2012-06-13|2012-07-10|NaT||||55.9||4|4|1|1|F|Black||17|Yes|Mother|28227|10|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|F|Black||47|28269|Bachelors Degree|Single|Law: Paralegal|28202|0|4|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|500243491|500188056|31|0|2|502919490|31|0|2|500619145|10|2|-2||2|1|500000294|-2||-2|0|4|||7464|9|||1||1766165378108010922|0
M123|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2337|Green||2010-09-30|2010-10-13|NaT||||76.8||1|1|1|1|F|Black||17|No|Mother|28269|12|Two Parent|Unknown||||Yes||Relative|General Community||Match Support|F|Multi-race (Asian & White)||33|28205|Masters Degree|Married|Finance: Economist|28223|7|0|Newspaper|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502172536|502172965|31|0|2|501279665|37|0|2|500475431|10|2|-2||2|1||-2||-2|0|3|||129|1|||1||2374609189072499123|0
M124|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1068|Green||2014-03-20|2014-04-04|NaT||||35.1||2|2|2|2|F|Black||17|Yes|Mother|28216|10|One Parent: Female|Unknown|||Y|Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|502180719|502181148|31|0|2|502391505|31|0|2|500755816|10|2|500003586||2|1|500000294|-2|500000294|-2|7016|11|||7438|1|||1||216500609169513656|0
M125|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1623|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-05-12|2011-05-20|2015-10-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||53.3||1|1|1|1|F|Black||17|No|Mother|28217|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||42|28210||Single|Business: Human Resources||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502551092|502551545|31|0|2|502366844|1|0|2|500536172|10|2|-2||4|2|500004640, 500005291|-2||-2|0|4|||10326|3|460|3|1|500004640, 500005291|5493246288421413675|0
M126|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1093|Green|Cabarrus County|2014-01-28|2014-03-10|NaT||||35.9||2|2|3|3|F|Black||17|No|Mother|28083|12|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|Black||41|28027|PHD|Single|Medical: Doctor, Provider|28075|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502670076|502670904|31|0|2|501391123|31|0|2|500745456|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|7659437100141520816|0
M127|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2976|Green||2008-12-08|2009-01-12|NaT||||97.8||2|2|1|1|M|Black||17|No|Mother|28215|8|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||32|28208|Associate Degree|Single|Service: Restaurant|28211|4|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500938154|500938424|31|0|1|501446421|1|0|1|500323753|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||6202343250032725030|0
M128|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|350|Green||2014-10-06|2014-10-06|2015-09-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||11.5||1|1|3|3|F|Hispanic||17|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Asian||32|28105|Bachelors Degree|Married|Librarian|28227|9|0|Neighbor/Friend|Neighbor/Friend|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500016847|504043289|504045307|3|0|2|502366876|4|0|2|500780880|10|1|500014504||4|1||-1|500014505, 500014506|-1|0|4|||7496|10|||1||702163000107564368|0
M129|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|461|Green||2015-12-02|2015-12-02|NaT||||15.1||2|2|4|4|F|Black||17|Yes|GrandMother|28273|10|Grandparents|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|501300013|500561354|31|0|2|500346193|31|0|2|500864495|10|2|-2||2|1|500000294|-2||-2|7294|13|||46|2|||1||5493390640808358320|0
M130|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|3100|Yellow||2008-09-03|2008-09-10|NaT||||101.8||3|3|1|1|F|Black||17|No|Mother|28227|5|One Parent: Female|$35,000 to $39,999||||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black|Other African|44|28212||Single|Consultant||1|5|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500970495|500970766|31|0|2|500965698|31|31|2|500285645|10|2|-2||3|2||-2||-2|7294|13|||46|2|||1||0|0
M131|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2351|Green|Amachi|2010-08-31|2010-09-29|NaT||||77.2||1|1|1|1|F|Black||17|Yes|Mother|28269||One Parent: Female|$30,000 to $34,999|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||61|28204||Divorced|Self-Employed, Entrepreneur||0|0|Billboard|Media|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|500970267|500970535|31|0|2|502084649|1|0|2|500468192|10|2|500003586||2|1|500000294|-2|500000294|-2|5635|9|||125|1|||1|500000294|0|0
M132|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1880|Green||2011-12-14|2012-01-13|NaT||||61.8||1|1|1|1|M|Black||17|No|Mother|28212|6|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|Black||45|28207|Masters Degree|Married|Tech: Management|28081|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502571727|502572181|31|0|1|502769619|31|0|1|500586830|10|2|-2||3|1||-2||-2|0|10|||7671|13|||1||0|0
M133|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3457|Green|Amachi, Cabarrus County|2007-09-05|2007-09-19|NaT||||113.6|Y|1|1|1|1|M|Black||17|Yes|Mother|28212|9|One Parent: Female|$40,000 to $44,999|||Y|No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|Black||62|28213||Married|Finance: Economist||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|500958307|500958577|31|0|1|500876132|31|0|1|500193868|10|2|500003586||2|1|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|500000294, 500016374|1766165378108010922|0
M134|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|751|Red||2013-11-13|2013-12-09|2015-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.7||1|1|1|1|F|White||17|No|Father|28269|9|Two Parent|$100,000 to $124,999|||Y|No||Relative|General Community||Match Support|F|White||29|28205|Some College|Single|Business: Mgt, Admin|29707|3|10|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|503417576|503419440|1|0|2|503594017|1|0|2|500730510|10|2|-2||4|3||-2|500000294|-2|0|3|||7464|9|||1||1652521212990559348|8243619853090168866
M135|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1034|Yellow||2013-07-16|2013-07-26|2016-05-25|Child: Lost interest|Child: Lost interest||34||1|1|2|3|M|Black||17|No|Mother|28216|11|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|Black||40|28202|Bachelors Degree|Single|Consultant|28281|4|5|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500013781|503255669|503257474|31|0|1|500188812|31|0|1|500703771|10|2|-2||4|2||-2|500000294|-2|0|10|||2238|7|||1||7301546317881317703|1283000929024117684
M136|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1623|Green||2011-11-28|2011-12-07|2016-05-17|Child: Lost interest|Child: Lost interest||53.3||1|1|1|1|F|Black||17|No|Mother|28269|9|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Sales||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|502674024|502674852|31|0|2|502660051|1|0|2|500581910|10|2|-2||4|1|500005291|-2||-2|0|10|||7496|10|||1||7301546317881317703|0
M137|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1300|Yellow||2012-06-12|2012-06-30|2016-01-21|Child: Lost interest|Child: Lost interest||42.7||3|4|1|1|F|Black||17||Relative: Other|28206|11|Grandparents|Unknown||||Yes||School|General Community|Amachi|Match Support|F|Black||37|28215|Masters Degree|Single|Education: Admin|28273|0|10|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500020752|501157075|501157349|31|0|2|502978065|31|0|2|500619009|10|2|-2||4|2|500000294|-2||-2|0|4|||7464|9|||1||2374609189072499123|0
M138|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|501|Red||2014-08-21|2014-09-15|2016-01-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.5||1|1|1|1|F|Black||17|No|Mother|28208|11|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Multi-race (Black & Hispanic)||59|28216|Some College|Divorced|Law: Legal Secretary|28202|14|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503804225|503805695|31|0|2|503881040|38|0|2|500773105|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1||253338316288302752|6993050796559809579
M139|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3098|Green|Amachi|2008-08-11|2008-09-12|NaT||||101.8||1|1|1|1|F|Black||17|Yes|Mother|28227|10|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||46|27704|Associate Degree|Divorced|Medical: Admin||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|501309634|501309912|31|0|2|501046221|31|0|2|500281317|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||7462|13|||1|500000294|1010189231295710785|0
M140|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|631|Green||2014-01-15|2014-02-26|2015-11-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.7||1|1|1|1|M|Black||17|No|Mother|28226|8|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||34|28210|Masters Degree|Married|Real Estate: Realtor|28202|2|3|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|503448711|503450577|31|0|1|503576769|1|0|1|500742906|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||9134125726462845918|3535616089900023359
M141|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green|mentor2.0, mentor2.0 2016|2015-10-26|2015-11-11|NaT||||15.8||1|1|1|1|M|White||17|No|Step-Mother|28217|9|Two Parent|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|White||59|28226|Masters Degree|Married|Business|28226|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504493589|504495874|1|0|1|504314218|1|0|1|500851954|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500016394|702163000107564368|0
M142|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1772|Green||2012-04-19|2012-04-30|NaT||||58.2||1|1|1|1|M|Black||17|No|Mother|28211|11|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Black||47|28227|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502885468|502886874|31|0|1|502954219|31|0|1|500610806|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||7501346876523517480|0
M143|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1954|Green||2011-10-20|2011-10-31|NaT||||64.2||1|1|2|2|M|Black||17|No|Mother|28206|11|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502371558|502371997|31|0|1|502528355|1|0|1|500568298|10|2|-2||2|1|500000294, 500005291|-2||-2|0|10|||132|8|||1||2374609189072499123|0
M144|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1669|Green|Amachi|2011-03-03|2011-03-21|2015-10-15|Child: Lost interest|Child: Lost interest||54.8||1|1|1|1|F|Black||17|No|Mother|28262|6|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||26|28031|Bachelors Degree|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|502275241|502275673|31|0|2|502394690|1|0|2|500521625|10|2|500003586||4|1|500000294|-2||-2|0|10|||7496|10|||1|500000294|0|0
M145|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1593|Green|Cabarrus County|2012-10-16|2012-10-26|NaT||||52.3||2|2|2|2|F|Black||17|No|GrandMother|28027|8|Grandparents|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|Black||42|28213|Bachelors Degree|Single|Finance: Banking|28202|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502129650|502130079|31|0|2|502598777|31|0|2|500646243|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|6353565629814722343|0
M146|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2542|Green||2009-10-13|2009-10-29|2016-10-14|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|9|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020910|501725162|501724831|39|0|1|501833178|1|0|1|500394157|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||7432163260389731024|0
M147|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|666|Green||2014-03-18|2014-03-31|2016-01-26|Volunteer: Moved|Volunteer: Moved||21.9||1|1|1|1|M|Black||17|No|Mother|28226|9|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|Multi-race (Black & White)||29|28215|Some College|Married|Student: College|28223|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503124706|503126373|31|0|1|503609606|36|0|1|500755317|10|2|-2||4|1||-2||-2|0|10|||46|2|||1||4102911263088044|6991424324982091759
M148|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1799|Green||2012-03-28|2012-04-03|NaT||||59.1||1|1|1|1|M|Black||17|No|Mother|28278|6|Two Mothers|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||32|28278|Bachelors Degree|Single|Medical|28208|3|5|Relative|Relative|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502526965|502527418|31|0|1|502881104|1|0|1|500606886|10|2|-2||2|1||-2||-2|0|10|||17161|11|||1||0|0
M149|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1238|Yellow||2012-08-03|2012-08-17|2016-01-07|Volunteer: Time constraint|Volunteer: Time constraint||40.7||2|2|1|1|F|Black||17|No|GrandMother|28208||One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|RTBM|F|White||41|28105|Bachelors Degree|Divorced|Business|28112|1|3|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502431187|502431630|31|0|2|503015009|1|0|2|500627361|7|2|-2||4|2|500005291|-2||-2|0|5|||46|2|||1||3038247238543299436|0
M150|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|178|Yellow|PERL 2014-2016|2014-09-04|2014-09-29|2015-03-26|Child: Severity of challenges|Child: Severity of challenges||5.8||1|1|2|2|M|Black||17|No|Mother|28216|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Asian||33|28204|Bachelors Degree|Married|Business: Engineer|28007|3|9|Man Up Campaign|Media|Big|General Community|Amachi, PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500015820|503546374|503548249|31|0|1|503890372|4|0|1|500774577|10|2|-2||4|2|500014681|-2|500000294, 500014681|-2|0|4|||17101|1|||1|500014681|0|6054903719040220574
M151|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2286|Green|Amachi|2009-04-01|2009-04-30|2015-08-03|Volunteer: Time constraint|Volunteer: Time constraint||75.1||2|2|1|1|F|Black||17|Yes|Mother|28227|9|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||31|28204|Bachelors Degree|Single|Business: Engineer|28269|0|2|TV|Media|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500011349|500271303|500271368|31|0|2|501291358|1|0|2|500354049|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||130|1|||1|500000294|3292090474897428830|0
M152|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|NaT||||16||1|1|1|1|M|Hispanic||17|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||31|28209|Masters Degree|Separated|Business: Marketing||5|5|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504447951|504450207|3|0|1|504272897|1|0|1|500846253|10|1|500014504||2|1||-1|500015184|-1|0|4|||17159|12|||1|500014505, 500015184|702163000107564368|0
M153|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3653|Green||2007-03-02|2007-03-07|NaT||||120||1|1|1|1|F|Black||17||Mother|28213|10|One Parent: Female|Less than $10,000|||Y|No||School|General Community||Match Support|F|Black||32|28214|Bachelors Degree|Married|Architect|28270|0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|500724632|500724899|31|0|2|500803551|31|0|2|500164708|10|2|-2||2|1||-2||-2|0|4|||46|2|||1||7432163260389731024|0
M154|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1443|Green||2013-03-25|2013-03-25|NaT||||47.4||2|2|2|2|F|Black||17|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502124485|502142970|31|0|2|501905673|31|0|2|500689671|10|2|-2||2|1||-2||-2|0|4|||7496|10|||1||702163000107564368|0
M155|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|882|Green|mentor2.0, mentor2.0 2014|2014-10-07|2014-10-07|NaT||||29||1|1|2|2|F|Black||17|Yes|Mother|28217||One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Asian||32|28209|PHD|Single|Business: Marketing|28223|1|2|Self|Self|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504042320|504044338|31|0|2|502779828|4|0|2|500781152|10|1|500014504||2|1||-1|500014505, 500014506|-1|0|4|||7464|9|||1|500014505, 500014506|702163000107564368|0
M156|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1429|Green|Project Big|2011-11-29|2011-11-30|2015-10-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||46.9||2|2|1|1|F|Black||17||Mother|28208|5|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28205|Bachelors Degree|Married|Business|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017777|502589869|502590381|31|0|2|502701252|1|0|2|500582617|10|2|500004641||4|1|500004640, 500005291|-2|500000294|-2|0|4|459|3|7496|10|||1|500004640|7869308672550505300|0
M157|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1534|Red||2012-03-23|2012-04-05|2016-06-17|Volunteer: Moved|Volunteer: Moved||50.4||1|1|1|1|F|Black||17|No|Mother|28216|10|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Business: Marketing|28203|0|8|Other Church Partner|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502912141|502913549|31|0|2|502932948|1|0|2|500605880|10|2|-2||4|3||-2||-2|34|2|||7453|7|||1||253338316288302752|3402014428779854546
M158|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2062|Green|2010-2012 OJJDP JJI|2011-02-04|2011-02-10|2016-10-03|Volunteer: Moved|Volunteer: Moved||67.7||1|1|1|1|M|Black||17|No|Mother|28212|7|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28202|Bachelors Degree|Single|Business: Sales|27560|1|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|1|0|1|0|277|60|598|500000170|500017732|502197477|502197915|31|0|1|502422929|1|0|1|500515536|10|2|-2||4|1|500005291|-2|500000294, 500004640|-2|0|4|||7464|9|||1|500005291|2811191761055817959|8113241890313112769
M159|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1349|Red|Amachi|2011-09-22|2011-10-13|2015-06-23|Child: Lost interest|Child: Lost interest||44.3||1|1|1|1|M|Black||17|Yes|GrandMother|28216|8|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||47|28216|Bachelors Degree|Married|Business: Engineer|28255|18|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500013781|502206673|502207102|31|0|1|502668179|1|0|1|500557233|10|2|500003586||4|3|500000294|-2||-2|0|10|||7464|9|||1|500000294|9134125726462845918|0
M160|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|336|Green||2014-10-08|2014-11-03|2015-10-05|Child/Family: Moved|Child/Family: Moved||11||1|1|2|2|F|Black||17|No|Mother|28273|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||39|28273|Masters Degree|Married|Business: Mgt, Admin|28208|2|0|BBBS National Site|Web Link|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043455|504045473|31|0|2|503972115|31|0|2|500781712|10|1|500014504||4|1||-1|500014506|-1|0|4|||46|2|||1||702163000107564368|0
M161|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green|mentor2.0, mentor2.0 2016|2015-10-25|2015-11-11|NaT||||15.8||1|1|1|1|M|Black||17|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Black||52|29708|Masters Degree|Single|Tech: Management||30|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454538|504456796|31|0|1|504311707|31|0|1|500851883|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||17159|12|||1|500014505, 500016394|702163000107564368|0
M162|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|136|Green|mentor2.0, mentor2.0 2015|2016-05-31|2016-05-31|2016-10-14|Child: Severity of challenges|Child: Severity of challenges||4.5||1|1|2|2|M|Black||17|No|GrandMother|28212|9|Grandparents|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|M|White||34|28210|Bachelors Degree|Married|Medical||3|6|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500021786|504513842|504516137|31|0|1|504431507|1|0|1|500895194|10|1|500014504||4|1|500015184|-1|500016394|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M163|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2965|Green|Amachi|2008-12-19|2009-01-23|NaT||||97.4||1|1|1|1|M|White||17|Yes|Mother|28227|9|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||54|28227|Bachelors Degree|Divorced|Business: Sales|28273|9|5|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|501361902|501249611|1|0|1|501307192|1|0|1|500328424|10|2|500003586||2|1|500000294|-2||-2|0|10|||46|2|||1|500000294|3292090474897428830|0
M164|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|580|Red||2013-09-10|2013-09-20|2015-04-23|Child: Lost interest|Child: Lost interest||19.1||1|1|1|1|M|Black||17|No|Mother|28212|9|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||63|28210|Bachelors Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503476243|503478109|31|0|1|503334174|1|0|1|500710120|10|2|-2||4|3||-2||-2|0|10|||7671|13|1561|2|1||2811191761055817959|887254134148570071
M165|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1714|Green||2012-06-15|2012-06-27|NaT||||56.3||1|1|1|1|M|Black||17|No|Mother|28217|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Black||41|28210|Bachelors Degree|Separated|Arts, Entertainment, Sports|28202|2|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502700505|502701350|31|0|1|503029324|31|0|1|500619505|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||194235582162093094|0
M166|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3012|Green||2008-06-23|2008-07-02|2016-09-30|Volunteer: Time constraint|Volunteer: Time constraint||99||3|3|1|1|F|Multi-Race (None of the above)||17||Mother|28215|11|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Match Support|F|Black||43|28208|Masters Degree|Single|Business: Sales|28078|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500545328|500545578|7|0|2|501033808|31|0|2|500274449|10|2|-2||4|1||-2||-2|0|10|||46|2|||1||1652521212990559348|0
M167|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3596|Red||2006-10-29|2006-10-29|2016-09-02|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||118.1|Y|1|1|1|1|M|Multi-Race (None of the above)||17||Mother|28215|10|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Match Support|M|Black||55|28214||Married|Clergy||12|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500545326|500545578|7|0|1|500697845|31|0|1|500134545|10|2|-2||4|3||-2||-2|0|10|||2238|7|||1||6875312010577189564|0
M168|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1651|Red||2012-01-11|2012-02-11|2016-08-19|Volunteer: Moved|Volunteer: Moved||54.2||1|1|1|1|F|Black||17|No|Mother|28083|7|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Cabarrus County|Match Support|F|Black||29|28027|Bachelors Degree|Single|Education: Teacher||1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500020753|502083429|502083853|31|0|2|502653045|31|0|2|500590992|10|2|-2||4|3|500016374|-2|500016374|-2|7016|11|||7464|9|||1||675996018716794055|0
M169|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2032|Red|Amachi|2009-06-24|2009-07-08|2015-01-30|Child/Family: Moved|Child/Family: Moved||66.8||1|1|1|1|F|Black||17|Yes|Mother|28212|3|One Parent: Female|Unknown||||Yes|YeaGod|Faith Organization|General Community|Amachi|Match Support|F|Black||51|28262|PHD|Married|Real Estate: Realtor||0|0|Weeping Willow|Faith Organization|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008321|501726201|501726541|31|0|2|501734664|31|0|2|500371036|10|2|-2||4|3|500000294|-2||-2|5634|9|||9218|7|||1|500000294|0|0
M170|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|625|Green||2014-04-30|2014-05-12|2016-01-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.5||1|1|1|1|F|Black||17|No|Mother|28208|8|Two Parent|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||38|28262|Masters Degree|Single|Finance|28262|0|6|Agency Sponsored|Special Event|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500018851|503833956|503835911|31|0|2|503635291|31|0|2|500761770|10|2|-2||4|1||-2|500000294|-2|34|2|||16426|8|||1||2611337051335117774|3630529025150538848
M171|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|883|Green||2014-09-17|2014-10-06|NaT||||29||4|4|1|1|M|Black||17|Yes|Mother|28213|11|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||39|28269|Bachelors Degree|Married|Arts, Entertainment, Sports|28202|15|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501786018|501786373|31|0|1|503914867|31|0|1|500776457|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||7301546317881317703|0
M172|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2476|Green||2009-03-19|2009-04-01|2016-01-11|Volunteer: Time constraint|Volunteer: Time constraint||81.3||1|1|3|4|F|Black||17|No|Mother|28216|10|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28269|||Business: Marketing||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|501376745|501377024|31|0|2|500725077|31|0|2|500350905|10|2|-2||4|1||-2||-2|6854|8|||46|2|||1||216500609169513656|682544529818549127
M173|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|883|Green|mentor2.0, mentor2.0 2014|2014-10-06|2014-10-06|NaT||||29||1|1|2|2|F|Black||17|No|Mother|28273|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||33|28215|Bachelors Degree|Single|Tech: Support, Writing|28204|6|0|Other|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504043477|504045495|31|0|2|501245666|31|0|2|500780765|10|1|500014504||2|1||-1|500014506|-2|0|4|||7671|13|||1|500014505, 500014506|702163000107564368|0
M174|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1235|Green||2013-10-09|2013-10-19|NaT||||40.6||1|1|2|2|F|Black||17|No|Mother|28216||One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503533026|503534897|31|0|2|502485670|31|0|2|500717656|10|2|-2||2|1||-2||-2|0|10|||7462|13|1204|3|1||3935539763241716148|1786514887916898235
M175|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2433|Green||2010-06-30|2010-07-09|NaT||||79.9||1|1|1|1|M|Black||17|No|Mother|29732|10|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||52|28270|Bachelors Degree|Married|Business: Mgt, Admin||4|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502067798|502074089|31|0|1|502062408|1|0|1|500459576|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||0|0
M176|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1169|Green||2011-11-28|2012-01-23|2015-04-06|Volunteer: Time constraint|Volunteer: Time constraint||38.4||2|2|1|1|F|Black||17|No|Mother|28216|8|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||48|28031|Some College|Divorced|Medical|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501529921|501530213|31|0|2|502554719|1|0|2|500581908|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||0|0
M177|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|350|Green||2014-10-06|2014-10-06|2015-09-21|Child/Family: Moved|Child/Family: Moved||11.5||1|1|2|2|F|Black||17|No|Mother|28214|9|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Site||Match Support|F|White||54|28210|Masters Degree|Married|Tech: Computer/Programmer|28202|1|10|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|502702827|502703671|31|0|2|503969458|1|0|2|500780876|10|1|500014504||4|1||-1|500014506|-1|0|10|||7671|13|||1||702163000107564368|7044657180546140448
M178|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|475|Green|mentor2.0, mentor2.0 2015|2015-11-06|2015-11-18|NaT||||15.6||1|1|1|1|F|Hispanic||17|No|Mother|28211|9|One Parent: Female|$10,000 to $14,999||||Yes||Relative|General Site||Match Support|F|White||31|28210|Bachelors Degree|Single|Business|33716|8|1|Self|Self|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504495905|504498190|3|0|2|504366540|1|0|2|500857036|10|1|500014504||2|1||-1|500015184|-1|0|3|||7464|9|||1|500014505, 500015184|702163000107564368|0
M179|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|336|Green||2014-10-14|2014-10-20|2015-09-21|Child: Changed school/site|Child: Changed school/site||11||2|2|1|1|M|Black||17||Mother|28208|9|One Parent: Female|Unknown|||Y|No||School|General Site|mentor2.0 2014|Match Support|M|Black||30|28273|Bachelors Degree|Single|Business||3|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500016847|501083790|501084064|31|0|1|503984623|31|0|1|500783501|10|1|500014504||4|1|500014506|-1|500014506|-1|0|4|||7462|13|||1||702163000107564368|0
M180|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2226|Green||2009-01-08|2009-01-21|2015-02-25|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||73.1||1|1|1|1|M|Black||17|No|Mother|28212||One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|White||53|15001|Masters Degree|Single|Consultant|28202|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501428903|501429188|31|0|1|501441245|1|0|1|500331206|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||0|0
M181|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|w|S|Completed|Match Support|336|Green|mentor2.0 2015|2015-10-25|2015-11-30|2016-10-31|Child/Family: Time constraints|Child/Family: Time constraints||11||1|1|1|1|F|Asian||17|No|Mother|28208||One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|White||26|28278|Masters Degree|Living w/ Significant Other|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|0|1|1|0|277|60|598|500000170|500017786|504445088|504447344|4|0|2|504368282|1|0|2|500851870|10|1|500014504||4|1|500015184|-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M182|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|343|Green|mentor2.0, mentor2.0 2015|2015-10-14|2015-11-06|2016-10-14|Child: Severity of challenges|Child: Severity of challenges||11.3||1|1|1|1|M|Black||17|Yes|Mother|28217|9|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Site|mentor2.0, mentor2.0 2015|Match Support|M|White||35|28210|Masters Degree|Married|Business: Sales|29708|8|0|Gala|Special Event|Big|General Site|mentor2.0 2015|Enrollment|0|1|1|0|277|60|598|500000170|500021786|502133283|502133712|31|0|1|504277979|1|0|1|500847663|10|1|500014504||4|1|500014505, 500015184|-1|500015184|-1|0|5|||7457|8|||1|500014505, 500015184|702163000107564368|5941760529237532868
M183|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1087|Green||2013-08-07|2013-08-26|2016-08-17|Child: Lost interest|Child: Lost interest||35.7||1|1|1|1|F|Black||17|No|Mother|28203|10|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||29|28110|Masters Degree|Single|Education: Teacher||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503014417|503015947|31|0|2|503518076|1|0|2|500706096|10|2|-2||4|1||-2||-2|0|10|||46|2|||1||2374609189072499123|7044657180546140448
M184|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|233|Yellow|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-17|2016-07-07|Child/Family: Moved|Child/Family: Moved||7.7||1|1|2|2|M|Hispanic||17|No|Mother|28209|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||30|28207||Single|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015, mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500021786|504447755|504450011|3|0|1|504434419|1|0|1|500846217|10|1|500014504||4|2||-1|500015184, 500016394|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M185|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2178|Green|Amachi, Project Big, Project Big AND Amachi|2011-03-02|2011-03-21|NaT||||71.6||1|1|1|1|F|Black||17|Yes|Mother|28205|9|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||53|28031||Divorced|Medical: Admin|28207|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502307585|502308017|31|0|2|501519450|1|0|2|500521250|10|2|500004772||2|1|500000294, 500004640, 500004901|-2||-2|0|4|||7446|3|||1|500000294, 500004640, 500004901|1766165378108010922|0
M186|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|396|Green|mentor2.0, mentor2.0 2014|2014-10-06|2014-10-06|2015-11-06|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||13||1|1|1|1|F|Black||17|Yes|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||28|28210|Masters Degree|Single|Tech: Management|28277|3|2|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043271|504045289|31|0|2|503974114|31|0|2|500780793|10|1|500014504||4|1||-1|500014506|-1|0|4|||7671|13|||1|500014505, 500014506|702163000107564368|0
M187|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1271|Yellow||2012-09-27|2012-10-29|2016-04-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||41.8||1|1|1|1|M|Black||17|No|Mother|28269|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||34|28203|Juris Doctorate (JD)|Single|Law: Lawyer||2|11|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|502920861|502922278|31|0|1|503097126|1|0|1|500639233|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1||967246839551912690|0
M188|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2126|Green|Project Big, 2010-2012 OJJDP JJI|2011-04-26|2011-04-30|2017-02-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||69.8||1|1|1|1|F|Black||17|No|Mother|28216|5|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||56|28226|Masters Degree|Married|Medical: Nurse|28217|34|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|1|0|1|0|277|60|598|500000170|500020910|502570188|502570642|31|0|2|502366830|1|0|2|500533448|10|2|500004641||4|1|500004640, 500005291|-2|500004640|-2|0|4|||10326|3|||1|500004640, 500005291|7869308672550505300|0
M189|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|332|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-17|2016-10-14|Child/Family: Time constraints|Child/Family: Time constraints||10.9||1|1|1|1|F|Black||17|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||36|28214|Masters Degree|Single|Arts, Entertainment, Sports|28202|1|3|BBBS National Site|Web Link|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504447916|504450172|31|0|2|504130536|31|0|2|500846243|10|1|500014504||4|1||-1|500015184|-1|0|4|||46|2|||1|500014505, 500015184|702163000107564368|0
M190|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|112|Green|PERL 2014-2016|2014-09-22|2014-09-23|2015-01-13|Child/Family: Moved|Child/Family: Moved||3.7||2|2|3|3|M|Black||17|No|Mother|28206|7|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|M|White||29|28202|Bachelors Degree|Single|Business: Engineer|28202|5|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503635703|500187462|31|0|1|503979778|1|0|1|500777350|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||16705|3|||1|500014681|7960300212314874874|0
M191|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2372|Red|Amachi|2010-03-10|2010-03-23|2016-09-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||77.9||2|2|1|1|M|Multi-race (Black & Hispanic)||17|Yes|Mother|28208|9|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Hispanic||28|28277|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501340097|501340376|38|0|1|501934966|3|0|1|500440292|10|2|500003586||4|3|500000294|-2||-2|0|10|||7464|9|||1|500000294|0|0
M192|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1789|Green|Project Big|2012-04-05|2012-04-13|NaT||||58.8||1|1|1|1|M|Black||17|No|GrandMother|28208|11|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community|Project Big|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502710796|502711683|31|0|1|502926804|1|0|1|500608316|10|2|500004641||2|1|500004640|-2||-2|6854|8|||7464|9|||1|500004640|2611337051335117774|0
M193|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|231|Yellow|mentor2.0 2015|2015-10-25|2015-11-17|2016-07-05|Child: Changed school/site|Child: Changed school/site||7.6||1|1|3|3|M|Black||17|No|Mother|28217|9|Two Parent|Unknown||||Yes||Relative|General Site|mentor2.0 2015|Match Support|M|Black||49|28027|Bachelors Degree|Married|Transport: Driver|28208|6|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|0|1|1|0|277|60|598|500000170|500017786|504426368|504428623|31|0|1|500863980|31|0|1|500851862|10|1|500014504||4|2|500015184|-1|500014505, 500014506|-1|0|3|||7671|13|||1|500015184|702163000107564368|0
M194|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|662|Red||2014-04-07|2014-05-31|2016-03-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.7||2|2|1|1|M|Black||17|Yes|Mother|28205|9|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community|Amachi|Match Support|M|White||29|28210|Bachelors Degree|Single|Finance||2|4|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500764138|500764404|31|0|1|503707921|1|0|1|500758491|10|2|-2||4|3|500000294|-2|500000294|-2|0|10|||7464|9|||1||7501346876523517480|0
M195|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|348|Green||2014-10-07|2014-10-08|2015-09-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||11.4||1|1|2|2|F|Black||17|No|Mother|28217||One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||34|28216|Masters Degree|Single|Business|28202|8|7|Self|Self|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043114|504045132|31|0|2|502261758|31|0|2|500781139|10|1|500014504||4|1||-1|500014505, 500014506|-1|0|4|||7464|9|||1||702163000107564368|0
M196|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|343|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|2016-10-14|Child: Lost interest|Child: Lost interest||11.3||1|1|1|1|M|Black||17|No|Mother|28216|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||36|28210||Married|Consultant|28211|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|0|1|1|0|277|60|598|500000170|500021786|504447778|504450034|31|0|1|504350981|1|0|1|500846247|10|1|500014504||4|1||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M197|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1809|Green|2010-2012 OJJDP JJI|2011-08-16|2011-08-29|2016-08-11|Child: Lost interest|Child: Lost interest||59.4||1|1|2|2|M|Black||17|No|Mother|28078|9|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|502097843|502098263|31|0|1|502643791|3|0|1|500550390|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|500005291|3455806768141331471|0
M198|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|882|Green|mentor2.0, mentor2.0 2014|2014-10-07|2014-10-07|NaT||||29||1|1|1|1|M|Black||17|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2014|Match Support|M|White||40|28205|Masters Degree|Married|Consultant|28202|0|4|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504043467|504045485|31|0|1|503971844|1|0|1|500781241|10|1|500014504||2|1|500014505, 500014506|-1|500014505, 500014506|-1|0|4|||7462|13|||1|500014505, 500014506|702163000107564368|0
M199|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|987|Green||2014-06-18|2014-06-24|NaT||||32.4||3|3|1|1|M|Black||17|No|Relative: Other|28208|10|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||29|28205||Single|Consultant|2210|2|10|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500340183|500340317|31|0|1|503868914|1|0|1|500766977|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1||0|0
M200|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|540|Yellow||2013-08-05|2013-08-20|2015-02-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.7||1|1|2|2|M|Black||17|No|Mother|28262|8|One Parent: Female|$25,000 to $29,999||||Yes||Relative|General Community||Match Support|M|Black||34|28213|Bachelors Degree|Single|Finance: Banking|28202|0|2|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503443162|503445028|31|0|1|500234684|31|0|1|500705816|10|2|-2||4|2||-2||-2|0|3|||7458|9|||1||1320477920662455183|7891205870025752229
M201|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1065|Red||2012-04-01|2012-04-30|2015-03-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||35||1|1|1|1|F|Multi-Race (None of the above)||17|No|Father|28214|6|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|White||33|28216|Bachelors Degree|Single|Business: Sales|28270|2|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502828131|502829415|7|0|2|502881454|1|0|2|500607446|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||6095563712459522926|0
M202|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2289|Green||2010-11-22|2010-11-30|NaT||||75.2||3|3|2|2|F|Black||17|No|Mother|28209||One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|F|White||39|28210|Masters Degree|Single|Education|28212|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|1|0|0|1|277|60|598|500000170|500020910|500829028|502254499|31|0|2|501978180|1|0|2|500498594|10|2|-2||2|1||-2|500000294, 500004640|-2|0|10|||7464|9|||1||7872663507285703533|0
M203|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1175|Green||2013-12-05|2013-12-18|NaT||||38.6||1|1|1|1|F|Black||17|No|Mother|28212|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||26|11237||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020753|502868969|502870370|31|0|2|503574667|1|0|2|500736904|10|2|-2||2|1||-2|500000294|-2|0|10|||46|2|||1||6381341368426079638|7044657180546140448
M204|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1840|Green||2012-01-27|2012-02-22|NaT||||60.5||1|1|1|1|M|Black||17|No|Mother|28269|5|One Parent: Female|$15,000 to $19,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||34|28269|Bachelors Degree|Single|Business: Human Resources|28025|2|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502469903|502470350|31|0|1|502868874|31|0|1|500594396|10|2|-2||2|1||-2||-2|0|5|||4748|14|1360|3|1||0|6147479637696055847
M205|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|883|Green|mentor2.0, mentor2.0 2014|2014-10-06|2014-10-06|NaT||||29||1|1|1|1|F|Black||17|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|F|Black||38|28216|Masters Degree|Married|Business|28255|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site||Match Support|1|0|0|1|277|60|598|500000170|500022907|504043252|504045270|31|0|2|503974167|31|0|2|500780750|10|1|500014504||2|1||-1||-1|0|3|||7462|13|||1|500014505, 500014506|702163000107564368|0
M206|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|232|Green|PERL 2014-2016|2014-10-27|2014-12-02|2015-07-22|Child: Changed school/site|Child: Changed school/site||7.6||1|1|1|1|F|Black||17|No|GrandMother|28208|8|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|Black||23|28262|High School Graduate|Single|Student: College|28278|0|0|Self|Self|Big|General Site|PERL 2014-2016|Enrollment|1|0|1|0|277|60|598|500000170|500016270|504059403|504061427|31|0|2|503658554|31|0|2|500788554|10|1|500000295|2128173561|4|1|500014681|-1|500014681|-1|0|4|||7464|9|||1|500014681|7960300212314874874|0
M207|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|913|Green||2014-08-21|2014-08-30|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||30||1|1|1|1|M|Black||17|No|Mother|28215|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|M|Black||38|28269||Single|Unemployed||0|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503813942|503815919|31|0|1|503873603|31|0|1|500773055|10|2|-2||4|1||-2||-2|0|3|||17101|1|||1||3148273126074974335|0
M208|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|752|Green|mentor2.0, mentor2.0 2014|2014-10-07|2014-10-07|2016-10-28|Child: Changed school/site|Child: Changed school/site||24.7||1|1|1|1|F|Hispanic||17|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2014|Match Support|F|White||28|28209|Masters Degree|Single|Finance: Accountant|28223|0|7|Self|Self|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504043100|504045118|3|0|2|503962672|1|0|2|500781120|10|1|500014504||4|1|500014505, 500014506|-1|500014506|-1|0|4|||7464|9|||1|500014505, 500014506|702163000107564368|0
M209|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|112|Green||2014-10-08|2014-10-16|2015-02-05|Child/Family: Moved|Child/Family: Moved||3.7||1|1|2|2|M|Black||17|Yes|Father|28208|9|One Parent: Male|Unknown||||No||School|General Site||Match Support|M|White||51|28277|Bachelors Degree|Married|Finance|28277|0|0|Igniting Breakfast|Special Event|Big|General Community|mentor2.0, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043445|504045463|31|0|1|503922166|1|0|1|500781673|10|1|-1||4|1||-1|500014505, 500014506|-2|0|4|||17266|8|||1||702163000107564368|0
M210|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1992|Green|Project Big, 2010-2012 OJJDP JJI|2011-08-29|2011-09-11|2017-02-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||65.4||1|1|1|1|M|Black||17|No|Mother|28208|5|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||51|28207|Masters Degree|Married|Business|28202|0|7|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020910|502602958|501480402|31|0|1|502578040|1|0|1|500552390|10|2|500004641||4|1|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291|5493246288421413675|0
M211|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|757|Green||2015-01-22|2015-02-09|NaT||||24.9||1|1|1|1|F|Black||17|No|Mother|28217|8|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Black||24|28273|Some College|Single|Finance: Accountant|28226|6|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|504169896|504172004|31|0|2|503987952|31|0|2|500809606|10|2|-2||2|1|500014681|-2||-2|0|4|||46|2|||1||7458247995093008174|0
M212|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3126|Green||2008-07-23|2008-08-15|NaT||||102.7||1|1|1|1|M|Black||17|No|Mother|28269|10|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Asian||35|28210|Bachelors Degree|Married|Business: Sales|28217|5|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501195410|501195684|31|0|1|501277677|4|0|1|500278978|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||0|8858586900346693884
M213|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|332|Green||2014-11-17|2014-11-24|2015-10-22|Child/Family: Moved|Child/Family: Moved||10.9||1|1|1|1|F|Black||17|No|Mother|28269|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||39|28078|Bachelors Degree|Single|Business: Sales|28117|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503873575|503875571|31|0|2|504004351|1|0|2|500796129|10|2|-2||4|1||-2||-2|0|10|||46|2|||1||932861092942387634|7044657180546140448
M214|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|876|Green||2014-10-07|2014-10-13|NaT||||28.8||1|1|1|1|M|Black||16|No|Mother|28213|8|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|Black||48|28262||Single|Retired||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503923102|503925109|31|0|1|503996589|31|0|1|500781196|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||3677730851176818072|1060411471255530133
M215|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0, mentor2.0 2015|2015-10-23|2015-11-17|NaT||||15.6||1|1|1|1|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||33|28078|Masters Degree|Married|Business: Human Resources|28078|7|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504426028|504428283|31|0|2|504357594|1|0|2|500851407|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||17159|12|||1|500014505, 500015184|702163000107564368|0
M216|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|421|Green||2014-08-12|2014-08-25|2015-10-20|Volunteer: Time constraint|Volunteer: Time constraint||13.8||1|1|1|1|F|Black||16|No|Mother|28227|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||30|28273|Bachelors Degree|Single|Business: Human Resources|28203|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503796616|503798593|31|0|2|503828896|1|0|2|500772098|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||0|7044657180546140448
M217|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1137|Green|Cabarrus County|2013-12-12|2014-01-25|NaT||||37.4||2|2|1|1|F|Black||16|No|Mother|28083|11|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||41|28027|Bachelors Degree|Married|Human Services|28025|0|9|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502761850|502762654|31|0|2|503632186|31|0|2|500738602|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|1557072896577419067|4058276550489173605
M218|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|245|Green||2014-10-07|2014-10-07|2015-06-09|Child: Lost interest|Child: Lost interest||8||3|3|1|1|M|Black||16|No|Aunt|28208|9|Other Relative|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||27|28216|Bachelors Degree|Living w/ Significant Other|Finance: Accountant|28202|0|11|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500016847|503216855|503218636|31|0|1|503969586|31|0|1|500781240|10|1|500014504||4|1||-1|500014506|-1|0|4|||7462|13|||1||702163000107564368|0
M219|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|374|Yellow||2014-01-14|2014-01-27|2015-02-05|Volunteer: Time constraint|Volunteer: Time constraint||12.3||1|1|3|3|M|Black||16|No|Mother|28215|8|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||26|28203|Bachelors Degree|Single|Finance: Banking|28213|0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503587930|503589807|31|0|1|500942257|1|0|1|500742670|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||0|2466453775578950862
M220|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2025|Green||2010-01-21|2010-01-26|2015-08-13|Child: Lost interest|Child: Lost interest||66.5||2|2|2|2|F|Black||16||GrandMother|28215|3|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||41|28277|Bachelors Degree|Single|Business: Mgt, Admin||9|0|General|Other Big|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500017732|501735420|501735760|31|0|2|500956022|1|0|2|500428818|10|2|-2||4|1||-2||-2|6854|8|||6450|12|||1||0|904091744937704216
M221|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2685|Green||2009-10-19|2009-10-30|NaT||||88.2||2|2|1|1|M|Black||16||Mother|28216|9|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28078|||Medical: Pharmacist|28210|10|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|500713817|500714084|31|0|1|501834795|1|0|1|500396466|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1||7301546317881317703|8947522103573893278
M222|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3094|Green||2008-09-11|2008-09-16|NaT||||101.7||1|1|1|1|F|Black||16|No|Mother|28216|8|Grandparents|Unknown||||No|TV|Media|General Community||Match Support|F|Black||42|28212|Bachelors Degree|Single|Unknown|28202|8|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501234606|501234882|31|0|2|501233675|31|0|2|500287478|10|2|-2||2|1||-2||-2|56|1|||7464|9|||1||7284449467126735125|0
M223|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1988|Green|Amachi|2011-09-21|2011-09-27|NaT||||65.3||2|2|1|1|F|Black||16|Yes|GrandMother|28213|12|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||24|28027|Some College|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|502221847|502222278|31|0|2|502654877|31|0|2|500556560|10|2|500003586||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294|932861092942387634|0
M224|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|244|Red||2014-08-13|2014-08-29|2015-04-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||8||2|2|1|1|F|Black||16|No|Mother|28269|8|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||34|28269|Masters Degree|Single|Medical|28025|1|7|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|502551045|502551498|31|0|2|503859553|1|0|2|500772207|10|2|-2||4|3||-2||-2|0|4|||17159|12|||1||3677730851176818072|0
M225|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|358|Green|mentor2.0 2015|2015-10-25|2015-11-05|2016-10-28|Child: Changed school/site|Child: Changed school/site||11.8||1|1|2|2|F|Black||16|Yes|Mother|28208|9|One Parent: Female|Unknown||||Yes||Relative|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||25|28203|Bachelors Degree|Single|Business|28201|1|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015, mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500017786|504454510|504456768|31|0|2|504357339|1|0|2|500851879|10|1|500014504||4|1|500014505, 500015184|-1|500014505, 500015184, 500016394|-1|0|3|||7462|13|||1|500015184|702163000107564368|0
M226|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|1220|Green||2012-02-01|2012-02-13|2015-06-17|Child: Changed school/site|Child: Changed school/site||40.1||1|1|1|1|F|Black||16|Yes|Mother|28205|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||49|28208|High School Graduate|Single|Business: Mgt, Admin||9|0|Recruitment Event|BBBS Board/Staff|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|502763473|502764385|31|0|2|502828246|31|0|2|500595333|10|1|500000295|2128173561|4|1||-1||-1|0|4|||7462|13|||1||7960300212314874874|0
M227|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|395|Green||2014-10-07|2014-10-07|2015-11-06|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||13||1|1|1|1|M|Hispanic||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||33|28207|Masters Degree|Single|Business||0|3|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504050643|504052667|3|0|1|503969686|1|0|1|500781223|10|1|500014504||4|1||-1|500014505, 500014506|-1|0|4|||7462|13|||1||702163000107564368|0
M228|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|371|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-10-26|2016-10-31|Child: Changed school/site|Child: Changed school/site||12.2||1|1|1|1|F|Black||16|No|Father|28217|9|One Parent: Male|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||46|28036|Bachelors Degree|Married|Business|28078|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504426151|504428406|31|0|2|504431643|1|0|2|500851863|10|1|500014504||4|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M229|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|756|Green|mentor2.0 2014|2014-10-06|2014-10-06|2016-10-31|Child: Changed school/site|Child: Changed school/site||24.8||1|1|1|1|F|Black||16|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||25|28202|Bachelors Degree|Single|Business|28202|1|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504043352|504045370|31|0|2|503969666|31|0|2|500780891|10|1|500014504||4|1||-1|500014506|-1|0|4|||7462|13|||1|500014506|702163000107564368|0
M230|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1710|Red|2010-2012 OJJDP JJI|2011-02-17|2011-02-28|2015-11-04|Volunteer: Moved|Volunteer: Moved||56.2||1|1|1|1|F|Black||16|No|Mother|28208|10|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28205|Masters Degree|Single|Medical: Doctor, Provider|28277|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501833031|501833394|31|0|2|502427342|1|0|2|500518294|10|2|-2||4|3|500005291|-2||-2|0|10|||7464|9|||1|500005291|702163000107564368|0
M231|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1924|Green||2011-10-28|2011-11-30|NaT||||63.2||1|1|1|1|F|Black||16||GrandMother|28269|8|Grandparents|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28269|Masters Degree|Single|Finance: Banking|28255|15|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502580335|502580838|31|0|2|502677590|31|0|2|500571804|10|2|-2||2|1|500005291|-2||-2|0|10|||7464|9|||1||0|0
M232|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|893|Green|PERL 2014-2016|2014-09-04|2014-09-19|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29.3||1|1|1|1|M|Black||16|No|Mother|28208|8|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||39|28262|Bachelors Degree|Single|Finance|28262|3|2|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500020752|503524036|503525911|31|0|1|503913408|31|0|1|500774440|10|2|-2||4|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681|7581500809034284566|3402014428779854546
M233|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|333|Green|mentor2.0 2015|2015-10-25|2015-11-30|2016-10-28|Child/Family: Moved|Child/Family: Moved||10.9||1|1|3|3|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|White||40|28078|Bachelors Degree|Single|Human Services: Social Worker|28277|0|9|Relative|Relative|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504454500|504456758|31|0|2|503529603|1|0|2|500851877|10|1|500014504||4|1|500015184|-1|500014505, 500015184|-1|0|4|||17161|11|||1|500015184|702163000107564368|0
M234|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|988|Green||2014-06-10|2014-06-23|NaT||||32.5||1|1|1|1|F|Black||16|No|Mother|28227|9|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||30|28205|Bachelors Degree|Single|Business|28262|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503767186|503769162|31|0|2|503788125|31|0|2|500766047|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||3292090474897428830|0
M235|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|830|Red|PERL 2014-2016|2014-11-12|2014-11-21|2017-02-28|Child/Family: Time constraints|Child/Family: Time constraints||27.3||1|1|1|1|F|Black||16|No|GrandMother|28269|9|One Parent: Female|Unknown|||Y|Yes||Foster Home|General Community|PERL 2014-2016|Match Support|F|Black||24|28217|Bachelors Degree|Single|Finance||0|2|AA Task Force|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500008321|504085882|503144847|31|0|2|503977000|31|0|2|500794719|10|2|-2||4|3|500014681|-2|500014681|-2|0|7|||9229|13|||1|500014681|4565518866290635873|8233867082779775199
M236|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|1072|Green|mentor2.0, mentor2.0 2015|2013-11-07|2013-11-07|2016-10-14|Volunteer: Time constraint|Volunteer: Time constraint||35.2||3|3|1|1|M|Black||16|No|Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||School|General Site|mentor2.0 2016|Match Support|M|Black||43|28216|Some College|Divorced|Consultant|28217|4|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500021786|503236129|503237920|31|0|1|503682677|31|0|1|500728645|10|1|500014504||4|1|500016394|-1||-1|0|4|||11247|3|||1|500014505, 500015184|3935539763241716148|0
M237|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green|mentor2.0 2016|2016-11-18|2016-11-18|NaT||||3.6||3|3|2|2|M|Black||16|No|Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||School|General Site|mentor2.0 2016|Match Support|M|White||30|28207||Single|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500021786|503236129|503237920|31|0|1|504434419|1|0|1|500929505|10|1|500014504||2|1|500016394|-1|500015184, 500016394|-1|0|4|||7462|13|||1|500016394|3935539763241716148|0
M238|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|1464|Green||2012-10-25|2012-10-25|2016-10-28|Child: Changed school/site|Child: Changed school/site||48.1||1|1|1|1|M|Black||16|No|Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Black||42|28269|Bachelors Degree|Married|Finance|28217|5|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|503236165|503237920|31|0|1|503163281|31|0|1|500651688|10|1|500014504||4|1|500014505, 500015184|-1||-1|0|4|||11247|3|1204|3|1||3935539763241716148|0
M239|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|965|Green||2014-06-27|2014-07-16|NaT||||31.7||3|3|1|1|F|Black||16|Yes|Mother|28206|10|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|Black||28|28223|Masters Degree|Single|Student: College|28223|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|501096791|501097065|31|0|2|503803014|31|0|2|500768008|10|2|-2||2|1||-2||-2|0|4|||46|2|||1||6286214584598985826|7044657180546140448
M240|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|756|Green|mentor2.0, mentor2.0 2014|2014-10-06|2014-10-06|2016-10-31|Child: Severity of challenges|Child: Severity of challenges||24.8||1|1|1|1|F|Native Hawaiian or Other Pacific Islander||16|No|Mother|28217||One Parent: Female|Unknown|||Y|Yes||Relative|General Site|mentor2.0, mentor2.0 2014|Match Support|F|White||24|28203|Bachelors Degree|Single|Finance: Banking||0|6|Self|Self|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504043184|504045202|5|0|2|504024311|1|0|2|500780788|10|1|500014504||4|1|500014505, 500014506|-1|500014505, 500014506|-1|0|3|||7464|9|||1|500014505, 500014506|702163000107564368|0
M241|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|883|Green|mentor2.0, mentor2.0 2014|2014-10-06|2014-10-06|NaT||||29||1|1|1|1|F|Black||16|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2014|Match Support|F|White||27|28210|Masters Degree|Married|Customer Service|28209|0|1|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504043120|504045138|31|0|2|503974816|1|0|2|500780896|10|1|500014504||2|1|500014505, 500014506|-1|500014506|-1|0|4|||17159|12|||1|500014505, 500014506|702163000107564368|0
M242|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1296|Green||2013-01-10|2013-01-30|2016-08-18|Child/Family: Moved|Child/Family: Moved||42.6||2|2|1|1|M|Black||16|No|Aunt|28213|8|One Parent: Female|$40,000 to $44,999||||Yes||School|General Community|Project Big|Match Support|M|White||33|28209|Associate Degree|Married|Business: Mgt, Admin||0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|502555551|502556004|31|0|1|503207140|1|0|1|500674218|10|2|-2||4|1|500004640|-2||-2|0|4|||7464|9|||1||5441374193599827162|0
M243|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|570|Green||2013-10-14|2013-11-25|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||18.7||1|1|1|1|M|Black||16|No|Mother|28206|7|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||33|28226|Bachelors Degree|Married|Business|28202|8|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503578835|503580712|31|0|1|503605630|1|0|1|500718994|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|7044657180546140448
M244|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3645|Green||2007-03-08|2007-03-15|NaT||||119.8||1|1|1|1|F|Black||16|No|Mother|28269|9|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||Match Support|F|White||34|28210|Bachelors Degree|Single|Education: Teacher|28226|0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|500824037|500824306|31|0|2|500789337|1|0|2|500165956|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||3960869250587139051|0
M245|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green|mentor2.0 2016|2016-11-18|2016-11-18|NaT||||3.6||1|1|2|2|F|Black||16|No|Mother|28217|11|Two Parent|$10,000 to $14,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||29|28216|Masters Degree|Single|Medical|30005|0|5|BBBS National Site|Web Link|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500022907|504842862|504845364|31|0|2|504300098|31|0|2|500929477|10|1|500014504||2|1|500014505, 500016394|-1|500015184|-1|0|4|||46|2|||1|500016394|702163000107564368|0
M246|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|753|Green|mentor2.0 2014|2014-10-06|2014-10-06|2016-10-28|Child: Changed school/site|Child: Changed school/site||24.7||1|1|1|1|F|Black||16|No|Mother|28208||One Parent: Female|Unknown|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||37|28203|Masters Degree|Divorced|Business|28202|10|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504043105|504045123|31|0|2|503969642|1|0|2|500780806|10|1|500014504||4|1|500014505, 500015184|-1|500014506|-1|0|4|||7462|13|||1|500014506|702163000107564368|0
M247|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-09-23|2015-10-26|NaT||||16.4||1|1|2|2|F|Black||16|No|Mother|28208|9|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||26|28205|Bachelors Degree|Single|Business|28255|1|3|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500022907|504180420|504182529|31|0|2|504001561|31|0|2|500841752|10|1|500014504||2|1|500014505, 500015184|-1|500014506|-1|34|2|||7671|13|||1|500014505, 500015184|6353565629814722343|8858586900346693884
M248|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|879|Yellow||2013-02-13|2013-02-28|2015-07-27|Child: Lost interest|Child: Lost interest||28.9||1|1|1|1|F|Black||16|No|GrandMother|28212|9|One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||46|28262|PHD|Single|Education: College Professor|28223|5|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|502581328|502581832|31|0|2|503144090|31|0|2|500681651|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1||1010189231295710785|645589252192201558
M249|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2115|Yellow||2010-10-11|2010-10-21|2016-08-05|Volunteer: Time constraint|Volunteer: Time constraint||69.5||1|1|1|1|M|White||16|No|Mother|28213|4|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community||Match Support|M|White||37|28205||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502063945|502064367|1|0|1|502295138|1|0|1|500478943|10|2|500004641||4|2||-2||-2|0|5|||7496|10|||1||0|0
M250|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2038|Yellow|Project Big|2010-10-20|2010-10-27|2016-05-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||67||1|1|1|1|F|Black||16||Mother|28212|5|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|F|White||33|28227|Bachelors Degree|Single|Unknown||9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|1|0|1|0|277|60|598|500000170|500008321|502338225|502338658|31|0|2|502312449|1|0|2|500483095|10|2|500004641||4|2|500004640|-2|500004640|-2|0|4|||7496|10|||1|500004640|7869308672550505300|0
M251|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1748|Green|Amachi|2012-05-15|2012-05-24|NaT||||57.4||2|3|1|1|M|Black||16|Yes|Mother|28216|9|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Match Support|M|White||34|28203|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500186245|500187840|31|0|1|502989318|1|0|1|500614903|10|2|500003586||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294|253338316288302752|1818964647027278255
M252|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1482|Green|Cabarrus County|2013-01-25|2013-02-14|NaT||||48.7||2|2|1|1|M|White||16|Yes|GrandMother|28083|9|Grandparents|Unknown|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||51|28117|Masters Degree|Divorced|Consultant|28117|12|11|Local Print|Media|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|501227649|501227925|1|0|1|503316978|1|0|1|500677437|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|10|||7439|1|||1|500016374|1557072896577419067|0
M253|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|121|Green||2014-10-07|2014-10-07|2015-02-05|Child/Family: Moved|Child/Family: Moved||4||1|1|3|3|M|Black||16|No|Father|28217|9|One Parent: Male|Unknown|||Y|Yes||School|General Site||Enrollment|M|Black||32|28216|Masters Degree|Single|Finance: Accountant|28280|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014, mentor2.0 2016|Match Support|1|0|1|0|277|60|598|500000170|500016847|504050627|504052651|31|0|1|503976447|31|0|1|500781229|5|1|-1||4|1||-1|500014505, 500014506, 500016394|-1|0|4|||7462|13|||1||702163000107564368|0
M254|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|333|Green|mentor2.0 2015|2015-10-23|2015-11-30|2016-10-28|Child: Lost interest|Child: Lost interest||10.9||1|1|3|3|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Black||31|28203|Juris Doctorate (JD)||Law: Lawyer|28203|1|0|Self|Self|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504445059|504447315|31|0|1|501631588|31|0|1|500851408|10|1|500014504||4|1|500014505, 500015184|-1|500015184|-1|0|4|||7464|9|||1|500015184|702163000107564368|0
M255|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3409|Yellow||2007-04-30|2007-04-30|2016-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||112||1|1|1|1|M|Black||16||Mother|28206|8|Two Parent|Less than $10,000|||Y|No||Self|General Community||Match Support|M|White||36|28203|||Retail: Sales|28226|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|500783100|500783368|31|0|1|500777047|1|0|1|500174449|10|2|-2||4|2||-2||-2|0|10|||46|2|||1||4863631750424600365|0
M256|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|754|Green||2013-03-11|2013-03-13|2015-04-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.8||1|1|1|1|M|Black||16|Yes|Mother|28273|8|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||43|29707|Bachelors Degree|Separated|Govt||10|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503296945|503298770|31|0|1|503381327|31|0|1|500687021|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||932861092942387634|880099004922011679
M257|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1916|Green||2011-11-18|2011-12-08|NaT||||62.9||1|1|1|1|F|Black||16|No|Mother|28205|7|One Parent: Female|$25,000 to $29,999|||Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||29|28120|Bachelors Degree|Single|Govt: Clerical||0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500021785|502760967|502761879|31|0|2|502666332|31|0|2|500579826|10|2|-2||2|1|500005291|-2||-2|2203|12|||7464|9|||1||8758769076374727509|0
M258|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|349|Green||2014-10-07|2014-10-07|2015-09-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||11.5||1|1|2|2|F|Black||16|Yes|Mother|28208|9|One Parent: Female|Less than $10,000|||Y|No||Self|General Site||Match Support|F|Black||37|28269|Masters Degree|Single|Human Services: Social Worker|28212|0|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|1|0|1|0|277|60|598|500000170|500016847|500905037|500905305|31|0|2|501564519|31|0|2|500781149|10|1|500014504||4|1||-1|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||702163000107564368|0
M259|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|752|Green|mentor2.0, mentor2.0 2014|2014-10-07|2014-10-07|2016-10-28|Child/Family: Moved|Child/Family: Moved||24.7||1|1|1|1|F|Black||16|No|Mother|28269|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2014|Match Support|F|White||26|28209|Bachelors Degree|Single|Finance: Accountant|28202|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504050561|504052585|31|0|2|503971898|1|0|2|500781118|10|1|500014504||4|1|500014505, 500014506|-1|500014506|-1|0|4|||7462|13|||1|500014505, 500014506|702163000107564368|0
M260|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2451|Green||2009-06-02|2009-06-17|2016-03-03|Volunteer: Moved|Volunteer: Moved||80.5||1|1|1|1|M|Black||16|No|Mother|28216|8|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Service: Hotel|28202|2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501631140|501631463|31|0|1|501628976|1|0|1|500367187|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||0|0
M261|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|775|Red||2013-05-13|2013-06-13|2015-07-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||25.5||1|1|1|1|F|Black||16|No|Mother|28262|7|One Parent: Female|$15,000 to $19,999|Yes: Active|Yes|Y|Yes|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||37|28269|Masters Degree|Single|Business: Human Resources|28262|1|3|Recruitment Event|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503149009|503150686|31|0|2|503199095|31|0|2|500696674|10|2|-2||4|3||-2||-2|6855|8|||7460|12|||1||3677730851176818072|8392423513746229127
M262|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1768|Yellow||2012-04-24|2012-05-04|NaT||||58.1||2|2|1|1|F|Black||16|No|Mother|28216|9|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community||Match Support|F|Asian||32|28216|Bachelors Degree|Single|Business: Mgt, Admin|28208|0|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500740296|500740560|31|0|2|502893901|4|0|2|500611525|10|2|-2||2|2||-2||-2|0|5|||7464|9|||1||253338316288302752|0
M263|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2414|Yellow|Project Big|2010-07-28|2010-07-28|NaT||||79.3||1|1|2|2|F|Black||16|No|GrandMother|28208|5|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community|Project Big|Match Support|F|Black||37|28216|Bachelors Degree|Single|Customer Service||8|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|0|1|277|60|598|500000170|500008321|502234504|502234935|31|0|2|502129464|31|0|2|500463451|10|2|500004641||2|2|500004640|-2||-1|0|4|||11247|3|1204|3|1|500004640|6458351142431041105|3402014428779854546
M264|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|122|Green||2014-10-06|2014-10-06|2015-02-05|Child/Family: Moved|Child/Family: Moved||4||1|1|2|2|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||26|28205|Bachelors Degree|Single|Business|28255|1|3|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043501|504045519|31|0|2|504001561|31|0|2|500780922|10|1|-1||4|1||-1|500014506|-1|0|4|||7671|13|||1||702163000107564368|0
M265|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|123|Yellow|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|2016-03-08|Child: Changed school/site|Child: Changed school/site||4||1|1|2|2|M|Black||16|Yes|Father|28217|10|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|M|Black||40|28104|Masters Degree|Divorced|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500016847|504454641|504456899|31|0|1|500800975|31|0|1|500846225|10|1|500014504||4|2||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M266|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|138|Green|mentor2.0 2015|2015-10-25|2015-11-11|2016-03-28|Child: Family structure changed|Child: Family structure changed||4.5||1|1|2|2|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|Black||45|28217|Bachelors Degree|Divorced|Education: Teacher|28226|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504425996|504428251|31|0|2|504272278|31|0|2|500851874|10|1|500014504||4|1|500015184|-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M267|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|172|Green|mentor2.0, mentor2.0 2015|2016-02-09|2016-02-13|2016-08-03|Child/Family: Moved|Child/Family: Moved||5.7||1|1|1|1|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|White||27|28215|Bachelors Degree|Single|Business|28273|0|2|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|RTBM|0|1|1|0|277|60|598|500000170|500017786|504494261|504496546|31|0|1|504423999|1|0|1|500878530|10|1|500014504||4|1|500014505, 500015184|-1|500014505, 500016394|-1|0|4|||7464|9|||1|500014505, 500015184|702163000107564368|0
M268|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|634|Green||2013-10-28|2013-11-15|2015-08-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.8||1|1|2|3|F|Black||16|Yes|Mother|28213|7|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||29|28209|Bachelors Degree|Single|Finance|28202|5|0|Duke Energy|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500016270|503602174|503604051|31|0|2|503615576|1|0|2|500724064|10|1|500009132|2128173561|4|1||-1||-2|0|4|||16705|3|||1||7960300212314874874|0
M269|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1852|Red|Amachi|2010-07-12|2010-07-30|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||60.8||1|1|1|1|M|Black||16|Yes|Mother|28269|8|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28214|Some College|Married|Medical||3|6|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500015820|502171910|502172339|31|0|1|502141964|31|0|1|500460627|10|2|500003586||4|3|500000294|-2|500000294|-2|0|5|||7464|9|||1|500000294|9134125726462845918|1202530717971184330
M270|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1749|Green||2012-05-15|2012-05-23|NaT||||57.5||1|1|1|1|M|Black||16|No|Mother|28270|6|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|White||29|28203|Bachelors Degree||Finance: Accountant||1|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502866475|502867876|31|0|1|502961396|1|0|1|500614954|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||5994075768656267011|0
M271|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|114|Yellow|mentor2.0, mentor2.0 2015|2015-10-12|2015-11-06|2016-02-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.7||1|1|1|1|F|Black||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||42|28134|Masters Degree|Single|Finance: Auditor|28211|2|1|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2015|Enrollment|0|1|1|0|277|60|598|500000170|500016847|504447927|504450183|31|0|2|503868542|31|0|2|500846710|10|1|500014504||4|2||-1|500014505, 500015184|-1|0|4|||17159|12|||1|500014505, 500015184|702163000107564368|0
M272|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|321|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|2016-09-22|Volunteer: Time constraint|Volunteer: Time constraint||10.5||2|2|2|2|F|Black||16|No|Mother|28208||One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||48|28079||Married|Finance|28255|4|2|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|0|1|1|0|277|60|598|500000170|500021786|504447891|504450147|31|0|2|503984584|31|0|2|500846223|10|1|500014504||4|1|500014505, 500015184|-1|500014506|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M273|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|48|Green||2016-10-11|2017-01-18|NaT||||1.6||2|2|1|1|F|Black||16|No|Mother|28208||One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||25|28262|Bachelors Degree|Single|Business||0|2|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500021786|504447891|504450147|31|0|2|504739188|31|0|2|500914300|10|1|500014504||2|1|500014505, 500015184|-1|500014505, 500016394|-1|0|4|||17159|12|||1||702163000107564368|0
M274|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|841|Green|PERL 2014-2016|2014-11-03|2014-11-17|NaT||||27.6||1|1|1|1|M|Black||16|Yes|GrandMother|28270|9|One Parent: Female|$15,000 to $19,999|||Y|No||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||48|28226|Juris Doctorate (JD)|Married|Law: Lawyer|28202|4|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020910|503983132|503985143|31|0|1|503995895|1|0|1|500791249|10|2|-2||2|1|500014681|-2|500014681|-2|0|5|||46|2|||1|500014681|1010189231295710785|0
M275|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2016|2015-10-09|2015-11-06|NaT||||16||1|1|1|1|M|Hispanic||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||57|29941|Bachelors Degree|Married|Self-Employed, Entrepreneur|28031|30|0|Igniting Breakfast|Special Event|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504440300|504442556|3|0|1|504313945|1|0|1|500846204|10|1|500014504||2|1||-1|500015184|-1|0|4|||17266|8|||1|500014505, 500016394|702163000107564368|0
M276|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|879|Green||2013-11-15|2013-12-06|2016-05-03|Volunteer: Moved|Volunteer: Moved||28.9||1|1|1|1|F|Black||16|No|Mother|28262|9|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Retail: Sales|28217|0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503597088|503598965|31|0|2|503642924|1|0|2|500731612|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||7432163260389731024|1198499568025045356
M277|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2140|Green|2010-2012 OJJDP JJI|2011-04-23|2011-04-28|NaT||||70.3||1|1|1|1|M|White||16|No|Mother|28277|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||54|28205|Some College|Separated|Self-Employed, Entrepreneur|28214|29|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|502478428|502478875|1|0|1|502555822|1|0|1|500533009|10|2|-2||2|1|500005291|-2||-2|0|10|||7464|9|||1|500005291|3966805366522644621|0
M278|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|611|Green||2013-09-03|2013-09-25|2015-05-29|Volunteer: Moved|Volunteer: Moved||20.1||1|1|1|1|M|Black||16|No|Mother|28273|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||28|28207|Bachelors Degree|Single|Education: Teacher||1|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503496889|503498757|31|0|1|503490051|1|0|1|500708903|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||194235582162093094|6507622620494997521
M279|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2741|Green|Amachi|2009-08-19|2009-09-04|NaT||||90.1||1|1|1|1|F|Black||16|Yes|Mother|28262|9|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||40|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28204|0|9|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501597228|501597548|31|0|2|501397328|31|0|2|500379964|10|2|500003586||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294|2374609189072499123|6168060654679577655
M280|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1058|Red||2012-03-30|2012-04-30|2015-03-24|Volunteer: Time constraint|Volunteer: Time constraint||34.8||1|1|1|1|M|Black||16|No|Mother|28214|6|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Bachelors Degree|Single|Finance|28216|3|0|Relative|Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502319984|502320419|31|0|1|502290677|1|0|1|500607367|10|2|-2||4|3|500005291|-2||-2|6854|8|||17161|11|||1||806697982905023857|3482130045776789614
M281|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|336|Green|mentor2.0 2015|2015-10-25|2015-11-30|2016-10-31|Child: Changed school/site|Child: Changed school/site||11||1|1|1|1|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown|||Y|No||School|General Site|mentor2.0 2015|Match Support|F|White||27|28203|Masters Degree|Living w/ Significant Other|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504426057|504428312|31|0|2|504363902|1|0|2|500851869|10|1|500014504||4|1|500015184|-1|500014505, 500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M282|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0 2015|2015-10-23|2015-11-17|NaT||||15.6||3|3|3|3|F|Black||16|No|Mother|28208|9|One Parent: Female|$15,000 to $19,999||||No||School|General Site||Match Support|F|Black||36|28078|Masters Degree|Married|Business: Marketing|28273|1|1|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500021786|502537469|502537922|31|0|2|502056302|31|0|2|500851387|10|1|500014504||2|1||-1|500014505, 500014506|-1|0|4|||7671|13|||1|500015184|702163000107564368|0
M283|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|751|Green||2013-06-26|2013-07-17|2015-08-07|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||24.7||3|3|2|2|F|Black||16|No|Mother|28208|9|One Parent: Female|$15,000 to $19,999||||No||School|General Site||Match Support|F|White||34|28078|Masters Degree|Single|Medical: Doctor, Provider|28001|0|2|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500017732|502537469|502537922|31|0|2|503323641|1|0|2|500702088|10|2|-2||4|1||-1|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||702163000107564368|0
M284|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|463|Green|mentor2.0 2015|2015-10-25|2015-11-30|NaT||||15.2||1|1|1|1|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|White||25|28036|Bachelors Degree|Single|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504419900|504422153|31|0|2|504351222|1|0|2|500851861|10|1|500014504||2|1|500015184|-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M285|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1550|Yellow||2012-05-01|2012-05-08|2016-08-05|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||50.9||3|3|1|1|F|Black||16||Mother|28213|5|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||28|28211|Bachelors Degree|Single|Human Services||2|0|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501143674|501143948|31|0|2|502958999|1|0|2|500612879|10|2|500004641||4|2||-2||-2|0|10|||132|8|||1||6713311931049891381|0
M286|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|201|Green||2014-09-04|2014-09-19|2015-04-08|Volunteer: Moved|Volunteer: Moved||6.6||4|4|1|1|F|Black||16|No|Mother|28213|8|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||RTBM|F|Black||30|28269|Masters Degree|Single|Medical||0|11|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500011349|500826100|500801835|31|0|2|503877762|31|0|2|500774526|7|2|-2||4|1||-2|500000294|-2|0|10|||46|2|||1||9134125726462845918|0
M287|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2815|Green||2009-06-15|2009-06-22|NaT||||92.5||1|1|1|1|M|Black||16|No|Mother|28214|9|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|M|White||46|28277||Married|Business: Mgt, Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500910037|500910307|31|0|1|500856100|1|0|1|500368834|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||216500609169513656|0
M288|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3039|Green|Amachi|2008-01-31|2008-02-21|2016-06-17|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||99.8||2|2|1|1|F|Black||16|Yes|Mother|28217|10|One Parent: Female|$15,000 to $19,999|||Y|No|TV|Media|General Community|Amachi|Match Support|F|Black||32|28269|Bachelors Degree|Single|Business: Marketing|28273|0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500843863|500844129|31|0|2|501078655|31|0|2|500241388|10|2|500003586||4|1|500000294|-2|500000294|-2|56|1|||2238|7|||1|500000294|702163000107564368|0
M289|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|371|Green|mentor2.0 2015|2015-10-25|2015-10-26|2016-10-31|Volunteer: Moved|Volunteer: Moved||12.2||1|1|1|1|M|Hispanic||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|M|White||59|28205|Bachelors Degree|Married|Business: Marketing|28205|15|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0|Match Support|0|1|1|0|277|60|598|500000170|500017786|504445029|504447285|3|0|1|504272155|1|0|1|500851866|10|1|500014504||4|1|500015184|-1|500014505|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M290|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2714|Green||2008-08-13|2008-08-27|2016-02-01|Volunteer: Moved|Volunteer: Moved||89.2||1|1|1|1|F|Black||16|No|Mother|28211|10|Two Parent|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||37|28027|PHD|Single|Education: College Professor|27411|1|8|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|501288021|501288299|31|0|2|501249338|31|0|2|500281778|10|2|-2||4|1||-2||-2|0|10|||46|2|||1||7501346876523517480|0
M291|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3101|Green||2007-11-29|2007-12-20|2016-06-16|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||101.9||1|1|2|2|M|Black||16|No|Mother|28227||One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||40|28210|Bachelors Degree|Married|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|1|0|1|0|277|60|598|500000170|500017732|500936718|500915629|31|0|1|501027885|1|0|1|500224574|10|2|-2||4|1||-2|500014505, 500015184|-1|34|2|||46|2|||1||7960300212314874874|0
M292|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|364|Green||2014-10-06|2014-10-06|2015-10-05|Child/Family: Moved|Child/Family: Moved||12||1|1|2|2|F|Black||16|No|Father|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||38|28209|Bachelors Degree|Single|Business|28202|13|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043155|504045173|31|0|2|503985283|1|0|2|500780911|10|1|500014504||4|1||-1|500014506|-1|0|4|||7462|13|||1||702163000107564368|0
M293|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|725|Green|mentor2.0, mentor2.0 2014|2014-11-03|2014-11-03|2016-10-28|Child/Family: Time constraints|Child/Family: Time constraints||23.8||1|1|1|1|F|Black||16|No|Mother|28208|9|Two Parent|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2014|Match Support|F|Black||53|28079|Masters Degree|Married|Finance|28202|18|4|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504099617|504101651|31|0|2|503984599|31|0|2|500791106|10|1|500014504||4|1|500014505, 500014506|-1|500014506|-1|0|4|||7462|13|||1|500014505, 500014506|702163000107564368|0
M294|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2587|Yellow|Amachi|2009-08-24|2009-08-24|2016-09-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||85||1|1|1|1|M|Black||16|Yes|Mother|28213|10|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||51|28214|Masters Degree|Married|Business: Sales|94108|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501825910|500188141|31|0|1|501196986|1|0|1|500380446|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7496|10|||1|500000294|7432163260389731024|0
M295|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|NaT||||16||1|1|1|1|M|Black||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||60|28270||Married|Finance||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504447802|504450058|31|0|1|504350780|1|0|1|500846222|10|1|500014504||2|1||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M296|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1807|Green||2012-03-01|2012-03-26|NaT||||59.4||1|1|1|1|F|Black||16|No|Mother|28217|11|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Asian||35|28210|Masters Degree|Married|Arts, Entertainment, Sports|28202|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502610186|502610737|31|0|2|502913393|4|0|2|500601697|10|2|-2||2|1||-2||-2|6854|8|||7671|13|||1||702163000107564368|0
M297|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-11-17|NaT||||15.6||1|1|1|1|F|Hispanic||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||25|28202|Bachelors Degree|Single|Business|28202|2|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504426106|504428361|3|0|2|504355965|1|0|2|500851867|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M298|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|767|Green||2014-05-07|2014-05-15|2016-06-20|Child/Family: Moved|Child/Family: Moved||25.2||1|1|1|1|M|White||16||Mother|28277|8|One Parent: Female|$40,000 to $44,999|||Y|No||Self|General Community||Match Support|M|White||60|28105|Bachelors Degree|Married|Tech: Research/Design|28277|4|0|Recruitment Event|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|503187841|503189585|1|0|1|503789478|1|0|1|500762532|10|2|-2||4|1||-2||-2|0|10|||7460|12|||1||5994075768656267011|1990673839571477301
M299|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Inactive|Match Support|481|Green|mentor2.0, mentor2.0 2015|2015-10-12|2015-11-12|NaT||||15.8||2|2|1|1|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||Self|General Site|Amachi|Match Support|M|White||26|28277|Bachelors Degree|Single|Business: Marketing|28273|0|4|Relative|Relative|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|501604887|501605207|31|0|1|503999324|1|0|1|500846761|10|1|500014504||3|1|500000294|-1|500014505, 500015184|-1|0|10|||17161|11|||1|500014505, 500015184|702163000107564368|0
M300|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3851|Yellow|Amachi|2006-08-15|2006-08-21|NaT||||126.5||1|1|1|1|M|Black||16|Yes|Mother|28262|10|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community|Amachi|Match Support|M|White||54|28226|Bachelors Degree|Married|Arts, Entertainment, Sports||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500465506|500465757|31|0|1|500496966|1|0|1|500118121|10|2|500003586||2|2|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294|7432163260389731024|0
M301|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|554|Green||2015-03-23|2015-03-25|2016-09-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.2||1|1|1|1|M|White||16|No|Mother|28078|9|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance|28412|1|4|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500021785|504104035|504106070|1|0|1|504214658|1|0|1|500820084|10|2|-2||4|1||-2||-2|0|5|||17159|12|||1||4565518866290635873|2141487034287122220
M302|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1924|Green|Amachi|2011-11-04|2011-11-30|NaT||||63.2||3|3|1|1|M|Black||16|No|Relative: Other|28205|9|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||33|28226|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|10|Relative|Relative|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501353940|501354219|31|0|1|502710990|1|0|1|500574615|10|2|500003586||2|1|500000294, 500005291|-2||-2|34|2|||17161|11|||1|500000294|1766165378108010922|0
M303|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|123|Green||2014-10-07|2014-10-23|2015-02-23|Child/Family: Moved|Child/Family: Moved||4||1|1|2|2|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||52|28105|Bachelors Degree|Married|Business||2|6|Local Print|Media|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500016847|504043305|504045323|31|0|1|503776239|1|0|1|500781246|10|1|500014504||4|1||-1|500014505, 500014506|-1|0|4|||7439|1|||1||702163000107564368|0
M304|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green|mentor2.0 2016|2016-11-18|2016-11-18|NaT||||3.6||2|2|3|3|M|Black||16|No|Mother|28217|9|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Site|mentor2.0, mentor2.0 2014|Match Support|M|Black||32|28216|Masters Degree|Single|Finance: Accountant|28280|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|501376223|501376502|31|0|1|503976447|31|0|1|500929506|10|1|500014504||2|1|500014505, 500014506|-1|500014505, 500014506, 500016394|-1|0|10|||7462|13|||1|500016394|702163000107564368|6108079083976570810
M305|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|737|Green|mentor2.0, mentor2.0 2014|2014-10-07|2014-10-22|2016-10-28|Volunteer: Moved|Volunteer: Moved||24.2||2|2|1|1|M|Black||16|No|Mother|28217|9|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Site|mentor2.0, mentor2.0 2014|Match Support|M|White||25|28203|Bachelors Degree|Single|Finance|28202|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|501376223|501376502|31|0|1|503969375|1|0|1|500781251|10|1|500014504||4|1|500014505, 500014506|-1|500014506|-1|0|10|||7462|13|||1|500014505, 500014506|702163000107564368|6108079083976570810
M306|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2391|Green||2010-07-26|2010-08-20|NaT||||78.6||1|1|2|2|M|Black||16|No|Mother|28217||One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|502064627|502065051|31|0|1|500773055|3|14|1|500462574|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||702163000107564368|2162928999922594413
M307|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|858|Yellow||2013-02-04|2013-02-11|2015-06-19|Child/Family: Moved|Child/Family: Moved||28.2||2|2|1|1|F|Black||16|No|Mother|28052|8|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||29|28277|Bachelors Degree|Single|Business|28217|2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|502482642|502391834|31|0|2|503118336|1|0|2|500679560|10|2|-2||4|2|500004640, 500005291|-2||-2|0|10|||7464|9|||1||0|0
M308|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2349|Red||2010-09-16|2010-09-22|2017-02-26|Child: Lost interest|Child: Lost interest||77.2||1|1|1|1|F|Hispanic||16|No|Mother|28211|4|One Parent: Female|Unknown||||Yes|Spanish Print|Media|General Community||Match Support|F|Hispanic||38|28202|Bachelors Degree|Single|Tech: Engineer|28202|12|0|Big Day|Special Event|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020753|502264006|502264438|3|0|2|502274748|3|0|2|500470897|10|2|-2||4|3||-2||-2|7063|1|||7456|8|||1||0|0
M309|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|577|Green||2013-10-18|2013-11-18|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19||1|1|1|1|F|Black||16||Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||29|28107|Bachelors Degree|Married|Business: Human Resources|28202|5|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|502766037|502766950|31|0|2|503605985|1|0|2|500720715|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M310|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2313|Green||2009-01-23|2009-02-16|2015-06-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||76||1|1|1|1|M|Black||16|No|Mother|28269|8|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28205|Some College|Married|Retail: Sales|28206|1|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|501525308|501525600|31|0|1|501536144|1|0|1|500335230|10|2|-2||4|1||-2||-2|6854|8|||7464|9|||1||3677730851176818072|4692800185712017442
M311|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|760|Green|PERL 2014-2016|2015-01-29|2015-02-06|NaT||||25||1|1|1|1|M|Black||16|No|Mother|28205|9|One Parent: Female|$10,000 to $14,999|||Y|Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|White||36|28269|Bachelors Degree|Married|Self-Employed, Entrepreneur|28269|7|5|Other|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504063426|504065453|31|0|1|504152304|1|0|1|500810827|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|56|1|||7671|13|||1|500014681|7987165241089060600|5081726734274569781
M312|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3263|Green|Amachi, Cabarrus County|2008-03-04|2008-03-31|NaT||||107.2||1|1|1|1|M|White||16|Yes|GrandMother|28025|10|Grandparents|Unknown||||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|White||46|28027|Bachelors Degree|Divorced|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|501074345|501074618|1|0|1|501158523|1|0|1|500250038|10|2|500003586||2|1|500000294, 500016374|-2|500016374|-2|5635|9|||46|2|||1|500000294, 500016374|3575183301237417432|0
M313|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|598|Red||2014-11-11|2014-12-08|2016-07-28|Child: Lost interest|Child: Lost interest||19.6||2|2|2|2|F|Hispanic||16|No|Mother|28262|10|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|F|White||26|28210|Bachelors Degree|Single|Medical: Admin|28209|1|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500013781|502753870|502751081|3|0|2|503869569|1|0|2|500794392|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||1652521212990559348|0
M314|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0 2016|2015-10-23|2015-11-17|NaT||||15.6||1|1|1|1|M|Hispanic||16|No|Mother|28217|4|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Hispanic||24|28273|Bachelors Degree|Single|Finance|28217|1|8|Self|Self|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|502531929|502532382|3|0|1|504397371|3|0|1|500851402|10|1|500014504||2|1||-1|500015184|-1|0|4|||7464|9|||1|500016394|702163000107564368|0
M315|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2077|Green|Amachi, Project Big, Project Big AND Amachi|2011-06-16|2011-06-30|NaT||||68.2||1|1|1|1|M|Black||16|Yes|Mother|28208|8|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|Amachi, PERL 2014-2016, Project Big, Project Big AND Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Business: Engineer|30357|6|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502549829|502550279|31|0|1|502594393|31|0|1|500541795|10|2|500004772||2|1|500000294, 500004640, 500004901, 500014681|-1||-2|0|4|||7464|9|||1|500000294, 500004640, 500004901|3935539763241716148|0
M316|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2454|Green|Amachi|2010-06-11|2010-06-18|NaT||||80.6||2|2|1|1|M|Black||16|Yes|Aunt|28216||One Parent: Female|Less than $10,000|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||34|20175|Bachelors Degree|Single|Business: Sales|28211|2|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|500934908|500935173|31|0|1|502107314|1|0|1|500456443|10|2|500003586||2|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294|0|0
M317|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|749|Green|PERL 2014-2016|2014-12-18|2015-02-17|NaT||||24.6||1|1|1|1|M|Black||16|No|Mother|28208|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||45|28273|Masters Degree|Married|Finance: Banking|28269|0|1|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|502552947|502553400|31|0|1|503881539|31|0|1|500804943|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||46|2|||1|500014681|702163000107564368|427143067147514567
M318|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1747|Green|Amachi|2012-05-09|2012-05-25|NaT||||57.4||2|2|1|1|F|Multi-race (Black & White)||16|Yes|Aunt|28269|4|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28078|Associate Degree|Married|Tech: Support, Writing|28210|2|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502393980|502394418|36|0|2|502928199|31|0|2|500613992|10|2|500003586||2|1|500005291|-2||-2|0|5|||7462|13|||1|500000294|7102230088759381237|0
M319|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|573|Yellow|mentor2.0, mentor2.0 2014|2014-10-07|2014-10-07|2016-05-02|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||18.8||1|1|1|1|M|Black||16|Yes|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||40|28210|Masters Degree|Married|Business|28281|3|1|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504043202|504045220|31|0|1|503971855|1|0|1|500781225|10|1|500014504||4|2||-1|500014506|-1|0|4|||7671|13|||1|500014505, 500014506|702163000107564368|0
M320|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|756|Green|mentor2.0 2014|2014-10-06|2014-10-06|2016-10-31|Child/Family: Moved|Child/Family: Moved||24.8||2|2|1|1|F|Black||16|No|Father|28217|9|One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|F|White||51|28269|Bachelors Degree|Married|Business|28217|3|0|Self|Self|Big|General Site|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|503712470|503714436|31|0|2|503952262|1|0|2|500780797|10|1|500014504||4|1||-1|500014506|-1|0|4|||7464|9|||1|500014506|702163000107564368|0
M321|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|395|Green||2014-10-07|2014-10-07|2015-11-06|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||13||1|1|2|2|M|American Indian or Alaska Native||16|Yes|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|M|White||34|28202||Married|Consultant||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014, mentor2.0 2016|Match Support|1|0|1|0|277|60|598|500000170|500016847|504050578|504052602|6|0|1|503969533|1|0|1|500781237|10|1|500014504||4|1||-1|500014506, 500016394|-1|0|3|||7462|13|||1||702163000107564368|0
M322|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|239|Green||2014-10-07|2014-10-07|2015-06-03|Child/Family: Moved|Child/Family: Moved||7.9||1|1|1|1|F|Hispanic||16|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||49|28104|Juris Doctorate (JD)|Single|Finance|28203|0|7|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500016847|504043211|504045229|3|0|2|503969563|31|0|2|500781135|10|1|500014504||4|1||-1|500014505, 500014506|-1|0|4|||7462|13|||1||702163000107564368|0
M323|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|124|Red|mentor2.0 2015|2015-10-25|2015-10-26|2016-02-27|Child: Changed school/site|Child: Changed school/site||4.1||1|1|2|2|M|Black||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||Self|General Site|Amachi|Match Support|M|White||40|28210|Bachelors Degree|Married|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|500395499|500395742|31|0|1|501027885|1|0|1|500851881|10|1|500014504||4|3|500000294|-1|500014505, 500015184|-1|0|10|||46|2|||1|500015184|702163000107564368|0
M324|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2429|Yellow|Amachi|2010-07-13|2010-07-13|NaT||||79.8||3|3|1|1|F|Black||16|Yes|Mother|28205|11|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|F|Black||30|28216|Bachelors Degree|Single|Human Services: Non-Profit|28216|0|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|500280148|500188151|31|0|2|502118494|31|0|2|500460767|10|2|500003586||2|2|500000294|-2||-2|0|3|||7464|9|||1|500000294|1010189231295710785|0
M325|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|554|Green||2014-11-07|2014-12-01|2016-06-07|Child: Changed school/site|Child: Changed school/site||18.2||1|1|1|1|M|Black||16|No|Mother|28217|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||32|28012||Single|Business||0|8|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|504089115|504091145|31|0|1|504081485|1|0|1|500793474|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M326|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|784|Green||2015-01-07|2015-01-13|NaT||||25.8||1|1|1|1|F|Black||16|No|Mother|28105|10|One Parent: Female|$35,000 to $39,999|||Y|Yes|Other|Faith Organization|General Community||Match Support|F|Black||27|28227|Bachelors Degree|Single|Finance: Banking|29715|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504090244|504092274|31|0|2|504121323|31|0|2|500806857|10|2|-2||2|1||-2||-2|5635|9|||46|2|||1||8029775806705219538|2359037990929827326
M327|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|157|Green|PERL 2014-2016|2015-11-17|2015-12-14|2016-05-19|Volunteer: Moved|Volunteer: Moved||5.2||1|1|1|1|F|Black||16|No|Mother|28215|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||25|28205|Bachelors Degree|Single|Business|28031|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500017777|503611723|503613600|31|0|2|504295160|1|0|2|500860670|5|2|-2||4|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681|6724463016047116758|0
M328|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|332|Green|mentor2.0, mentor2.0 2015|2015-11-17|2015-11-17|2016-10-14|Child: Changed school/site|Child: Changed school/site||10.9||1|1|1|1|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|M|Black||34|28205|Bachelors Degree|Married|Business: Clerical||3|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|0|1|1|0|277|60|598|500000170|500021786|504449675|504451931|31|0|1|504461244|31|0|1|500860453|10|1|500014504||4|1|500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M329|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|371|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-10-26|2016-10-31|Child: Changed school/site|Child: Changed school/site||12.2||1|1|2|2|M|Black||16|No|Father|28217|9|One Parent: Male|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Black||58|28216|Bachelors Degree|Married|Business: Mgt, Admin|27701|30|0|AA Task Force|Special Event|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504426315|504428570|31|0|1|503796728|31|0|1|500851855|10|1|500014504||4|1|500014505, 500015184|-1|500015184|-1|0|4|||11098|8|||1|500014505, 500015184|702163000107564368|0
M330|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2020|Yellow||2011-07-28|2011-08-19|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||66.4||1|1|1|1|F|Black||16|No|Mother|28208|6|Two Parent|$35,000 to $39,999|||Y|Yes||Relative|General Community||Match Support|F|Hispanic||26|28217|Bachelors Degree|Single|Service: Restaurant||3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502593613|502594130|31|0|2|502601730|3|0|2|500547881|10|2|-2||4|2||-2||-2|0|3|||7464|9|||1||7581500809034284566|0
M331|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1173|Red||2013-02-08|2013-03-08|2016-05-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38.5||1|1|1|1|F|White||16|No|Mother|28082|8|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|White||33|28138|Associate Degree|Divorced|Insurance||2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020753|503225805|503227593|1|0|2|503317460|1|0|2|500680855|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1||0|0
M332|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|NaT||||16||1|1|1|1|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||37|28210|Masters Degree|Single|Business: Mgt, Admin|28203|0|7|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454746|504457004|31|0|2|504339857|1|0|2|500846250|10|1|500014504||2|1||-1|500015184|-1|0|4|||17159|12|||1|500014505, 500015184|702163000107564368|0
M333|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|456|Green||2014-06-30|2014-06-30|2015-09-29|Child: Graduated|Child: Graduated||15||2|2|5|5|M|Black||16|No|Father|28208|8|One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||49|28278|Bachelors Degree|Separated|Finance|28217|7|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|503212298|503824721|31|0|1|500189616|31|0|1|500768234|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M334|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1282|Yellow||2013-02-15|2013-02-27|2016-09-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||42.1||2|2|1|1|M|White||16|No|Mother|28277|7|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||47|28277|Bachelors Degree|Married|Business|28217|20|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502304267|502304699|1|0|1|503343217|1|0|1|500682425|10|2|-2||4|2||-2||-2|0|10|||7671|13|||1||3966805366522644621|7023993708128426307
M335|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|472|Green||2015-10-14|2015-11-13|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||15.5||1|1|1|1|F|Black||16|No|Mother|28216|9|Two Parent|Unknown||||Yes||School|General Community||Match Support|F|White||31|28203|Bachelors Degree|Married|Business: Mgt, Admin|28255|0|9|Other|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|504269922|504272121|31|0|2|504285435|1|0|2|500847702|10|2|-2||4|1||-2||-2|0|4|||18267|3|||1||0|3260639349613832803
M336|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3361|Green||2007-05-10|2007-05-17|2016-07-29|Child: Graduated|Child: Graduated||110.4||1|1|1|1|M|Black||16|No|Mother|28216|8|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|Black||46|28269|||Human Services: Non-Profit||0|0|BBBS National Site|Web Link|Big|General Community|VOL - Adjudicated, VOL - Cultural Comp, VOL - PreMatch|Match Support|1|0|1|0|277|60|598|500000170|500008321|500727291|500727558|31|0|1|500857838|31|0|1|500176403|10|2|-2||4|1||-2|500007913, 500007920, 500011311|-2|0|10|||46|2|||1||0|0
M337|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1832|Red|Project Big|2010-07-20|2010-07-25|2015-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||60.2||1|1|1|1|F|Black||16|No|Mother|28213|4|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|Black||34|28269||Single|Student: College||0|0|UNCC|College Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502179379|502179808|31|0|2|502161458|31|0|2|500461681|10|2|-2||4|3|500004640|-2||-2|0|10|||9221|5|||1|500004640|7376591015108056209|2862823696767408751
M338|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|784|Green||2015-01-07|2015-01-13|NaT||||25.8||1|1|1|1|M|Black||16|No|Mother|28227|8|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community||Match Support|M|White||30|28202|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504034181|504036199|31|0|1|504053608|1|0|1|500806936|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||2129686509389594346|3402014428779854546
M339|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|333|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-10-26|2016-09-23|Child: Changed school/site|Child: Changed school/site||10.9||1|1|2|2|F|Black||16|No|Mother|28208||One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||29|28216|Masters Degree|Single|Medical|30005|0|5|BBBS National Site|Web Link|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504454486|504456744|31|0|2|504300098|31|0|2|500851880|10|1|500014504||4|1|500014505, 500015184|-1|500015184|-1|0|4|||46|2|||1|500014505, 500015184|702163000107564368|0
M340|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|501|Green||2013-11-04|2013-11-15|2015-03-31|Child: Lost interest|Child: Lost interest||16.5||1|1|3|3|M|Black||16|No|Mother|28206|7|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||28|28204|Bachelors Degree|Single|Tech: Computer/Programmer|28204|3|0|Duke Energy|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503624220|503626109|31|0|1|503605851|31|0|1|500727093|10|1|500009132|2128173561|4|1||-1|500014505, 500016394|-1|0|4|||16705|3|||1||7960300212314874874|0
M341|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1384|Green|Cabarrus County|2013-05-17|2013-05-23|NaT||||45.5||1|1|1|1|M|Black||16||Mother|28027|6|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||51|28269|Bachelors Degree|Married|Business: Sales||6|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|503379566|503381423|31|0|1|503407492|1|0|1|500697331|10|2|500016307||2|1|500016374|-2|500016374|-2|34|2|||46|2|||1|500016374|6353565629814722343|8876904578828505776
M342|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Inactive|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-11-06|2015-11-06|NaT||||16||1|1|1|1|M|Black||16|No|Mother|28211|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||27|28120|Masters Degree|Married|Business|28202|3|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504495937|504498222|31|0|1|504355841|1|0|1|500856978|10|1|500014504||3|1||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M343|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3263|Yellow||2006-09-14|2006-09-18|2015-08-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||107.2||1|1|2|2|M|Black||16||Mother|28215|7|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||43|28215|Bachelors Degree|Single|Finance: Banking|28262|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500382177|500382427|31|0|1|500188566|31|0|1|500122093|10|2|-2||4|2||-2||-2|0|10|||7496|10|||1||5741767063897867874|0
M344|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|672|Green||2013-07-08|2013-07-26|2015-05-29|Child/Family: Moved|Child/Family: Moved||22.1||1|1|1|1|F|Black||16|Yes|Mother|28214|7|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||25|28223|Some College|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503472839|503474705|31|0|2|503503841|31|0|2|500702872|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||7089569121628268952|7044657180546140448
M345|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|594|Green||2014-01-22|2014-02-21|2015-10-08|Volunteer: Moved|Volunteer: Moved||19.5||1|1|1|1|M|Black||16|No|Mother|28212|8|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28204|Masters Degree|Single|Finance: Accountant|28202|4|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503395663|503397520|31|0|1|503735537|1|0|1|500744097|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1||2811191761055817959|4912398592230479482
M346|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1582|Red|Project Big, 2010-2012 OJJDP JJI|2011-06-30|2011-06-30|2015-10-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||52||1|1|1|1|M|Black||16|No|Mother|28208|4|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Black||40|28037|Bachelors Degree|Married|Medical: Doctor, Provider||2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502589865|502590381|31|0|1|502625828|31|0|1|500544108|10|2|500004641||4|3|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291|7869308672550505300|0
M347|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|789|Green||2013-11-07|2013-11-07|2016-01-05|Child: Graduated|Child: Graduated||25.9||1|1|2|2|F|Black||16|No|Mother|28202|7|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||41|28025|Some College|Single|Business|28217|4|0|LPL Financial|Workplace Partner|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500017786|503681619|503683584|31|0|2|503680923|31|0|2|500728684|10|1|500009132|2128207319|4|1||-1|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||11247|3|||1||3935539763241716148|0
M348|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-10-26|NaT||||16.4||1|1|2|2|F|Black||16|No|Mother|28208|9|Two Parent|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||38|28209|Bachelors Degree|Single|Business|28202|13|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500021786|504419831|504422084|31|0|2|503985283|1|0|2|500851859|10|1|500014504||2|1|500014505, 500015184|-1|500014506|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M349|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-10-23|2015-10-26|NaT||||16.4||1|1|2|2|F|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||39|28273|Masters Degree|Married|Business: Mgt, Admin|28208|2|0|BBBS National Site|Web Link|Big|General Site|mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500021786|504426322|504428577|31|0|2|503972115|31|0|2|500851410|10|1|500014504||2|1|500014505, 500015184|-1|500014506|-1|0|4|||46|2|||1|500014505, 500015184|702163000107564368|0
M350|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|491|Green|mentor2.0, mentor2.0 2016|2015-10-25|2015-11-02|NaT||||16.1||1|1|1|1|M|Black||16|No|Father|28217|9|One Parent: Male|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Multi-race (Asian & White)||36|28203|Bachelors Degree|Married|Finance||0|11|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504425700|504427955|31|0|1|504445539|37|0|1|500851875|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500016394|702163000107564368|0
M351|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|621|Green|PERL 2014-2016|2015-06-12|2015-06-25|NaT||||20.4||1|1|1|1|M|Black||16|No|Mother|28208|7|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Hispanic||26|28203|Bachelors Degree|Single|Business: Sales|53073|0|5|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503955527|503957535|31|0|1|504285092|3|0|1|500830048|10|2|-2||2|1|500014681|-2||-2|0|5|||17159|12|||1|500014681|8568001799025358453|3380017483853696343
M352|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|349|Green|mentor2.0 2015|2015-10-25|2015-11-17|2016-10-31|Child: Lost interest|Child: Lost interest||11.5||1|1|1|1|M|Hispanic||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||38|28214|Bachelors Degree|Married|Tech: Computer/Programmer||2|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504426175|504428430|3|0|1|504445758|31|0|1|500851856|10|1|500014504||4|1||-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M353|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|833|Green||2014-11-17|2014-11-25|NaT||||27.4||1|1|1|1|M|Black||16|No|Mother|28212||One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|White||35|28211|Masters Degree|Single|Finance: Accountant|28202|2|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503934189|503936197|31|0|1|503918487|1|0|1|500796401|10|2|-2||2|1||-2||-2|0|4|||17101|1|||1||1010189231295710785|6178126991714892144
M354|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|980|Green||2013-11-04|2013-11-04|2016-07-11|Child: Changed school/site|Child: Changed school/site||32.2||1|1|1|1|F|Black||16|No|Mother|28208|8|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||31|28278|Associate Degree|Single|Customer Service|28217|0|8|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|503678291|503680256|31|0|2|503680714|31|0|2|500726845|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M355|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|637|Yellow||2014-01-06|2014-01-10|2015-10-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.9||1|1|3|3|M|Black||16|No|Mother|28269|8|One Parent: Female|$50,000 to $59,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500017777|503556065|503557940|31|0|1|501284751|31|0|1|500741332|10|2|-2||4|2||-2|500007920, 500011315, 500011316|-2|34|2|||132|8|||1||0|3634914038612765160
M356|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|460|Green||2015-01-27|2015-01-29|2016-05-03|Child: Lost interest|Child: Lost interest||15.1||1|1|1|1|F|Black||16|No|Mother|28212|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|Black||26|28213|Bachelors Degree|Single|Finance|28269|2|1|TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500021785|503441463|501290021|31|0|2|504122275|31|0|2|500810468|10|2|-2||4|1||-2||-2|0|4|||130|1|||1||2811191761055817959|7044657180546140448
M357|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0 2015|2015-10-25|2015-11-17|NaT||||15.6||1|1|1|1|M|Black||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|White||57|28211|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504460043|504462301|31|0|1|504314082|1|0|1|500851884|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M358|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-31|2016-11-02|NaT||||4.1||1|1|3|3|M|Black||16|No|Father|28217|9|One Parent: Male|$20,000 to $24,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|Black||28|28204|Bachelors Degree|Single|Tech: Computer/Programmer|28204|3|0|Duke Energy|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831646|504834148|31|0|1|503605851|31|0|1|500921844|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||16705|3|||1||702163000107564368|6641222291370253715
M359|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|910|Green||2013-01-25|2013-01-31|2015-07-30|Volunteer: Moved|Volunteer: Moved||29.9||2|2|1|1|M|Black||16||Mother|28273|7|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|White||32|28273|Bachelors Degree|Single|Business: Mgt, Admin|28217|3|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|502193174|502193603|31|0|1|503100143|1|0|1|500677433|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1||0|0
M360|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1241|Red||2013-02-27|2013-03-05|2016-07-28|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||40.8||2|2|1|1|F|Black||16|No|GrandMother|28206|7|Grandparents|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Multi-race (Asian & White)||28|60654|Bachelors Degree|Single|Business: Mgt, Admin|60601|3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502876870|502878273|31|0|2|503104166|37|0|2|500684838|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||4863631750424600365|0
M361|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|477|Green||2013-12-04|2013-12-09|2015-03-31|Child/Family: Moved|Child/Family: Moved||15.7||1|1|1|1|M|Black||16|No|Mother|28208|8|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||41|28226|Masters Degree|Married|Consultant|28202|8|0|Duke Energy|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503690133|503692098|31|0|1|503605679|1|0|1|500736453|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||5424205421938369753|0
M362|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|925|Red||2013-08-07|2013-08-26|2016-03-08|Child: Lost interest|Child: Lost interest||30.4||1|1|1|1|M|White||16|No|Mother|28273|9|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||63|28226|Masters Degree|Widowed|Business: Marketing||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503484186|503486052|1|0|1|503355490|1|0|1|500706097|10|2|-2||4|3||-2||-2|0|10|||7671|13|1561|2|1||3960869250587139051|1202530717971184330
M363|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2533|Green||2010-03-16|2010-03-31|NaT||||83.2||1|1|1|1|M|Black||16|No|Mother|28212|9|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||26|28215|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|501434147|501434432|31|0|1|501926474|31|0|1|500441566|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||7284449467126735125|2730899240024631792
M364|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2689|Green||2009-06-11|2009-06-22|2016-11-01|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||88.3||1|1|1|1|M|Black||16|No|Mother|28208|8|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||59|28269|Masters Degree|Married|Clergy||0|0|Coca Cola|Workplace Partner|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500020752|501721760|501722098|31|0|1|501755476|1|0|1|500368545|10|2|-2||4|1||-2|500000294|-2|0|10|||9610|3|||1||1227369534771287213|0
M365|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1693|Green||2012-06-20|2012-07-18|NaT||||55.6||2|2|1|1|F|Black||16|No|Mother|28214|4|Two Parent|$40,000 to $44,999|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28210|Masters Degree|Single|Medical: Healthcare Worker||1|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502591898|502592415|31|0|2|503002003|31|0|2|500620503|10|2|-2||2|1|500004640, 500005291|-2||-2|0|4|||7496|10|||1||2611337051335117774|0
M366|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1279|Green||2013-04-11|2013-04-30|2016-10-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||42||1|1|1|1|F|Black||16|No|Mother|28227|4|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||41|28105|High School Graduate|Divorced|Business: Mgt, Admin|28207|6|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502787401|502788587|31|0|2|503122442|1|0|2|500692539|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||8979408036987322141|7044657180546140448
M367|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|549|Green||2014-09-17|2014-09-28|2016-03-30|Volunteer: Time constraint|Volunteer: Time constraint||18||2|2|1|1|F|Black||16|No|Mother|28215|8|Two Parent|$50,000 to $59,999||||No||Self|General Community||Match Support|F|White||26|28202|Bachelors Degree|Single|Business||11|10|Current/Previous Big|Other Big|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500013781|503326540|503328374|31|0|2|503852999|1|0|2|500776439|10|2|-2||4|1||-2||-2|0|10|||17159|12|||1||0|5823903291619049470
M368|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|463|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-11-30|NaT||||15.2||1|1|1|1|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Some Other Race||26|28262|Bachelors Degree|Single|Tech: Engineer|29707|2|5|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504419824|504422077|31|0|1|504455318|41|0|1|500851854|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M369|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green|mentor2.0 2015|2015-10-23|2015-11-11|NaT||||15.8||1|1|1|1|F|Black||16|No|Father|28208|9|One Parent: Male|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||36|29708|Juris Doctorate (JD)|Married|Law|28202|8|8|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504425599|504427854|31|0|2|504349061|1|0|2|500851392|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M370|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|848|Green||2014-10-13|2014-11-10|NaT||||27.9||1|1|1|1|F|Black||16|No|Mother|28262|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||26|28269|Masters Degree|Single|Human Services: Social Worker|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|504004117|504006132|31|0|2|503929259|31|0|2|500783097|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||932861092942387634|0
M371|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|945|Green||2013-11-07|2013-11-11|2016-06-13|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31||1|1|1|1|M|Black||16|No|Mother|28208|7|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||42|28273|High School Graduate|Married|Customer Service|28217|1|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|503681650|503683615|31|0|1|503661517|31|0|2|500728598|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M372|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1503|Green||2013-01-22|2013-01-24|NaT||||49.4||2|2|1|1|F|Black||16|No|Mother|28208|5|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||32|28210|High School Graduate|Single|Business: Sales|28277|0|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502980965|502982410|31|0|2|503091130|1|0|2|500676334|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||2324686837245224089|0
M373|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1694|Green||2012-06-19|2012-07-17|NaT||||55.7||1|1|1|1|M|Black||16|No|Mother|28208|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Sales|28273|2|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502980958|502982410|31|0|1|503008664|1|0|1|500620394|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||932861092942387634|0
M374|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|119|Green|mentor2.0 2015|2015-10-23|2015-11-30|2016-03-28|Child/Family: Moved|Child/Family: Moved||3.9||1|1|2|2|M|Hispanic||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Hispanic||42|28209|Masters Degree|Married|Finance: Banking|28255|12|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504456568|504458826|3|0|1|504380428|3|0|1|500851403|10|1|500014504||4|1||-1|500015184|-1|0|4|||17159|12|||1|500015184|702163000107564368|0
M375|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1868|Yellow|Amachi|2012-01-18|2012-01-25|NaT||||61.4||2|2|1|1|F|Black||16|Yes|Mother|28227|9|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||52|28227|Bachelors Degree|Married|Insurance|28277|14|0|AA Task Force|Special Event|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500847570|500188056|31|0|2|502542379|31|0|2|500592215|10|2|500003586||2|2|500000294|-2|500000294|-2|0|10|||11098|8|||1|500000294|1766165378108010922|0
M376|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-10-23|2015-10-26|NaT||||16.4||1|1|1|1|F|Black||16|Yes|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||35|28203|Masters Degree|Single|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504426348|504428603|31|0|2|504363925|1|0|2|500851384|10|1|500014504||2|1|500014505, 500015184|-1|500014505, 500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M377|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1453|Yellow||2011-06-21|2011-06-27|2015-06-19|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||47.7||2|2|2|2|M|Black||16|No|Mother|28216|8|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|White||53|28117|Bachelors Degree|Married|Real Estate: Realtor|28031|0|0|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|1|0|1|0|277|60|598|500000170|500015820|501842678|501843047|31|0|1|502335257|1|0|1|500542227|10|2|-2||4|2||-2|500000294, 500004901|-2|0|10|||7464|9|||1||6267183121733002735|0
M378|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1065|Yellow||2013-02-15|2013-03-12|2016-02-10|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||35||1|1|1|1|M|Black||16||Mother|28211|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||29|28211|Bachelors Degree||Construction|28208|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502979759|502981210|31|0|1|503234517|1|0|1|500682418|10|2|-2||4|2||-2||-2|0|10|||46|2|||1||4440360203097874486|8247408236389589972
M379|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|554|Yellow||2013-07-16|2013-08-06|2015-02-11|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.2||3|3|2|2|F|Black||16|No|Mother|28226|3|Two Parent|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|F|Black||34|28215|Some College|Single|Finance: Banking|28270|1|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|500826603|500826861|31|0|2|502672644|31|0|2|500703783|10|2|-2||4|2||-2||-2|0|5|||7464|9|||1||4903779310522421428|0
M380|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|579|Green||2014-11-06|2014-11-06|2016-06-07|Child: Changed school/site|Child: Changed school/site||19||2|2|1|1|F|Black||16|No|Mother|28208|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||34|28269|Masters Degree|Single|Business|28217|0|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|503681628|503683593|31|0|2|504024551|31|0|2|500792596|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M381|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|117|Green||2016-10-26|2016-11-04|2017-03-01|Child/Family: Moved|Child/Family: Moved||3.8||1|1|1|1|M|Black||16|Yes|Mother|28208|9|Two Parent|Unknown|||Y|Yes||Relative|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||30|28205|Bachelors Degree|Single|Finance|28202|0|2|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Enrollment|0|1|0|1|277|60|598|500000170|500022907|504888350|504890870|31|0|1|503599329|1|0|1|500920234|10|1|500014504||4|1|500014505, 500016394|-1|500014505, 500016394|-1|0|3|||7464|9|||1||702163000107564368|0
M382|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|481|Green|mentor2.0, mentor2.0 2015|2015-10-12|2015-11-12|NaT||||15.8||1|1|3|3|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||32|28210|Bachelors Degree|Single|Tech: Sales, Mktg|28202|7|6|Duke Energy|Workplace Partner|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454736|504456994|31|0|1|503605671|31|0|1|500846714|10|1|500014504||2|1||-1|500015184|-1|0|4|||16705|3|||1|500014505, 500015184|702163000107564368|0
M383|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|115|Yellow|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|2016-02-29|Child/Family: Moved|Child/Family: Moved||3.8||1|1|1|1|M|Hispanic||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||46|28211|Masters Degree|Married|Finance|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site||Enrollment|0|1|1|0|277|60|598|500000170|500016847|504451240|504453496|3|0|1|504432323|1|0|1|500846210|10|1|500014504||4|2||-1||-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M384|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2093|Green|Project Big, 2010-2012 OJJDP JJI|2011-05-27|2011-06-02|2017-02-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||68.8||1|1|1|1|M|Black||16|No|GrandMother|28208|8|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||36|28205|Masters Degree|Living w/ Significant Other|Journalist/Media|28202|3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020910|502552438|502552891|31|0|1|502549491|1|0|1|500538826|10|2|-2||4|1|500004640, 500005291|-2||-2|0|10|||7464|9|||1|500004640, 500005291|1653226628427425023|0
M385|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|317|Green|mentor2.0, mentor2.0 2015|2015-12-02|2015-12-02|2016-10-14|Child: Lost interest|Child: Lost interest||10.4||1|1|1|1|M|Black||16|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||39|28277|Masters Degree|Married|Business: Mgt, Admin|28273|1|2|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504447817|504450073|31|0|1|504422986|1|0|1|500864580|10|1|500014504||4|1||-1|500015184|-1|0|4|||17159|12|||1|500014505, 500015184|702163000107564368|0
M386|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|81|Yellow||2015-10-16|2015-10-31|2016-01-20|Child: Severity of challenges|Child: Severity of challenges||2.7||1|1|2|2|M|Black||16|No|Mother|28202|8|Two Parent|Unknown||||Yes||Relative|General Site||Match Support|F|Black||44|28216|Bachelors Degree|Single|Business||2|0|LPL Financial|Workplace Partner|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500015820|504416080|504418332|31|0|1|504349689|31|0|2|500848793|10|1|500009132|2128207319|4|2||-1||-1|0|3|||11247|3|||1||3935539763241716148|0
M387|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|620|Red|PERL 2014-2016|2014-10-31|2014-11-17|2016-07-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.4||1|1|1|1|F|Black||16|No|Mother|28277|7|One Parent: Female|$40,000 to $44,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||31|28209|Juris Doctorate (JD)|Single|Law|28210|1|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500008321|503746685|503755760|31|0|2|503961087|1|0|2|500790718|10|2|-2||4|3|500014681|-2|500014681|-2|34|2|||17159|12|||1|500014681|7883015200677941272|0
M388|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2427|Green||2009-02-19|2009-02-26|2015-10-20|Volunteer: Moved|Volunteer: Moved||79.7||1|1|1|1|M|Black||16|No|Mother|28227|7|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||33|10019|Bachelors Degree|Single|Business: Marketing|28202|2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|500765381|500739190|31|0|1|501579025|1|0|1|500342803|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||8202428416367135871|0
M389|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|290|Red|PERL 2014-2016|2015-01-20|2015-02-13|2015-11-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||9.5||1|1|1|1|M|Black||16|No|Mother|28212|8|One Parent: Female|$35,000 to $39,999||||Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|White||57|28226|Some College|Single|Business: Sales|28134|10|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500008321|504129007|504131049|31|0|1|504137446|1|0|1|500809001|10|2|-2||4|3|500014681|-2|500014681|-2|56|1|||17159|12|||1|500014681|2811191761055817959|2197933814735019388
M390|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1155|Green||2012-04-01|2012-04-30|2015-06-29|Child/Family: Moved|Child/Family: Moved||37.9||1|1|1|1|F|Multi-Race (None of the above)||16|No|Father|28214|5|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher|28078|0|8|Self|Self|Big|General Community|Project Big|Match Support|1|0|1|0|277|60|598|500000170|500008321|502828137|502829415|7|0|2|502446364|31|0|2|500607445|10|2|-2||4|1||-2|500004640|-2|0|10|||7464|9|||1||7089569121628268952|0
M391|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1686|Green|2010-2012 OJJDP JJI|2011-05-05|2011-05-17|2015-12-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||55.4||1|1|1|1|M|Black||16|No|Mother|28215|6|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28215||Single|Law: Police Officer||14|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502402515|502402953|31|0|1|502537081|31|0|1|500535130|10|2|-2||4|1|500005291|-2||-2|34|2|||7464|9|||1|500005291|5741767063897867874|0
M392|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2239|Green|2010-2012 OJJDP JJI|2011-01-14|2011-01-19|NaT||||73.6||1|1|2|2|F|Black||16|No|Mother|28216|7|Two Parent|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28209|Bachelors Degree|Single|Law|28273|5|0|Relative|Relative|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500021785|502244776|502245202|31|0|2|502143351|1|0|2|500511171|10|2|-2||2|1|500005291|-2|500000294|-2|0|4|||17161|11|||1|500005291|1653226628427425023|0
M393|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|NaT||||16||1|1|2|2|M|Hispanic||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||31|28269|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|3|Neighbor/Friend|Neighbor/Friend|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500021786|504440280|504442536|3|0|1|503028265|1|0|1|500846203|10|1|500014504||2|1||-1|500014505, 500014506|-1|0|4|||7496|10|||1|500014505, 500015184|702163000107564368|0
M394|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-27|2016-11-04|NaT||||4||1|1|1|1|F|Hispanic||15|No|Mother|28217|9|Two Parent|Less than $10,000||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Hispanic||29|28206|Masters Degree|Single|Architect|28204|1|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831472|504833974|3|0|2|504339626|3|0|2|500920558|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500015184|-1|0|4|||17159|12|||1||702163000107564368|0
M395|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1149|Green||2013-12-05|2014-01-06|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||37.7||1|1|1|1|F|Black||15|Yes|Mother|28216|7|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||32|28270|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503606415|503608292|31|0|2|503665457|1|0|2|500736909|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1||8758769076374727509|4206170845868125206
M396|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|363|Green|mentor2.0 2015|2016-03-08|2016-03-09|NaT||||11.9||1|1|1|1|F|Black||15|No|Father|28208|9|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|F|Black||45|28211|Masters Degree|Divorced|Finance: Auditor|28255|1|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504447831|504450087|31|0|2|504349089|31|0|2|500883507|10|1|500014504||2|1||-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M397|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|578|Green||2013-10-18|2013-11-15|2015-06-16|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19||1|1|3|3|F|Black||15|No|Mother|28205|9|One Parent: Female|Unknown|||Y|Yes||School|General Community||Enrollment|F|White||29|28209|Bachelors Degree|Single|Business|28202|6|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503635439|503637389|31|0|2|503605799|1|0|2|500720716|5|1|500009132|2128173561|4|1||-2|500014681|-1|0|4|||16705|3|||1||6286214584598985826|0
M398|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1240|Green||2013-08-16|2013-08-26|2017-01-17|Volunteer: Moved|Volunteer: Moved||40.7||1|1|1|1|F|Black||15|No|Mother|28216|6|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||37|28078|Bachelors Degree|Single|Medical|46285|6|5|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503503500|503505371|31|0|2|503390470|1|0|2|500706999|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||5441374193599827162|0
M399|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|343|Green|mentor2.0, mentor2.0 2015|2015-10-12|2015-11-06|2016-10-14|Volunteer: Time constraint|Volunteer: Time constraint||11.3||1|1|1|1|M|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|RTBM|M|Asian||49|28210|Masters Degree|Married|Business||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504445105|504447361|31|0|1|504447607|4|0|1|500846715|7|1|500014504||4|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M400|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-17|NaT||||15.6||1|1|1|1|F|Hispanic||15|Yes|Mother|28273|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||35|28204|Bachelors Degree|Single|Business: Sales|28202|1|7|AA Task Force|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454672|504456930|3|0|2|503885836|1|0|2|500846237|10|1|500014504||2|1||-1|500014505, 500015184|-1|0|4|||9223|3|||1|500014505, 500015184|702163000107564368|0
M401|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|963|Green||2014-06-23|2014-07-18|NaT||||31.6||2|2|1|1|F|Multi-Race (None of the above)||15|No|Mother|28213|8|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||32|28209|Bachelors Degree|Single|Business: Sales|45236|0|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|501725168|501724831|7|0|2|503828482|1|0|2|500767445|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||6381341368426079638|0
M402|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|672|Green||2015-04-28|2015-05-05|NaT||||22.1||1|1|1|1|F|White||15|No|Mother|28227|8|One Parent: Female|$35,000 to $39,999||||Yes||School|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Law: Paralegal|28211|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504235352|504237484|1|0|2|504200139|1|0|2|500825073|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||1421169092898167719|8961132295198487522
M403|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-10-14|2015-11-06|NaT||||16||1|1|1|1|M|Hispanic||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|M|White||40|28226|Bachelors Degree|Married|Finance||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504449679|504451935|3|0|1|504447687|1|0|1|500847841|10|1|500014504||2|1|500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M404|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1245|Green||2013-09-10|2013-09-27|2017-02-23|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||40.9||1|1|1|1|M|Black||15|No|Mother|28215|10|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||47|28215|Bachelors Degree|Married|Finance: Banking|28269|13|6|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020910|503318447|503320281|31|0|1|503537303|31|0|1|500709889|10|2|-2||4|1||-2||-2|0|10|||7458|9|||1||675142027733303647|6178126991714892144
M405|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green|mentor2.0 2016|2015-10-23|2015-11-11|NaT||||15.8||1|1|1|1|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||35|28273|Bachelors Degree|Single|Business: Engineer|28273|0|8|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504425892|504428147|31|0|2|504352616|31|0|2|500851391|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||17159|12|||1|500016394|702163000107564368|0
M406|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|354|Green|mentor2.0 2015|2015-10-12|2015-10-26|2016-10-14|Child: Lost interest|Child: Lost interest||11.6||1|1|1|1|F|Hispanic||15|Yes|Mother|28217||One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|White||34|28204|Bachelors Degree|Married|Finance: Banking|28204|2|2|Other|Workplace Partner|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504451307|504453563|3|0|2|504356262|1|0|2|500846709|10|1|500014504||4|1|500015184|-1|500015184|-1|0|4|||18267|3|||1|500015184|702163000107564368|0
M407|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|448|Green|PERL 2014-2016|2015-11-30|2015-12-15|NaT||||14.7||1|1|1|1|F|Black||15|No|Mother|28215|9|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||26|28213|Bachelors Degree|Single|Business: Mgt, Admin|28105|2|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500021785|504393421|504395660|31|0|2|504395484|31|0|2|500863556|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||46|2|||1|500014681|414551800606805272|5081726734274569781
M408|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|617|Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2015-05-20|2015-06-29|NaT||||20.3||1|1|1|1|F|Hispanic||15|No|Mother|28215|9|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|White||45|28205|Associate Degree|Married|Tech: Computer/Programmer|28202|10|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|504154291|504156341|3|0|2|503862054|1|0|2|500827743|10|2|-2||2|1|500011312, 500014681|-2|500014681|-2|0|10|||17159|12|||1|500011312, 500014681|0|0
M409|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|860|Green||2014-10-23|2014-10-29|NaT||||28.3||1|1|1|1|F|Black||15|No|Mother|28262||One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||37|28208|Bachelors Degree|Single|Tech: Research/Design|28202|3|8|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|504031334|503917391|31|0|2|503882331|1|0|2|500787330|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||0|8283117761446993531
M410|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|206|Green||2014-11-07|2014-11-07|2015-06-01|Child: Lost interest|Child: Lost interest||6.8||3|3|1|1|F|Black||15|No|Mother|28217|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||34|28269|Masters Degree|Single|Customer Service|28269|1|2|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|503216820|503218601|31|0|2|504024735|31|0|2|500793488|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M411|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-10-26|NaT||||16.4||1|1|1|1|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||25|28204|Masters Degree|Single|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504419837|504422090|31|0|2|504368264|31|0|2|500851860|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M412|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|579|Green||2013-10-14|2013-11-15|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19||1|1|2|2|M|Hispanic||15|Yes|Father|28216|7|One Parent: Female|Unknown||||Yes||School|General Community|VOL - Mentoring Hispanic Youth|Enrollment|M|White||34|28202|Masters Degree|Single|Business: Engineer|28202|4|5|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503602228|503612230|3|0|1|503605726|1|0|1|500719010|5|1|500009132|2128173561|4|1|500011312|-2||-1|0|4|||16705|3|||1||7960300212314874874|0
M413|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2039|Yellow|2010-2012 OJJDP JJI|2011-02-17|2011-03-02|2016-09-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||67||1|1|1|1|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28205|Masters Degree|Single|Education: Teacher|2122|1|5|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501833026|501833394|31|0|2|502451325|1|0|2|500518305|10|2|-2||4|2|500005291|-2|500000294|-2|0|10|||7464|9|||1|500005291|702163000107564368|0
M414|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|463|Green|mentor2.0, mentor2.0 2016|2015-10-23|2015-11-30|NaT||||15.2||1|1|1|1|M|Hispanic||15|Yes|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Hispanic||24|28202|Bachelors Degree|Living w/ Significant Other|Finance: Banking|28255|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504444913|504447169|3|0|1|504272227|3|0|1|500851395|10|1|500014504||2|1||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500016394|702163000107564368|0
M415|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Pending Match|399|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-17|2016-12-20|Volunteer: Moved|Volunteer: Moved||13.1||1|2|1|1|M|Hispanic||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0|Pending Match|M|White||27|28202|Bachelors Degree|Single|Finance: Banking|28202|1|9|Neighbor/Friend|Neighbor/Friend|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504447870|504450126|3|0|1|504320091|1|0|1|500846235|9|1|500014504||4|1|500014505|-1|500015184|-1|0|4|||7496|10|||1|500014505, 500015184|702163000107564368|0
M416|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|981|Green||2014-06-19|2014-06-30|NaT||||32.2||4|4|1|1|M|White||15|No|Mother|28031|6|One Parent: Female|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28031|Bachelors Degree|Separated|Business: Mgt, Admin|28206|20|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500796261|500796529|1|0|1|503790153|1|0|1|500767163|10|2|-2||2|1|500005291|-2||-2|34|2|||7496|10|||1||2798582775385400033|0
M417|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|343|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|2016-10-14|Child: Lost interest|Child: Lost interest||11.3||1|1|2|2|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Asian||49|28210|Masters Degree|Married|Education: Teacher||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504440272|504442528|31|0|2|503281135|4|0|2|500846208|10|1|500014504||4|1||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M418|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1356|Green||2013-06-10|2013-06-20|NaT||||44.6||2|2|1|1|M|Black||15|No|Mother|28215|10|One Parent: Female|$40,000 to $44,999||||Yes||Self|General Community||Match Support|M|Black||30|28205|Bachelors Degree|Single|Self-Employed, Entrepreneur|28206|5|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501194563|501194837|31|0|1|503477116|31|0|1|500700141|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||6875312010577189564|5832494112856974468
M419|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|491|Green|mentor2.0 2015|2015-10-25|2015-11-02|NaT||||16.1||1|1|1|1|F|Black||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|White||28|28269|Masters Degree|Single|Business|28202|4|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504444978|504447234|31|0|2|504357304|1|0|2|500851864|10|1|500014504||2|1|500015184|-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M420|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1678|Red||2012-07-06|2012-07-24|2017-02-26|Child: Lost interest|Child: Lost interest||55.1||1|1|1|1|M|Multi-race (Black & Hispanic)||15||Mother|28270|8|One Parent: Female|$25,000 to $29,999|||Y|No||Therapist/Counselor|General Community||Match Support|M|White||51|28173|Bachelors Degree|Married|Consultant|28173|1|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020753|503005868|503007379|38|0|1|502935610|1|0|1|500623124|10|2|-2||4|3||-2||-2|0|5|||7671|13|||1||5994075768656267011|6580743739284115546
M421|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3057|Yellow|Amachi, Cabarrus County|2008-10-14|2008-10-23|NaT||||100.4||2|2|1|1|M|White||15|Yes|Mother|28083||One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|Amachi, Cabarrus County|Match Support|M|White||35|28083|Masters Degree|Single|Business: Mgt, Admin|28027|2|3|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|500496598|500496849|1|0|1|501383928|1|0|1|500299090|10|2|500003586||2|2|500000294, 500016374|-2|500016374|-2|34|2|||7464|9|||1|500000294, 500016374|0|8022741264464756696
M422|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|658|Green||2015-05-07|2015-05-19|NaT||||21.6||1|1|1|1|F|Black||15|No|Mother|28214|9|Two Parent|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|Black||22|28223||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504023342|504060686|31|0|2|504173078|31|0|2|500826184|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||216500609169513656|0
M423|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|132|Green||2015-06-11|2015-08-20|2015-12-30|Child/Family: Moved|Child/Family: Moved||4.3||1|1|1|1|F|Black||15|No|Mother|28215|8|Two Parent|Unknown||||Yes||Self|General Community||Match Support|F|Multi-race (Black & Asian)||23|28206|High School Graduate|Single|Business|28273|1|6|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500020990|504207073|504025357|31|0|2|504201268|39|0|2|500829987|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||9076057728106637014|6720484407795402036
M424|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|340|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|2016-10-11|Child: Changed school/site|Child: Changed school/site||11.2||1|1|2|2|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||34|28262|Bachelors Degree|Single|Insurance|28277|0|4|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Enrollment|0|1|1|0|277|60|598|500000170|500021786|504440264|504442520|31|0|2|504267500|31|0|2|500846201|10|1|500014504||4|1||-1|500014505, 500016394|-1|0|4|||17159|12|||1|500014505, 500015184|702163000107564368|0
M425|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|331|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-18|2016-10-14|Child: Lost interest|Child: Lost interest||10.9||1|1|3|3|M|Hispanic||15|Yes|Father|28208|9|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|M|Black||28|28204|Bachelors Degree|Single|Tech: Computer/Programmer|28204|3|0|Duke Energy|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500021786|504454695|504456953|3|0|1|503605851|31|0|1|500846245|10|1|500014504||4|1||-1|500014505, 500016394|-1|0|4|||16705|3|||1|500014505, 500015184|702163000107564368|0
M426|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|330|Red|PERL 2014-2016|2015-05-05|2015-06-02|2016-04-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.8||1|1|1|1|M|Black||15|No|Mother|28273|8|One Parent: Female|$35,000 to $39,999||||No|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||30|28208|Bachelors Degree|Single|Self-Employed, Entrepreneur|28078|2|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500013781|504159888|504161941|31|0|1|504240720|1|0|1|500825834|10|2|-2||4|3|500014681|-2|500014681|-2|34|2|||17159|12|||1|500014681|6505995099520362521|8491998754880714879
M427|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|476|Green|PERL 2014-2016, Cabarrus County|2015-11-10|2015-11-17|NaT||||15.6||1|1|1|1|M|White||15|Yes|Mother|28025|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28025|High School Graduate|Single|Business: Sales|28025|5|0|Local TV|Media|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|503821678|503823656|1|0|1|504468148|1|0|1|500858177|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7438|1|||1|500014681, 500016374|6750834084344455219|7044657180546140448
M428|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||1|1|1|1|F|Hispanic||15|No|Mother|28209|9|Two Parent|$15,000 to $19,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||22|28208|Bachelors Degree|Single|Journalist/Media|27413|0|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504883840|504886360|3|0|2|504742660|31|0|2|500921974|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M429|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|412|Green||2015-04-29|2015-05-27|2016-07-12|Child: Changed school/site|Child: Changed school/site||13.5||1|1|2|2|M|Black||15|No|Mother|28214|8|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||33|28216|Bachelors Degree|Single|Customer Service||2|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504287270|504289471|31|0|1|504024992|1|0|1|500825343|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M430|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|579|Green||2014-02-20|2014-02-27|2015-09-29|Child: Graduated|Child: Graduated||19||1|1|2|2|F|Black||15|No|Mother|28208|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Multi-Race (None of the above)||34|28134|Some College|Single|Business|28217|2|4|LPL Financial|Workplace Partner|Big|General Site||RTBM|1|0|1|0|277|60|598|500000170|500017786|503805173|503807150|31|0|2|503799347|7|0|2|500750061|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M431|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|31|Green|mentor2.0 2015|2015-10-23|2015-11-30|2015-12-31|Child: Changed school/site|Child: Changed school/site||1||1|1|2|2|F|Black||15|No|Mother|28208||One Parent: Female|Unknown||||Yes||Relative|General Site|mentor2.0 2015|Match Support|F|Black||28|28216|Bachelors Degree|Single|Business|28120|0|6|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500017786|504425766|504428021|31|0|2|504287751|31|0|2|500851406|10|1|500014504||4|1|500015184|-1|500016394|-1|0|3|||17159|12|||1|500015184|702163000107564368|0
M432|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|NaT||||16||1|1|1|1|F|Black||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||37|28202|Bachelors Degree|Living w/ Significant Other|Personal Trainer/Coach|28202|4|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504445152|504447408|31|0|2|504355816|1|0|2|500846231|10|1|500014504||2|1||-1|500014505, 500015184|-1|0|4|||7462|13|||1|500014505, 500015184|0|0
M433|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|927|Green|Cabarrus County|2014-08-18|2014-08-23|NaT||||30.5||1|1|1|1|F|Black||15|Yes|GrandMother|28075|9|Grandparents|$10,000 to $14,999|||Y|Yes||Relative|General Community|Amachi, Cabarrus County|Match Support|F|Black||33|28269|PHD|Single|Education: Admin|28081|4|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|503532788|503534663|31|0|2|503939365|31|0|2|500772617|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|3|||17159|12|||1|500016374|4764211246455367412|7044657180546140448
M434|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|333|Green|mentor2.0 2015|2015-10-23|2015-11-30|2016-10-28|Child: Changed school/site|Child: Changed school/site||10.9||1|1|1|1|M|Hispanic||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|Asian||30|28202|Bachelors Degree|Single|Finance|28202|1|9|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504426069|504428324|3|0|1|504350928|4|0|1|500851385|10|1|500014504||4|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500015184|702163000107564368|0
M435|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1077|Red||2013-08-19|2013-08-30|2016-08-11|Child/Family: Moved|Child/Family: Moved||35.4||2|2|1|1|F|Multi-race (Black & Hispanic)||15|Yes|Mother|28217|9|Two Parent|$35,000 to $39,999||||Yes||Self|General Community||Match Support|F|Black||28|28269|Bachelors Degree|Single|Business||0|7|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502990571|502992028|38|0|2|503400909|31|0|2|500707095|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||1227369534771287213|447407360804656930
M436|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-10-26|NaT||||16.4||1|1|1|1|M|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|White||38|28210|Masters Degree|Single|Education|28273|0|4|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504444999|504447255|31|0|1|504448559|1|0|1|500851865|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M437|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|475|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-18|NaT||||15.6||1|1|2|2|F|Hispanic||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||54|28210|Masters Degree|Married|Tech: Computer/Programmer|28202|1|10|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500021786|504445133|504447389|3|0|2|503969458|1|0|2|500846238|10|1|500014504||2|1||-1|500014506|-1|0|4|||7671|13|||1|500014505, 500015184|702163000107564368|0
M438|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green|mentor2.0|2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|F|Black||15|No|Mother|28216|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||28|28216|Bachelors Degree|Single|Business|28120|0|6|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500021786|504425789|504428044|31|0|2|504287751|31|0|2|500929526|10|1|500014504||2|1|500014505, 500015184|-1|500016394|-1|0|4|||17159|12|||1|500014505|702163000107564368|0
M439|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|352|Green|mentor2.0 2015|2015-10-23|2015-11-11|2016-10-28|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||11.6||2|2|2|2|F|Black||15|No|Mother|28216|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||24|28202||Single|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504425789|504428044|31|0|2|504353872|1|0|2|500851389|10|1|500014504||4|1|500014505, 500015184|-1|500014505, 500015184|-1|0|4|||17159|12|||1|500015184|702163000107564368|0
M440|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|189|Green||2016-08-15|2016-08-30|NaT||||6.2||1|1|1|1|M|Multi-race (Black & Hispanic)||15|No|Mother|28269|8|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|M|White||33|28203|Juris Doctorate (JD)|Married|Law: Lawyer|28202|2|7|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504148143|504125727|38|0|1|504559007|1|0|1|500903465|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||2811191761055817959|887254134148570071
M441|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1269|Red|Project Big, Project Big AND Amachi|2011-12-16|2012-02-08|2015-07-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||41.7||1|1|2|2|M|Black||15|No|Mother|28214|4|One Parent: Female|Unknown||||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|M|White||33|28214|Associate Degree|Single|Law: Security Officer|28208|2|9|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502317500|502317931|31|0|1|502658498|1|0|1|500587614|10|2|-2||4|3|500004640, 500004901|-2||-2|0|4|||7464|9|||1|500004640, 500004901|7089569121628268952|0
M442|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1356|Green|Amachi|2013-06-13|2013-06-20|NaT||||44.6||2|2|1|1|F|Black||15|Yes|Mother|28270|9|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||35|28205|Bachelors Degree|Married|Business: Mgt, Admin|28217|5|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501224282|501224558|31|0|2|503347558|1|0|2|500700583|10|2|-2||2|1|500000294|-2||-2|5635|9|||46|2|||1|500000294|0|0
M443|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|326|Green|PERL 2014-2016|2014-11-07|2014-11-07|2015-09-29|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||10.7||2|2|1|1|F|Black||15|No|Mother|28208|7|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|Black||41|29715|Bachelors Degree|Married|Business|28217|1|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|504089161|504091191|31|0|2|504078362|31|0|2|500793380|10|1|500009132|2128207319|4|1|500014681|-1||-1|0|4|||11247|3|||1|500014681|3935539763241716148|0
M444|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|255|Green|PERL 2014-2016|2015-10-16|2015-10-30|2016-07-11|Child: Changed school/site|Child: Changed school/site||8.4||2|2|1|1|F|Black||15|No|Mother|28208|7|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|White||36|28031|Bachelors Degree|Single|Business: Human Resources|28217|1|0|LPL Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500015820|504089161|504091191|31|0|2|504393611|1|0|2|500848778|10|1|500009132|2128207319|4|1|500014681|-1|500014681|-1|0|4|||11247|3|||1|500014681|3935539763241716148|0
M445|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3192|Red|Amachi|2007-04-26|2007-04-30|2016-01-25|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||104.9||1|1|1|1|M|Black||15|Yes|Mother|28215|7|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|M|White||34|29708|Bachelors Degree|Single|Self-Employed, Entrepreneur|29708|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500545470|501750989|31|0|1|500815012|1|0|1|500173957|10|2|500003586||4|3|500000294|-2|500000294|-2|0|3|||2238|7|||1|500000294|2811191761055817959|0
M446|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|219|Yellow||2014-07-22|2014-07-29|2015-03-05|Volunteer: Time constraint|Volunteer: Time constraint||7.2||1|1|1|1|M|White||15|No|Mother|28226|7|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||RTBM|M|White||73|28277|High School Graduate|Married|Arts, Entertainment, Sports||0|0|Radio|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503834613|503836592|1|0|1|503790527|1|0|1|500770182|7|2|-2||4|2||-2||-2|0|10|||131|1|||1||384008102559124244|5465455237646252584
M447|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|391|Green|PERL 2014-2016|2015-05-29|2015-05-29|2016-06-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.8||1|1|1|1|F|Black||15|No|Mother|28227|8|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||22|28262||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504081466|504083495|31|0|2|504098772|1|0|2|500828761|10|2|-2||4|1|500014681|-2||-2|34|2|||17159|12|||1|500014681|1421169092898167719|4786128411006480901
M448|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|1455|Green||2011-10-03|2011-10-11|2015-10-05|Child: Changed school/site|Child: Changed school/site||47.8||4|4|1|1|M|Black||15||Mother|28213|6|One Parent: Female|Unknown||||No||School|General Site|2010-2012 OJJDP JJI|Match Support|M|Black||29|28269|Bachelors Degree|Single|Tech: Computer/Programmer|28269|0|4|Other|BBBS Board/Staff|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|501076082|501076355|31|0|1|502687269|31|0|1|500560406|10|1|500000295|2128173561|4|1|500005291|-1||-1|0|4|||7671|13|||1||7960300212314874874|0
M449|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|495|Green||2013-10-14|2013-10-24|2015-03-03|Volunteer: Moved|Volunteer: Moved||16.3||1|1|1|1|M|Black||15|No|Mother|28216|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||RTBM|M|Black||27|28216|Bachelors Degree|Single|Business: Engineer|28202|0|1|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|503533022|503534897|31|0|1|503534544|31|0|1|500718872|7|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||7883015200677941272|1786514887916898235
M450|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|380|Green|PERL 2014-2016|2015-03-05|2015-03-09|2016-03-23|Volunteer: Time constraint|Volunteer: Time constraint||12.5||1|1|1|1|F|Black||15|No|Mother|28208|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||28|28204|Bachelors Degree|Single|Finance: Accountant|28277|0|3|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500018851|504075196|504048929|31|0|2|504108003|1|0|2|500817229|10|2|-2||4|1|500014681|-2|500014681|-2|0|4|||46|2|||1|500014681|932861092942387634|7044657180546140448
M451|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|82|Yellow||2015-10-16|2015-10-30|2016-01-20|Child/Family: Moved|Child/Family: Moved||2.7||1|1|2|2|M|Black||15|No|Mother|28217|8|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site||Match Support|M|White||27|29710|Bachelors Degree|Married|Business: Human Resources|28217|3|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504428620|504430875|31|0|1|504035546|1|0|1|500848781|10|1|500009132|2128207319|4|2||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M452|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1564|Green|VOL - PreMatch|2012-11-12|2012-11-24|NaT||||51.4||2|2|1|1|F|Black||15|No|GrandMother|28205|5|Grandparents|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||31|28209|Associate Degree|Married|Retail: Mgt|28134|4|3|UNCC|College Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502859187|500187987|31|0|2|503090888|1|0|2|500658723|10|2|-2||2|1||-2||-2|0|10|||9221|5|||1|500007920|7960300212314874874|0
M453|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2533|Green||2010-03-03|2010-03-31|NaT||||83.2||1|1|1|1|M|White||15|No|Mother|29710|8|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Community||Match Support|M|White||38|28210|||Business||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502030263|502030662|1|0|1|501923553|1|0|1|500438867|10|2|-2||2|1||-2||-2|6855|8|||7464|9|||1||0|0
M454|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|579|Green||2013-10-14|2013-11-15|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19||1|1|3|3|M|Black||15|No|Mother|28205|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||30|29707|Bachelors Degree|Married|Business: Engineer|28202|6|2|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503634083|503636024|31|0|1|503605644|1|0|1|500719001|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M455|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2206|Green|2010-2012 OJJDP JJI, Cabarrus County|2011-02-03|2011-02-21|NaT||||72.5||2|2|1|1|F|White||15|No|Father|28025||One Parent: Male|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|White||43|28027|Associate Degree|Married|Student: College||4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|501247269|500341682|1|0|2|501914025|1|0|2|500515263|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7496|10|||1|500005291, 500016374|0|0
M456|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|349|Green|mentor2.0 2015|2015-10-25|2015-11-17|2016-10-31|Volunteer: Moved|Volunteer: Moved||11.5||1|1|1|1|M|Hispanic||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|M|White||23|28203|Bachelors Degree|Single|Law: Lawyer|28202|0|1|Recruitment Event|Workplace Partner|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017786|504444952|504447208|3|0|1|504284272|1|0|1|500851876|10|1|500014504||4|1|500015184|-1|500015184|-1|0|4|||7446|3|||1|500015184|702163000107564368|0
M457|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1530|Yellow|Amachi|2012-04-05|2012-04-12|2016-06-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||50.3||1|1|1|1|F|Black||15|Yes|Mother|28208|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Multi-race (Black & White)||33|28269|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502809446|502810724|31|0|2|502909383|36|0|2|500608444|10|2|500003586||4|2|500000294|-2||-2|0|10|||7462|13|||1|500000294|5424205421938369753|0
M458|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1324|Green||2013-07-17|2013-07-22|NaT||||43.5||4|5|2|2|F|Black||15||Aunt|28213|8|Two Parent|Unknown||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||24|28262|Some College|Single|Student: College|28216|0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|500570756|500214349|31|0|2|502889143|31|0|2|500703847|10|2|-2||2|1|500004640, 500005291|-2||-2|0|4|||7464|9|||1||6381341368426079638|0
M459|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|343|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-06|2016-10-14|Volunteer: Time constraint|Volunteer: Time constraint||11.3||1|1|1|1|M|Black||15|No|Father|28208|9|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|M|White||24|28270|Bachelors Degree|Single|Business|28217|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504440287|504442543|31|0|1|504382284|1|0|1|500846211|10|1|500014504||4|1||-1|500014505, 500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M460|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|394|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment, PERL 2014-2016|2015-12-22|2016-01-30|2017-02-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||12.9||1|1|2|2|M|Black||15|No|Mother|28269|8|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||32|28202|Masters Degree|Single|Finance: Accountant|28202|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020910|504397554|504399794|31|0|1|504206321|1|0|1|500869278|10|2|-2||4|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||17159|12|||1|500007920, 500011315, 500011316, 500014681|3677730851176818072|5898021503604846505
M461|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-17|NaT||||15.6||1|1|1|1|M|Black||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||Relative|General Site||Match Support|M|White||32|28211||Married|Student: College||0|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454712|504456970|31|0|1|504214615|1|0|1|500846252|10|1|500014504||2|1||-1|500014505|-1|0|3|||17159|12|||1|500014505, 500015184|702163000107564368|0
M462|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|650|Yellow|Cabarrus County|2015-05-05|2015-05-27|NaT||||21.4||1|1|1|1|F|Black||15|No|Mother|28027|9|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community|2010-2012 OJJDP JJI, Cabarrus County|Match Support|F|White||27|28262|Associate Degree|Single|Self-Employed, Entrepreneur|28217|3|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502501997|502502446|31|0|2|504227306|1|0|2|500825847|10|2|500016307||2|2|500005291, 500016374|-2|500016374|-2|0|10|||17159|12|||1|500016374|1557072896577419067|2581014289501540602
M463|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2016|2015-10-09|2015-11-06|NaT||||16||1|1|1|1|M|Hispanic||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||67|28210||Married|Retired||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504440292|504442548|3|0|1|504364944|1|0|1|500846206|10|1|500014504||2|1||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500016394|702163000107564368|0
M464|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1621|Green|Amachi, Project Big, Project Big AND Amachi|2011-11-08|2011-12-02|2016-05-10|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||53.3||2|2|1|1|F|Black||15|Yes|Mother|28217|4|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||47|28226|Bachelors Degree|Single|Education: Teacher||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502247579|502248010|31|0|2|502681447|31|0|2|500575685|10|2|500003586||4|1|500000294, 500004640, 500004901|-2||-2|0|10|||2238|7|||1|500000294, 500004640, 500004901|5493246288421413675|0
M465|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|187|Green||2015-07-30|2015-07-30|2016-02-02|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||6.1||1|1|1|1|M|Black||15|No|Mother|28215|7|One Parent: Female|$60,000 to $74,999||||No||School|General Community||Match Support|M|Black||52|28273|Bachelors Degree|Single|Self-Employed, Entrepreneur||25|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|501401583|501401868|31|0|1|504338671|31|0|1|500834950|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1||1421169092898167719|3003539216843226222
M466|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1421|Yellow|Amachi|2013-04-01|2013-04-16|NaT||||46.7||1|1|1|1|F|Black||15|Yes|Mother|28216|7|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||31|28262|Bachelors Degree|Single|Finance|28281|5|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502051702|501977740|31|0|2|503378835|31|0|2|500690864|10|2|-2||2|2|500000294|-2||-2|0|10|||7464|9|||1|500000294|1653226628427425023|0
M467|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|247|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-11-30|2016-08-03|Child/Family: Moved|Child/Family: Moved||8.1||1|1|2|2|F|Black||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||65|28205|Masters Degree|Divorced|Business|28255|40|5|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500017786|504425918|504428173|31|0|2|504383897|1|0|2|500851857|10|1|500014504||4|1|500014505, 500015184|-1|500014505, 500016394|-1|0|4|||46|2|||1|500014505, 500015184|702163000107564368|0
M468|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|36|Green||2015-01-26|2015-01-28|2015-03-05|Child: Lost interest|Child: Lost interest||1.2||1|1|1|1|F|Black||15|No|Mother|28273|8|One Parent: Male|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|Black||37|28273|Masters Degree|Single|Business|29715|3|0|Current/Previous Big|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500013781|504174131|504143662|31|0|2|503997551|31|0|2|500810212|10|2|-2||4|1||-2||-2|0|4|||17159|12|||1||194235582162093094|0
M469|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|255|Green||2015-10-16|2015-10-30|2016-07-11|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||8.4||1|1|1|1|M|Black||15|No|Mother|28208|8|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|M|White||38|28173|Bachelors Degree|Married|Finance|28217|0|2|Recruitment Event|BBBS Board/Staff|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504416061|504418313|31|0|1|504465459|1|0|1|500848780|10|1|500009132|2128207319|4|1||-1||-1|0|4|||7462|13|||1||3935539763241716148|0
M470|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3056|Green|Amachi|2008-08-21|2008-10-24|NaT||||100.4||1|1|2|2|M|Black||15|Yes|Mother|28230|10|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||37|28203|Masters Degree|Single|Medical: Doctor, Provider|28211|6|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501253195|501253471|31|0|1|500395148|1|0|1|500282924|10|2|500003586||2|1||-2||-2|0|10|||7464|9|||1|500000294|0|0
M471|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|441|Red|PERL 2014-2016|2015-11-30|2015-12-15|2017-02-28|Volunteer: Time constraint|Volunteer: Time constraint||14.5||1|1|1|1|M|Black||15||Mother|28209|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||31|28207|Masters Degree|Married|Finance: Accountant|28202|7|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020753|504289347|504291548|31|0|1|504428167|1|0|1|500863609|10|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|500014681|4440360203097874486|7044657180546140448
M472|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|120|Green||2016-10-30|2016-10-31|2017-02-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.9||2|3|2|3|F|Black||15|No|Mother|28217|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016, PERL 2014-2016|Match Support|F|Black||29|28209||Single|Customer Service|28217|0|6|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500022907|504416147|504418399|31|0|2|504212639|31|0|2|500921518|10|1|500014504||4|1|500014505, 500014681, 500016394|-1|500014505, 500016394|-1|0|4|||17159|12|||1||702163000107564368|0
M473|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|448|Green||2013-11-27|2013-12-19|2015-03-12|Child/Family: Moved|Child/Family: Moved||14.7||1|1|1|1|F|Black||15|No|Mother|2649|8|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||31|28203|Doctor of Medicine (MD)|Living w/ Significant Other|Medical|28112|1|2|other|College Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500015820|503569117|503570990|31|0|2|503583743|1|0|2|500735247|10|2|-2||4|1||-2||-2|0|10|||7670|5|||1||4440360203097874486|7674215580094440446
M474|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|272|Green|mentor2.0, mentor2.0 2015|2015-10-23|2015-11-05|2016-08-03|Child: Lost interest|Child: Lost interest||8.9||1|1|2|2|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|Black||23|28117|Bachelors Degree|Single|Business|28117|0|3|Duke Energy|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500017786|504454572|504456830|31|0|2|504359810|31|0|2|500851404|10|1|500014504||4|1|500015184|-1|500014505, 500016394|-1|0|4|||16705|3|||1|500014505, 500015184|702163000107564368|0
M475|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-11-17|NaT||||15.6||4|4|2|2|F|Black||15|Yes|Mother|28208|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||48|28211|Bachelors Degree|Single|Consultant|28278|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|502549826|502550279|31|0|2|501223094|31|0|2|500851882|10|1|500014504||2|1|500014505, 500015184|-1|500014505, 500015184|-1|0|4|||7462|13|||1|500014505, 500015184|3935539763241716148|0
M476|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1379|Green||2013-04-19|2013-05-28|NaT||||45.3||4|4|1|1|F|Black||15|Yes|Mother|28208|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||38|28215|Bachelors Degree|Single|Business: Mgt, Admin|28210|11|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502549826|502550279|31|0|2|503431300|31|0|2|500693780|10|2|-2||3|1|500014505, 500015184|-1||-2|0|4|||7464|9|||1||3935539763241716148|0
M477|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|572|Green||2014-11-07|2014-11-13|2016-06-07|Child: Changed school/site|Child: Changed school/site||18.8||4|4|2|2|F|Black||15|Yes|Mother|28208|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||31|28216|Masters Degree|Single|Customer Service|28217|1|6|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|502549826|502550279|31|0|2|504037091|31|0|2|500793483|10|1|500009132|2128207319|4|1|500014505, 500015184|-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M478|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|523|Green||2014-08-13|2014-08-21|2016-01-26|Volunteer: Time constraint|Volunteer: Time constraint||17.2||1|1|1|1|M|Black||15|No|Mother|28227|8|One Parent: Female|$60,000 to $74,999||||No|AARTF|BBBS Board/Staff|General Community||Match Support|M|Black||23|28227|Some College|Single|Student: College|28078|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503831166|503833145|31|0|1|503861120|31|0|1|500772203|10|2|-2||4|1||-2||-2|7294|13|||7496|10|||1||8202428416367135871|0
M479|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|593|Green||2015-07-23|2015-07-23|NaT||||19.5||1|1|1|1|M|Black||15|No|Mother|28215|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|White||31|28202|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504220177|504222291|31|0|1|504309758|1|0|1|500834242|10|2|-2||2|1||-2||-2|0|4|||46|2|||1||0|2876415545463317777
M480|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|861|Green|PERL 2014-2016|2014-10-15|2014-10-28|NaT||||28.3||2|2|1|1|F|Black||15|No|Mother|28208|8|One Parent: Female|Unknown||||No||School|General Community|PERL 2014-2016, Project Big|Match Support|F|Black||50|28278|Bachelors Degree|Single|Finance: Banking|29715|15|2|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020752|502699353|502700198|31|0|2|503945609|31|0|2|500783805|10|2|-2||2|1|500004640, 500014681|-2|500000294, 500014681|-2|0|4|||7496|10|||1|500014681|9076057728106637014|0
M481|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1408|Yellow||2012-10-04|2012-10-22|2016-08-30|Child/Family: Moved|Child/Family: Moved||46.3||2|2|1|1|M|Black||15|No|Mother|28273|3|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28273|Juris Doctorate (JD)|Single|Law: Lawyer||0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|501989028|502425720|31|0|1|503039778|31|0|1|500641725|10|2|-2||4|2|500005291|-2||-2|6855|8|||7496|10|635|1|1||0|0
M482|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-11-17|NaT||||15.6||1|1|1|1|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||Relative|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||36|28081|Bachelors Degree|Living w/ Significant Other|Business|28078|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504425672|504427927|31|0|2|504448500|1|0|2|500851858|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|3|||7462|13|||1|500014505, 500015184|702163000107564368|0
M483|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1376|Green||2013-04-15|2013-05-31|NaT||||45.2||1|1|1|1|M|Black||15|No|Mother|28269|9|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||33|28278|Bachelors Degree|Single|Arts, Entertainment, Sports|28269|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503023832|503025372|31|0|1|503139766|1|0|1|500692957|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1||1652521212990559348|3006000722566969828
M484|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|225|Yellow||2014-10-27|2014-11-17|2015-06-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.4||1|1|2|2|M|Black||15|Yes|Mother|28269|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|Hispanic||31|28209|High School Graduate|Single|Finance|28262|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503831971|503833950|31|0|1|504011759|3|0|1|500788190|10|2|-2||4|2|500000294|-2||-2|0|10|||46|2|||1||3677730851176818072|0
M485|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2118|Red||2010-10-28|2010-11-08|2016-08-26|Volunteer: Moved|Volunteer: Moved||69.6||1|1|1|1|M|Hispanic||15||Mother|28212|3|One Parent: Female|Unknown||||No|Spanish Radio|Media|General Community||Match Support|M|White||33|28226|Bachelors Degree|Single|Education: Teacher||3|0|Spanish Print|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502255225|502255655|3|0|1|502312682|1|0|1|500487118|10|2|-2||4|3||-2||-2|7068|1|||11662|1|||1||0|0
M486|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|354|Green|mentor2.0, mentor2.0 2015|2015-10-12|2015-10-26|2016-10-14|Volunteer: Time constraint|Volunteer: Time constraint||11.6||1|1|1|1|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|F|Black||40|28269|PHD|Single|Human Services: Psychologist|28027|4|1|BBBS National Site|Web Link|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500021786|504440275|504442531|31|0|2|504342087|31|0|2|500846705|10|1|500014504||4|1|500015184|-1|500015184|-1|0|4|||46|2|||1|500014505, 500015184|702163000107564368|0
M487|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|266|Green|PERL 2014-2016|2014-09-15|2014-09-25|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||2|2|1|1|M|Black||15|No|Mother|28206|6|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|M|White||25|28270|Bachelors Degree|Single|Finance|28202|0|1|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|501904523|500909693|31|0|1|503979230|1|0|1|500776009|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||16705|3|||1|500014681|7960300212314874874|0
M488|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1245|Red||2012-03-28|2012-04-19|2015-09-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||40.9||1|1|1|1|M|Black||15|No|Mother|28202|4|One Parent: Male|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28277||Single|Business||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502845758|502847118|31|0|1|502944923|1|0|1|500606912|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1||4726905079488957916|8858586900346693884
M489|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green|mentor2.0, mentor2.0 2015|2015-10-23|2015-11-11|NaT||||15.8||1|1|1|1|F|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||24|28202|Bachelors Degree|Single|Business|28202|0|2|BBBS National Site|Web Link|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454594|504456852|31|0|2|504249944|1|0|2|500851409|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||46|2|||1|500014505, 500015184|702163000107564368|0
M490|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2554|Green|Cabarrus County|2010-02-23|2010-03-10|NaT||||83.9||1|1|1|1|F|Black||15|No|Mother|28027|9|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||60|28213||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|501811395|501811730|31|0|2|500876892|31|0|2|500436702|10|2|500016307||2|1|500016374|-2|500016374|-2|6854|8|||2238|7|||1|500016374|370020301266015142|0
M491|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-10-26|NaT||||16.4||1|1|1|1|M|Hispanic||15|No|Mother|28210|9|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||28|28207|Bachelors Degree|Single|Business|28224|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504440268|504442524|3|0|1|504315884|1|0|1|500846213|10|1|500014504||2|1||-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M492|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Inactive|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||1|1|2|2|M|Multi-race (Black & Hispanic)||15|No|Mother|28217||One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||34|28210|Bachelors Degree|Married|Medical||3|6|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831598|504834100|38|0|1|504431507|1|0|1|500921878|10|1|500014504||3|1|500014505, 500016394|-1|500016394|-1|0|4|||7462|13|||1||702163000107564368|0
M493|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2669|Green|Amachi|2009-09-11|2009-09-29|2017-01-19|Child: Severity of challenges|Child: Severity of challenges||87.7||1|1|1|1|M|Black||15|Yes|GrandMother|28213|3|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||46|28227|High School Graduate|Single|Medical: Healthcare Worker|28269|4|0|Coworker|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500020752|501332658|501332937|31|0|1|501814288|1|0|1|500384166|10|2|-2||4|1|500000294|-2||-2|6854|8|||7447|3|||1|500000294|0|0
M494|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2118|Green|2010-2012 OJJDP JJI|2011-04-19|2011-05-20|NaT||||69.6||1|1|1|1|M|White||15|No|Mother|28226|9|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||55|28210|Bachelors Degree|Married|Finance|28203|1|6|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|1|0|0|1|277|60|598|500000170|500018851|502495501|502495950|1|0|1|502508181|1|0|1|500531873|10|2|-2||2|1|500005291|-2|500005291|-2|0|10|||7464|9|||1|500005291|1227369534771287213|0
M495|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|845|Green||2014-10-13|2014-11-13|NaT||||27.8||1|1|1|1|M|Black||15|No|Mother|28208|10|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Some Other Race||33|28056|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28204|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503803718|503805695|31|0|1|503930530|41|0|1|500783205|10|2|-2||2|1||-2||-2|34|2|||46|2|||1||6381341368426079638|6993050796559809579
M496|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1152|Yellow|Amachi|2012-12-11|2012-12-15|2016-02-10|Volunteer: Time constraint|Volunteer: Time constraint||37.8||1|1|1|1|M|Black||15|Yes|Mother|28205|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Amachi|Match Support|M|White||27|28203|Bachelors Degree|Single|Business||0|2|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|502983808|502985262|31|0|1|503140432|1|0|1|500668771|10|2|-2||4|2|500000294|-2|500000294|-2|0|4|||7464|9|||1|500000294|976372749760822282|3351268171347533976
M497|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|65|Green||2015-10-16|2015-10-31|2016-01-04|Volunteer: Time constraint|Volunteer: Time constraint||2.1||2|2|2|2|M|Black||15|No|Mother|28208|8|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||58|29715||Widowed|Business|28217|0|6|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504416042|504418294|31|0|1|504072039|1|0|2|500848785|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M498|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|168|Green||2016-01-04|2016-01-25|2016-07-11|Child: Changed school/site|Child: Changed school/site||5.5||2|2|2|2|M|Black||15|No|Mother|28208|8|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|M|White||40|28273||Married|Finance|28217|10|0|LPL Financial|Workplace Partner|Big|General Site|VOL - PreMatch|Match Support|0|1|1|0|277|60|598|500000170|500015820|504416042|504418294|31|0|1|504557665|1|0|1|500870050|10|1|500009132|2128207319|4|1||-1|500007920|-1|0|4|||11247|3|||1||3935539763241716148|0
M499|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1603|Yellow||2012-09-26|2012-10-16|NaT||||52.7||1|1|1|1|M|Black||15|No|Mother|28214|9|One Parent: Female|$45,000 to $49,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28207|Masters Degree|Married|Finance|28273|1|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503041998|503043639|31|0|1|503110820|1|0|1|500638908|10|2|-2||2|2||-2||-2|34|2|||7464|9|||1||216500609169513656|3962350215736335346
M500|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1042|Green||2014-04-23|2014-04-30|NaT||||34.2||1|1|2|2|F|Black||15|No|Mother|28214|9|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||45|28227|Bachelors Degree|Married|Customer Service|28262|18|0|Big For A Day|Special Event|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|502146600|502932575|31|0|2|503483337|31|0|2|500760757|10|2|-2||2|1||-2|500000294|-2|6854|8|||16422|8|||1||8029775806705219538|0
M501|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1996|Green|2010-2012 OJJDP JJI|2011-09-15|2011-09-19|NaT||||65.6||2|2|1|1|M|Black||15|No|Mother|28213|5|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28213|Bachelors Degree|Married|Tech: Support, Writing|28273|11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|501604446|501604760|31|0|1|502664359|31|0|1|500555050|10|2|-2||2|1|500005291|-2||-2|0|10|||7462|13|||1|500005291|4013586283864837776|0
M502|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|287|Yellow|mentor2.0, mentor2.0 2015|2015-10-12|2015-10-26|2016-08-08|Child: Lost interest|Child: Lost interest||9.4||1|1|3|3|M|Black||15|No|Father|28217|9|One Parent: Male|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|M|Black||32|28216|Masters Degree|Single|Finance: Accountant|28280|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014, mentor2.0 2016|Match Support|0|1|1|0|277|60|598|500000170|500021786|504451288|504453544|31|0|1|503976447|31|0|1|500846708|10|1|500014504||4|2|500015184|-1|500014505, 500014506, 500016394|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M503|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|579|Green||2013-10-18|2013-11-15|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19||1|1|2|2|F|Asian||15|No|Father|28206|6|Two Parent|Unknown|||Y|Yes||School|General Community||Enrollment|F|White||29|28031|Masters Degree|Married|Tech: Support, Writing|28202|2|5|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503635399|504018995|4|0|2|503605621|1|0|2|500720718|5|1|500009132|2128173561|4|1||-2|500014681|-1|0|4|||16705|3|||1||7960300212314874874|0
M504|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|247|Red|PERL 2014-2016|2014-12-08|2015-01-12|2015-09-16|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||8.1||5|5|1|1|M|Black||15|No|Mother|28203|7|One Parent: Female|$15,000 to $19,999||||Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||22|28210|Some College|Single|Customer Service|28208|0|1|Man Up Campaign|Media|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500008321|501068963|501069236|31|0|1|503906067|31|0|1|500801900|10|2|-2||4|3|500014681|-2|500014681|-2|0|4|||17101|1|||1|500014681|8568001799025358453|7044657180546140448
M505|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|456|Red||2015-06-18|2015-06-29|2016-09-27|Child/Family: Time constraints|Child/Family: Time constraints||15||2|2|1|1|F|Some Other Race||15|No|Aunt|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||36|28210|Masters Degree|Single|Finance: Accountant|28202|6|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502612404|500188044|41|0|2|504226710|1|0|2|500830721|10|2|-2||4|3||-2||-2|0|10|||17159|12|||1||1421169092898167719|6156547733130613405
M506|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|233|Red|PERL 2014-2016|2014-08-28|2014-10-06|2015-05-27|Volunteer: Moved|Volunteer: Moved||7.7||2|2|1|1|F|Some Other Race||15|No|Aunt|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||26|28217|Bachelors Degree|Single|Business|28277|0|8|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500013781|502612404|500188044|41|0|2|503790988|31|0|2|500773744|10|2|-2||4|3||-2|500014681|-2|0|10|||46|2|||1|500014681|1421169092898167719|6156547733130613405
M507|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1469|Green||2013-02-25|2013-02-27|NaT||||48.3||1|1|1|1|M|Black||15|No|Mother|28212|7|Two Parent|$35,000 to $39,999|Yes: Active|Yes||No||Relative|General Community||Match Support|M|White||30|28105|Bachelors Degree|Single|Business: Sales|17001|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502663937|502664764|31|0|1|503296990|1|0|1|500684232|10|2|-2||2|1||-2||-2|0|3|||7496|10|||1||0|0
M508|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|476|Green|mentor2.0, mentor2.0 2015|2015-10-09|2015-11-17|NaT||||15.6||1|1|1|1|M|Black||15|No|Mother|28217|10|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||30|28209|Masters Degree|Single|Business: Engineer|28202|7|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454656|504456914|31|0|1|504387544|1|0|1|500846233|10|1|500014504||2|1||-1|500014505, 500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M509|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|275|Green||2016-05-10|2016-05-24|2017-02-23|Volunteer: Moved|Volunteer: Moved||9||1|1|1|1|M|Black||15|No|Mother|28208|9|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|PHD|Single|Self-Employed, Entrepreneur|30604|4|0|Local Print|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020910|504347348|504349572|31|0|1|504566830|1|0|1|500892524|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|34|2|||7439|1|||1||2374609189072499123|7044657180546140448
M510|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green|mentor2.0, mentor2.0 2015|2015-10-25|2015-11-11|NaT||||15.8||1|1|1|1|M|Black||15|No|Mother|28208|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|M|White||28|28269||Married|Business: Engineer|28078|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454566|504456824|31|0|1|504448602|1|0|1|500851873|10|1|500014504||2|1|500014505, 500015184|-1|500015184|-1|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M511|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2231|Green||2009-06-01|2009-06-24|2015-08-03|Volunteer: Time constraint|Volunteer: Time constraint||73.3||1|1|1|1|M|Black||15|No|Mother|28269|8|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Multi-race (Asian & White)||34|28205|Bachelors Degree|Single|Tech: Research/Design|28255|3|1|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500011349|501641325|501641648|31|0|1|501715652|37|0|1|500366872|10|2|-2||4|1|500000294|-2|500000294|-2|6854|8|||7464|9|||1||9134125726462845918|7124320636013019662
M512|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|392|Red||2014-08-27|2014-09-15|2015-10-12|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12.9||2|2|1|1|M|Black||15|No|Mother|28215|2|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||40|28217|Masters Degree|Single|Finance: Accountant|28034|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|501627668|501627988|31|0|1|503921388|1|0|1|500773645|10|2|-2||4|3||-2||-2|0|10|||17159|12|||1||0|4715213876709649683
M513|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2113|Green|Amachi|2011-05-18|2011-05-25|NaT||||69.4||2|2|1|1|F|Black||15|Yes|Mother|28212|3|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||34|28203|Masters Degree|Single|Business: Mgt, Admin|28273|0|7|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502270499|502231230|31|0|2|502510107|1|0|2|500536754|10|2|500003586||2|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294|0|0
M514|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1220|Green||2013-09-10|2013-10-22|2017-02-23|Volunteer: Time constraint|Volunteer: Time constraint||40.1||2|2|1|1|M|Black||15|No|Mother|28215|7|One Parent: Female|Less than $10,000||||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|White||41|28269|Bachelors Degree|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501010684|503560069|31|0|1|503491643|1|0|1|500710107|10|2|-2||4|1|500005291|-2||-2|7016|11|||7464|9|||1||6724463016047116758|1786514887916898235
M515|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1888|Green||2010-10-11|2010-10-20|2015-12-21|Child/Family: Moved|Child/Family: Moved||62||2|2|1|1|F|Black||15|No|Mother|28227|1|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||48|28210|Some College|Single|Human Services||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501123191|500915629|31|0|2|502153920|1|0|2|500478644|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||0|0
M516|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|49|Green|mentor2.0, mentor2.0 2016|2017-01-05|2017-01-17|NaT||||1.6||1|1|2|2|F|Black||15|No|Mother|28208|9|Two Parent|$20,000 to $24,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||25|28203|Bachelors Degree|Single|Business|28201|1|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831621|504834123|31|0|2|504357339|1|0|2|500938318|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500015184, 500016394|-1|0|4|||7462|13|||1|500014505, 500016394|702163000107564368|6960968151966841272
M517|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|449|Green|Amachi, PERL 2014-2016|2015-11-20|2015-12-14|NaT||||14.8||1|1|1|1|F|Black||15|Yes|Mother|28215|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi, PERL 2014-2016|Match Support|F|White||30|28203|Bachelors Degree|Single|Business|60611|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|503611732|503613600|31|0|2|504421910|1|0|2|500862006|10|2|-2||2|1|500000294, 500014681|-2|500014681|-2|0|10|||17159|12|||1|500000294, 500014681|6724463016047116758|0
M518|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|924|Red||2013-11-13|2013-11-26|2016-06-07|Child: Changed school/site|Child: Changed school/site||30.4||1|1|2|2|F|Hispanic||15|No|Mother|28202|7|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Asian||38|28215|Some College|Married|Finance|28217|5|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|503681630|503683595|3|0|2|503162750|4|0|2|500730752|10|1|500009132|2128207319|4|3||-1||-1|0|4|||11247|3|1204|3|1||3935539763241716148|0
M519|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green||2016-11-18|2016-11-28|NaT||||3.3||1|1|2|2|F|Black||15|Yes|Mother|28217|9|One Parent: Female|Less than $10,000||||Yes||School|General Site|mentor2.0|Match Support|F|Black||23|28117|Bachelors Degree|Single|Business|28117|0|3|Duke Energy|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831552|504834054|31|0|2|504359810|31|0|2|500929516|10|1|500014504||2|1|500014505|-1|500014505, 500016394|-1|0|4|||16705|3|||1||702163000107564368|0
M520|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2259|Green|Amachi, Project Big, Project Big AND Amachi|2010-12-13|2010-12-30|NaT||||74.2|Y|2|2|2|2|M|Black||15|Yes|Mother|28216|7|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|502180724|502181148|31|0|1|502391505|31|0|2|500505039|10|2|500004772||2|1|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7438|1|||1|500000294, 500004640, 500004901|46835895261850668|0
M521|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|826|Red||2013-09-09|2013-10-01|2016-01-05|Volunteer: Time constraint|Volunteer: Time constraint||27.1||2|2|1|1|M|Black||15|No|Mother|28216|9|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community||Match Support|M|Black||32|28277|Bachelors Degree|Single|Construction|28211|0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500784687|500784955|31|0|1|503531111|31|0|1|500709609|10|2|-2||4|3||-2||-2|0|5|||7464|9|||1||0|1786514887916898235
M522|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|532|Green|PERL 2014-2016|2015-02-20|2015-03-17|2016-08-30|Volunteer: Moved|Volunteer: Moved||17.5||2|2|1|1|M|Black||15||GrandMother|28227|3|One Parent: Female|Unknown|||Y|Yes|AARTF|BBBS Board/Staff|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||25|28202|Bachelors Degree|Single|Finance: Banking|28202|0|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500018851|502287066|502287498|31|0|1|504056150|1|0|1|500814738|5|2|-2||4|1|500005291|-2|500014681|-2|7294|13|||17159|12|||1|500014681|0|0
M523|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|58|Green||2017-01-06|2017-01-08|NaT||||1.9||1|1|2|2|M|Black||15|No|Father|28208|8|Two Parent: Not Married|Unknown||||Yes||School|General Site||Match Support|M|White||23|28202|Bachelors Degree|Single|Business|28202|0|9|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504976123|504978668|31|0|1|504685043|1|0|1|500938699|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M524|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|372|Green|PERL 2014-2016|2016-02-18|2016-02-29|NaT||||12.2||1|1|1|1|M|Black||15|No|Mother|28209|7|One Parent: Female|$25,000 to $29,999||||Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||29|28209|Masters Degree|Single|Law: Lawyer|28202|0|4|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|500917189|500917459|31|0|1|504538036|1|0|1|500880191|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||7464|9|||1|500014681|7276767778509034039|2719955880210213907
M525|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|280|Green||2016-05-16|2016-05-31|NaT||||9.2||1|1|1|1|F|Black||15|No|Mother|28212|8|One Parent: Female|$40,000 to $44,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||48|28212|Associate Degree|Single|Finance||11|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504473782|504476056|31|0|2|504550297|1|0|2|500893115|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1||8202428416367135871|2806833304218536184
M526|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-11|2016-11-02|NaT||||4.1||1|1|1|1|F|Hispanic||15|No|Mother|28217|9|Two Parent|$10,000 to $14,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||36|28269|Juris Doctorate (JD)|Single|Finance|28262|1|0|Self|Self|Big|General Site|mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504834787|504837289|3|0|2|504808345|31|0|2|500914305|10|1|500014504||2|1|500014505, 500016394|-1|500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M527|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|76|Green||2016-12-05|2016-12-21|NaT||||2.5||1|1|1|1|M|Black||15|No|Mother|28227|8|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||25|28277|Bachelors Degree|Single|Business|28208|1|8|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504662357|504664784|31|0|1|504791469|31|0|1|500933117|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1||7883015200677941272|3557919386369667257
M528|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1329|Green||2013-06-12|2013-07-17|NaT||||43.7||1|1|1|1|F|Black||15|No|Mother|28215|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|Black||39|28214|Bachelors Degree|Single|Govt||1|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|503230648|502841119|31|0|2|503169561|31|0|2|500700323|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||0|3714886275549507192
M529|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2475|Green||2010-05-03|2010-05-28|NaT||||81.3||1|1|1|1|M|Black||15|No|Mother|28262|7|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black|Other African|32|28262||Married|Law: Police Officer||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501611456|501611776|31|0|1|501876475|31|31|1|500450969|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||806697982905023857|4701122331973296331
M530|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|165|Red|PERL 2014-2016|2015-04-16|2015-04-27|2015-10-09|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||5.4||2|2|2|2|F|Black||15|No|Mother|28262|8|One Parent: Female|$45,000 to $49,999||||No||School|General Community|PERL 2014-2016|Match Support|F|Black||38|28269|Masters Degree|Single|Business|28262|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500017777|503974135|503598965|31|0|2|503860995|31|0|2|500823546|10|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|500014681|1320477920662455183|1198499568025045356
M531|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|312|Green||2016-03-14|2016-04-29|NaT||||10.3||2|2|1|1|F|Black||15|No|Mother|28262|8|One Parent: Female|$45,000 to $49,999||||No||School|General Community|PERL 2014-2016|Match Support|F|Black||20|28213||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503974135|503598965|31|0|2|504341793|31|0|2|500884595|10|2|-2||2|1|500014681|-2||-2|0|4|||46|2|||1||1320477920662455183|1198499568025045356
M532|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-31|2016-11-02|NaT||||4.1||1|1|1|1|F|Black||15|No|Mother|28217|9|Two Parent|$10,000 to $14,999|||Y|Yes||Relative|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||38|28269|Masters Degree|Single|Business: Mgt, Admin|28213|2|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504842890|504845392|31|0|2|504780315|31|0|2|500921750|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|3|||7464|9|||1||702163000107564368|5081726734274569781
M533|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1141|Green|Amachi|2013-03-27|2013-04-10|2016-05-25|Volunteer: Moved|Volunteer: Moved||37.5||1|1|1|1|M|Black||15|No|Mother|28212|5|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||27|28209|Bachelors Degree|Single|Finance|28255|1|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|503246887|503248691|31|0|1|503253208|1|0|1|500690197|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||46|2|||1|500000294|2762897743412756173|0
M534|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|488|Green|mentor2.0 2015|2015-10-25|2015-11-05|NaT||||16||1|1|1|1|M|Hispanic||15|Yes|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0 2015|Match Support|M|Hispanic||32|28273||Married|Customer Service|28037|0|1|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504454583|504456841|3|0|1|504274695|3|0|1|500851871|10|1|500014504||2|1|500015184|-1|500015184|-1|0|4|||17159|12|||1|500015184|702163000107564368|0
M535|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-26|2016-11-04|NaT||||4||1|1|2|2|F|Black||15|No|Mother|28208|9|One Parent: Female|$10,000 to $14,999||||Yes||Relative|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||35|28213|Masters Degree|Single|Business||4|0|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504842854|504845356|31|0|2|500953330|31|0|2|500920220|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|3|||46|2|||1||702163000107564368|8696376245285900472
M536|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|326|Green||2014-11-07|2014-11-07|2015-09-29|Child: Changed school/site|Child: Changed school/site||10.7||1|1|2|2|F|Black||15|No|Mother|28217|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||58|29715||Widowed|Business|28217|0|6|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|504089143|504091173|31|0|2|504072039|1|0|2|500793456|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M537|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1269|Yellow||2012-10-01|2012-10-31|2016-04-22|Child/Family: Moved|Child/Family: Moved||41.7||2|2|2|2|M|Black||15|No|Mother|28215|1|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|M|White||31|28269|Masters Degree|Single|Insurance|28262|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501372080|501372359|31|0|1|502500246|1|0|1|500640327|10|2|-2||4|2||-2||-2|0|3|||7496|10|||1||314687390558932914|8166272525880133677
M538|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|445|Yellow||2014-11-07|2014-11-13|2016-02-01|Child/Family: Moved|Child/Family: Moved||14.6||1|1|1|1|M|Black||15|No|Father|28217|8|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|M|White||22|28270|Masters Degree|Married|Business|28217|3|3|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|504089098|504091128|31|0|1|504037139|1|0|1|500793480|10|1|500009132|2128207319|4|2||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M539|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2769|Green||2009-07-22|2009-08-07|NaT||||91||1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28216|5|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||49|28031|Bachelors Degree|Married|Transport: Pilot|40223|9|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|501809541|501809896|36|0|1|501620528|1|0|1|500375025|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||0|0
M540|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|784|Yellow|PERL 2014-2016|2015-01-09|2015-01-13|NaT||||25.8||1|1|1|1|F|Black||15|Yes|Mother|28212|9|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||25|28213|Bachelors Degree|Single|Retail: Mgt||0|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504076406|504078432|31|0|2|503831499|31|0|2|500807374|10|2|-2||2|2|500014681|-2|500014681|-2|0|5|||17159|12|||1|500014681|3292090474897428830|7044657180546140448
M541|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|403|Green|mentor2.0, mentor2.0 2016|2016-01-04|2016-01-29|NaT||||13.2||2|2|2|2|F|Black||15|Yes|Mother|28208|9|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||50|28262||Married|Business: Sales|28217|5|5|LPL Financial|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504416180|504418432|31|0|2|503630789|31|0|2|500870097|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||11247|3|||1|500014505, 500016394|702163000107564368|0
M542|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|65|Yellow||2015-10-16|2015-10-31|2016-01-04|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||2.1||2|2|1|1|F|Black||15|Yes|Mother|28208|9|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||40|28210|Bachelors Degree|Married|Consultant|28217|0|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504416180|504418432|31|0|2|504399592|31|0|2|500848805|10|1|500009132|2128207319|4|2|500014505, 500016394|-1||-1|0|4|||11247|3|||1||702163000107564368|0
M543|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-26|2016-11-02|NaT||||4.1||1|1|1|1|M|Multi-race (Asian & White)||15|No|Mother|28217|9|One Parent: Female|Less than $10,000||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||31|28217|Bachelors Degree|Married|Business|28278|3|0|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504834756|504837258|37|0|1|504767391|1|0|1|500920166|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||46|2|||1||702163000107564368|3677141092383031375
M544|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1532|Green|2010-2012 OJJDP JJI|2011-07-25|2011-08-03|2015-10-13|Volunteer: Time constraint|Volunteer: Time constraint||50.3||1|1|1|1|M|Black||15||GrandMother|28227|3|Grandparents|Unknown||||No||Self|General Community|PERL 2014-2016|RTBM|M|White||27|28205|Associate Degree|Single|Law: Police Officer||0|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|1|0|1|0|277|60|598|500000170|500017777|502252828|502253254|31|0|1|502602451|1|0|1|500547383|7|2|-2||4|1|500014681|-2|500005291|-2|0|10|||7496|10|||1|500005291|0|0
M545|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|293|Green||2015-09-16|2015-10-08|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.6||1|1|2|2|M|Black||15|Yes|Mother|28208|7|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site||Match Support|M|Black||48|28205|Masters Degree|Single|Finance|28202|3|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504423117|504425370|31|0|1|504359583|31|0|1|500840442|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M546|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2533|Red|Cabarrus County|2010-02-18|2010-03-02|2017-02-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||83.2||1|1|1|1|M|Black||15|No|Mother|28083||One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||52|28075||Married|Medical: Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500022817|501716720|501716992|31|0|1|501878786|31|0|1|500435676|10|2|500016307||4|3|500016374|-2|500016374|-2|6854|8|||7464|9|||1|500016374|0|0
M547|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|578|Yellow|Amachi|2014-05-14|2014-05-22|2015-12-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||19||1|1|2|2|M|Black||15|Yes|Mother|28227|7|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||30|28213|Masters Degree|Single|Education|28217|0|7|Recruitment Event|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500018851|503728057|503730029|31|0|1|503788318|31|0|1|500763247|10|2|-2||4|2||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7458|9|||1|500000294|5604470640552265812|7825731075480167876
M548|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-26|2016-11-04|NaT||||4||1|1|1|1|F|Black||15|No|Mother|28209|9|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||27|28215|Masters Degree|Single|Business||0|8|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831502|504834004|31|0|2|504775164|31|0|2|500920214|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||17159|12|||1||702163000107564368|0
M549|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|911|Green||2014-07-21|2014-07-30|2017-01-26|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||29.9||1|1|1|1|M|Black||15|No|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||38|28269|Some College|Married|Tech: Management|28273|3|1|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503899239|503901239|31|0|1|503871007|1|0|1|500770094|10|2|-2||4|1||-2||-2|0|10|||17101|1|||1||253338316288302752|7044657180546140448
M550|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|543|Green||2014-04-11|2014-04-24|2015-10-19|Volunteer: Moved|Volunteer: Moved||17.8||2|2|1|1|F|Multi-race (Black & White)||15|No|Mother|28134|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||55|28217|Some College|Married|Retail: Mgt|28217|14|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503722616|503724588|36|0|2|503707316|1|0|2|500759403|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||7872663507285703533|3402014428779854546
M551|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|374|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-22|2016-02-27|NaT||||12.3||2|2|1|1|F|Multi-race (Black & White)||15|No|Mother|28134|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||30|28226|Bachelors Degree|Single|Business|28202|4|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|503722616|503724588|36|0|2|504343006|31|0|2|500880706|10|2|-2||3|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|500007920, 500011315, 500011316|7872663507285703533|3402014428779854546
M552|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|266|Green|PERL 2014-2016|2014-09-18|2014-09-25|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||2|2|1|1|F|Black||15|No|Mother|28205|7|One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|F|White||31|28203|Bachelors Degree|Single|Consultant|28202|2|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|RTBM|1|0|1|0|277|60|598|500000170|500016270|503623969|503625858|31|0|2|503976684|1|0|2|500776599|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||16705|3|||1|500014681|7960300212314874874|0
M553|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|547|Green||2013-10-14|2013-11-18|2015-05-19|Child/Family: Moved|Child/Family: Moved||18||1|1|1|1|M|Black||15|No|Mother|28052|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||30|28216|Masters Degree|Married|Finance: Accountant|28202|2|7|Duke Energy|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503635425|503637375|31|0|1|503606058|1|0|1|500718999|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M554|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|129|Green||2016-09-16|2016-10-17|2017-02-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.2||1|1|1|1|M|Black||15|No|Mother|28211|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||34|28209||Married|Business: Sales||0|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020910|504039275|504041293|31|0|1|504461897|1|0|1|500908017|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||675142027733303647|0
M555|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|159|Green||2016-01-25|2016-02-03|2016-07-11|Child: Changed school/site|Child: Changed school/site||5.2||2|2|2|2|F|Black||15|No|Mother|28208|8|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|Black||44|28216|Bachelors Degree|Single|Business||2|0|LPL Financial|Workplace Partner|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500015820|504526221|504528553|31|0|2|504349689|31|0|2|500875232|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M556|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|49|Yellow||2015-11-17|2015-12-02|2016-01-20|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||1.6||2|2|1|1|F|Black||15|No|Mother|28208|8|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|Multi-race (Black & Hispanic)||33|28215|Bachelors Degree|Married|Consultant|28217|0|5|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504526221|504528553|31|0|2|504396970|38|0|2|500860672|10|1|500009132|2128207319|4|2||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M557|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|416|Green||2014-04-25|2014-04-28|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||13.7||2|2|1|1|F|Black||15|Yes|Mother|28205|6|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|Match Support|F|Black||43|28078|Masters Degree|Single|Business: Human Resources|28202|7|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503633871|503635812|31|0|2|503855574|31|0|2|500761186|10|1|500009132|2128173561|4|1|500000294|-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M558|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|48|Green||2015-02-02|2015-02-11|2015-03-31|Child/Family: Moved|Child/Family: Moved||1.6||2|2|1|1|F|Black||15|No|Mother|28208|9|Two Parent|$15,000 to $19,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||37|28120|Masters Degree|Married|Finance: Accountant|28202|12|0|Duke Energy|Workplace Partner|Big|General Site||Enrollment|0|1|1|0|277|60|598|500000170|500016270|504183446|504185555|31|0|2|503979203|1|0|2|500811396|10|1|500009132|2128173561|4|1|500014505, 500016394|-1||-1|0|4|||16705|3|||1||702163000107564368|0
M559|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-27|2016-11-04|NaT||||4||2|2|1|1|F|Black||15|No|Mother|28208|9|Two Parent|$15,000 to $19,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||26|28202|Bachelors Degree|Single|Business: Mgt, Admin|28226|2|9|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500022907|504183446|504185555|31|0|2|504267362|1|0|2|500920575|10|1|500014504||2|1|500014505, 500016394|-1|500015184|-1|0|4|||17159|12|||1||702163000107564368|0
M560|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|3100|Green||2008-05-05|2008-05-14|2016-11-08|Volunteer: Time constraint|Volunteer: Time constraint||101.8||1|1|1|1|M|White||15|No|Father|28025|4|One Parent: Male|Unknown||||No||Self|General Community|Cabarrus County|Enrollment|M|White||49|27103|Masters Degree|Single|Education: Teacher|27282|0|0|Other|Service Organization|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500020753|501247286|500341682|1|0|1|501247141|1|0|1|500264655|5|2|-2||4|1|500016374|-2|500016374|-2|0|10|||7452|6|||1||1345826867198613426|0
M561|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|523|Green|mentor2.0, mentor2.0 2016|2015-05-27|2015-05-27|2016-10-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||17.2||2|2|4|4|M|Black||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|Black||44|29732|High School Graduate|Married|Business|28217|5|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500022907|504312104|504314322|31|0|1|503754104|31|0|1|500828440|10|1|500009132|2128207319|4|1|500014505, 500016394|-1||-1|0|4|||11247|3|||1|500014505, 500016394|702163000107564368|0
M562|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||2|2|1|1|M|Black||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|Black||36|28203|Bachelors Degree|Single|Tech: Computer/Programmer|28202|10|11|TV|Media|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504312104|504314322|31|0|1|504766848|31|0|1|500921866|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||130|1|||1||702163000107564368|0
M563|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|98|Green||2016-11-08|2016-11-29|NaT||||3.2||1|1|1|1|F|Black||15|No|Mother|28211|9|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||47|28215|Masters Degree|Married|Education|28202|5|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504471621|504473895|31|0|2|504580592|31|0|2|500925801|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||7501346876523517480|1545381051186164660
M564|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|311|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-04-13|2016-04-30|NaT||||10.2||1|1|1|1|M|Black||15|No|Mother|28120|6|One Parent: Female|Less than $10,000||||Yes||Relative|General Community|PERL 2014-2016|Match Support|M|White||28|28214|Bachelors Degree|Married|Business|28214|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|503782093|503784070|31|0|1|504545677|1|0|1|500888935|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|3|||17159|12|||1|500007920, 500011315, 500011316|7872663507285703533|0
M565|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2931|Green|Amachi|2009-02-18|2009-02-26|NaT||||96.3||1|1|1|1|M|Black||15|Yes|Mother|28206|7|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Single|Tech: Computer/Programmer||0|5|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|501390344|501390617|31|0|1|501380163|1|0|1|500342682|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294|4863631750424600365|5161383151676749743
M566|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1764|Green|Amachi|2012-04-11|2012-05-08|NaT||||58||2|2|1|1|M|Black||15|Yes|Mother|28206|7|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||35|28206|Bachelors Degree|Single|Business: Sales|28117|4|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|501390345|501390617|31|0|1|502966998|1|0|1|500609269|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294|4863631750424600365|5161383151676749743
M567|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|628|Green|PERL 2014-2016|2015-06-10|2015-06-18|NaT||||20.6||1|1|1|1|F|Black||15|No|Mother|28212|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||31|28204|Masters Degree|Single|Student: College||0|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500017732|502979699|502981150|31|0|2|504127445|1|0|2|500829841|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||7464|9|||1|500014681|7883015200677941272|415738029281868742
M568|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|736|Green||2015-02-23|2015-03-02|NaT||||24.2||1|1|1|1|M|Black||15|No|Mother|28105|7|One Parent: Female|$40,000 to $44,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||45|28226|Bachelors Degree|Single|Insurance|28226|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503413167|503415024|31|0|1|504190868|1|0|1|500815087|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1||2129686509389594346|3714886275549507192
M569|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1504|Green||2012-07-18|2012-08-03|2016-09-15|Child/Family: Moved|Child/Family: Moved||49.4||1|1|1|1|M|Black||15|No|Mother|28205|4|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance: Banking|28202|0|7|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500020910|503044619|503046265|31|0|1|503021454|1|0|1|500624634|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1||5822146217251000296|7044657180546140448
M570|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|61|Green||2016-10-31|2016-11-04|2017-01-04|Child/Family: Moved|Child/Family: Moved||2||3|3|2|2|F|Black||15|Yes|GrandMother|28208|9|Grandparents|Unknown||||Yes||School|General Site|Amachi, mentor2.0, mentor2.0 2016|Match Support|F|Black||34|28262|Bachelors Degree|Single|Insurance|28277|0|4|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Enrollment|0|1|1|0|277|60|598|500000170|500022907|502821865|502823144|31|0|2|504267500|31|0|2|500921744|10|1|500014504||4|1|500000294, 500014505, 500016394|-1|500014505, 500016394|-1|0|4|||17159|12|||1||702163000107564368|0
M571|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|249|Green||2015-11-02|2015-11-05|2016-07-11|Child: Changed school/site|Child: Changed school/site||8.2||2|2|5|5|M|Black||15|No|Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||49|28278|Bachelors Degree|Separated|Finance|28217|7|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|503678239|503680204|31|0|1|500189616|31|0|1|500855262|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M572|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|721|Green||2013-11-11|2013-11-11|2015-11-02|Volunteer: Time constraint|Volunteer: Time constraint||23.7||2|2|1|1|M|Black||15|No|Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||39|28210|Masters Degree|Married|Finance|28217|6|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|503678239|503680204|31|0|1|503689039|1|0|1|500729623|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M573|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2716|Green|Amachi|2009-09-24|2009-09-29|NaT||||89.2||1|1|2|3|F|Black||15|Yes|Mother|28215|6|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||38|28273||Single|Tech: Engineer||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501831581|501831944|31|0|2|500715453|31|0|2|500387624|10|2|500003586||2|1|500000294|-2||-2|0|10|||46|2|||1|500000294|6724463016047116758|0
M574|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1619|Green||2012-08-17|2012-09-30|NaT||||53.2||1|1|1|1|M|Black||15|No|Mother|28216|8|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||28|28269|Some College|Single|Business: Clerical||0|3|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503071479|503069483|31|0|1|503051382|1|0|1|500629193|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1||7679812394383646966|7291948965517877884
M575|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-22|2015-10-01|NaT||||17.2||1|1|3|3|M|Black||15|Yes|Mother|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|White||29|28202|Bachelors Degree|Single|Business: Engineer|28202|5|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504410184|504412435|31|0|1|503979778|1|0|1|500841354|10|1|500009132|2128212899|2|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M576|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2377|Green||2010-08-12|2010-08-27|2017-02-28|Volunteer: Time constraint|Volunteer: Time constraint||78.1||2|2|1|1|F|Black||15|No|Mother|28216|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||30|28209|Bachelors Degree|Single|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501529924|501530213|31|0|2|502199360|1|0|2|500465517|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||0|0
M577|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|21|Yellow||2015-12-09|2015-12-18|2016-01-08|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||0.7||1|1|1|1|F|Black||15|No|Mother|28269|8|One Parent: Female|$30,000 to $34,999||||Yes||School|General Community|VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|F|White||26|28078|Masters Degree|Single|Business: Marketing|28269|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500017777|504458036|504460294|31|0|2|504416792|1|0|2|500866388|5|2|-2||4|2|500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||7276767778509034039|3086452374500817499
M578|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2107|Green|Amachi, 2010-2012 OJJDP JJI|2011-05-19|2011-05-31|NaT||||69.2||1|1|1|1|F|Black||15|Yes|Mother|28206|3|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||40|28269|Masters Degree|Single|Tech: Engineer|77058|6|6|Relative|Relative|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502569117|502569571|31|0|2|502538689|31|0|2|500536957|10|2|500003586||2|1|500005291|-2||-2|0|10|||17161|11|||1|500000294, 500005291|8979408036987322141|7106634858630667125
M579|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-26|2016-11-02|NaT||||4.1||1|1|1|1|F|Black||15|Yes|GrandMother|28217|9|Grandparents|$10,000 to $14,999||||Yes||School|General Site|Amachi, mentor2.0, mentor2.0 2016|Match Support|F|Black||38|29720|Bachelors Degree|Married|Business: Mgt, Admin|28209|14|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504859855|504834054|31|0|2|504784459|31|0|2|500920225|10|1|500014504||2|1|500000294, 500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M580|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|251|Yellow||2015-10-16|2015-11-03|2016-07-11|Child: Severity of challenges|Child: Severity of challenges||8.2||1|1|2|2|F|Black||15|No|Mother|28208|8|Two Parent|$15,000 to $19,999||||Yes||Relative|General Site||Match Support|F|Multi-Race (None of the above)||34|28134|Some College|Single|Business|28217|2|4|LPL Financial|Workplace Partner|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500015820|504416166|504418418|31|0|2|503799347|7|0|2|500848808|10|1|500009132|2128207319|4|2||-1||-1|0|3|||11247|3|||1||3935539763241716148|0
M581|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2994|Red|Cabarrus County|2008-11-26|2008-11-26|2017-02-06|Child: Severity of challenges|Child: Severity of challenges||98.4||3|3|1|1|F|White||15||Father|28025|1|One Parent: Male|Unknown||||No||School|General Site|Cabarrus County|Match Support|F|White||44|28037|Bachelors Degree|Married|Business: Sales|28027|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500022817|501536733|501537025|1|0|2|501418563|1|0|2|500320917|10|2|500016307||4|3|500016374|-1|500016374|-2|0|4|||7464|9|||1|500016374|0|1466298645186383139
M582|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-21|2016-10-31|NaT||||4.2||1|1|1|1|M|Black||15|No|Mother|28105|9|One Parent: Female|Less than $10,000|||Y|Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|Black||30|28105|Bachelors Degree|Married|Business|28078|0|7|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504698283|504700711|31|0|1|504765309|31|0|1|500918562|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|56|1|||7464|9|||1||0|7044657180546140448
M583|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2810|Green||2008-06-06|2008-06-23|2016-03-03|Child: Family structure changed|Child: Family structure changed||92.3|Y|1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28227|6|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||45|28211||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|501185592|501185866|36|0|1|501255830|1|0|1|500270254|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1||8452412398369747552|0
M584|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2709|Green||2009-08-19|2009-09-29|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||89||1|1|1|1|F|Black||15|No|Mother|28269|1|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||31|28262|Bachelors Degree|Single|Medical: Admin|28216|0|8|Recruitment Event|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501771263|501741899|31|0|2|501622704|31|0|2|500379993|10|2|-2||4|1||-2||-2|0|10|||7443|2|||1||0|0
M585|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-27|2016-11-04|NaT||||4||1|1|1|1|F|Multi-Race (None of the above)||15|No|Mother|28217|9|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||45|28269|Masters Degree|Married|Unknown|28206|0|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831667|504834169|7|0|2|504780301|31|0|2|500920538|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|4200792623487537971
M586|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-27|2016-11-04|NaT||||4||2|2|2|2|F|Black||15|No|Mother|28208|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016, PERL 2014-2016|Match Support|F|White||65|28205|Masters Degree|Divorced|Business|28255|40|5|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504089123|504091153|31|0|2|504383897|1|0|2|500920566|10|1|500014504||2|1|500014505, 500014681, 500016394|-1|500014505, 500016394|-1|0|4|||46|2|||1||702163000107564368|0
M587|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|678|Green|PERL 2014-2016|2014-11-13|2014-11-25|2016-10-03|Child: Changed school/site|Child: Changed school/site||22.3||2|2|2|2|F|Black||15|No|Mother|28208|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016, PERL 2014-2016|Match Support|F|Black||29|28262||Married|Customer Service|28217|1|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|504089123|504091153|31|0|2|503680769|31|0|2|500795303|10|1|500009132|2128207319|4|1|500014505, 500014681, 500016394|-1||-1|0|4|||11247|3|||1|500014681|702163000107564368|0
M588|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||2|2|1|1|M|Black||15|Yes|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||Self|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||25|28207|Bachelors Degree|Single|Finance|28269|0|0|Recruitment Event|Self|Big|General Site|mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|503624276|503626165|31|0|1|504786758|1|0|1|500922054|10|1|500014504||2|1|500014505, 500016394|-1|500016394|-1|0|10|||7458|9|||1||702163000107564368|0
M589|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|366|Green||2014-04-25|2014-04-29|2015-04-30|Volunteer: Time constraint|Volunteer: Time constraint||12||1|1|1|1|M|White||15|No|Mother|28211|7|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||63|28105|Bachelors Degree|Married|Self-Employed, Entrepreneur|28105|7|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503770826|503772799|1|0|1|503820142|1|0|1|500761166|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1||2811191761055817959|7044657180546140448
M590|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1189|Green||2013-11-20|2013-12-04|NaT||||39.1||1|1|1|1|M|Black||15|No|Mother|28213|9|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||31|28203||Single|Law|28202|3|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|503328958|503330792|31|0|1|503574852|1|0|1|500733114|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||7432163260389731024|514301162572611567
M591|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1436|Green||2012-05-07|2012-06-11|2016-05-17|Volunteer: Time constraint|Volunteer: Time constraint||47.2||3|3|1|1|F|Black||15|Yes|Mother|28216|7|One Parent: Female|$35,000 to $39,999|||Y|No||Self|General Community|Amachi|Enrollment|F|Black||34|28215|Some College|Single|Customer Service||0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|501253965|503287812|31|0|2|502985911|31|0|2|500613577|5|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1||9134125726462845918|0
M592|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|630|Green|PERL 2014-2016|2015-06-09|2015-06-16|NaT||||20.7||1|1|1|1|M|Black||15|No|GrandMother|28208|7|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|3|10|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|503944459|503946467|31|0|1|504260502|1|0|1|500829606|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||7462|13|||1|500014681|3935539763241716148|7044657180546140448
M593|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|360|Yellow||2014-11-07|2014-11-07|2015-11-02|Child/Family: Moved|Child/Family: Moved||11.8||1|1|2|2|M|Black||15|No|Mother|28217|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||63|28216|Some College|Single|Business|28217|1|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|504089059|504091089|31|0|1|504024774|31|0|1|500793445|10|1|500009132|2128207319|4|2||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M594|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|493|Green|mentor2.0, mentor2.0 2016|2015-10-16|2015-10-31|NaT||||16.2||1|1|1|1|F|Black||15|No|Mother|28207|9|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||38|28273|Bachelors Degree|Married|Business|28217|14|0|LPL Financial|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504416202|504418454|31|0|2|504394234|1|0|2|500848807|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||11247|3|||1|500014505, 500016394|702163000107564368|6780434725479563638
M595|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|221|Green|PERL 2014-2016|2016-01-11|2016-01-21|2016-08-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.3||1|1|1|1|M|Black||15|No|Mother|28269|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Multi-race (Black & White)||27|28115|Bachelors Degree|Single|Business|28115|4|4|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500017777|504268284|504270481|31|0|1|503172653|36|0|1|500871097|10|2|-2||4|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500014681|2798582775385400033|2378213070582218846
M596|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|518|Green|PERL 2014-2016|2015-02-10|2015-02-10|2016-07-12|Child: Changed school/site|Child: Changed school/site||17||1|1|3|3|M|Black||15|No|Mother|28217|8|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|M|Black||31|29710|Bachelors Degree|Married|Consultant|28217|3|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504207081|504209193|31|0|1|504060437|31|0|1|500812949|10|1|500009132|2128207319|4|1|500014681|-1||-1|0|4|||11247|3|||1|500014681|3935539763241716148|0
M597|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3480|Green|Amachi|2007-08-02|2007-08-27|NaT||||114.3||1|1|2|2|F|Black||15|Yes|Mother|28227|9|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||51|28216|Bachelors Degree|Divorced|Business: Clerical|28204|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500961274|500934638|31|0|2|500403000|31|0|2|500186952|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|4565518866290635873|0
M598|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|433|Green||2014-04-08|2014-04-30|2015-07-07|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||14.2||1|1|1|1|M|Black||15|No|Mother|28206|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Enrollment|M|Black||35|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28202|3|6|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503770380|503772356|31|0|1|503833456|31|0|1|500758739|5|1|500000295|2128173561|4|1||-1||-1|0|4|||7464|9|||1||7960300212314874874|0
M599|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1076|Green||2014-03-24|2014-03-27|NaT||||35.4||1|1|1|1|M|Black||15|No|Mother|28215|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Black||30|28202|Bachelors Degree|Single|Consultant|28281|2|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503758675|503760648|31|0|1|503792275|31|0|1|500756323|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||2129686509389594346|7044657180546140448
M600|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|493|Green|mentor2.0, mentor2.0 2016|2015-10-16|2015-10-31|NaT||||16.2||1|1|1|1|F|Black||15|No|Mother|28208|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0 2016|Match Support|F|Black||32|28269|Masters Degree|Single|Finance: Auditor|28217|1|0|LPL Financial|Workplace Partner|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504428649|504430904|31|0|2|504396801|31|0|2|500848796|10|1|500014504||2|1|500016394|-1|500014505, 500016394|-1|0|4|||11247|3|||1|500014505, 500016394|702163000107564368|0
M601|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|881|Green|PERL 2014-2016|2014-09-18|2014-10-08|NaT||||28.9||1|1|1|1|M|Black||15|No|Mother|28273|6|One Parent: Female|$20,000 to $24,999||||No||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28277|Bachelors Degree|Single|Business: Marketing|29067|0|3|Man Up Campaign|Media|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020910|503704573|503706538|31|0|1|503883049|1|0|1|500776636|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||17101|1|||1|500014681|3935539763241716148|2676951287175971833
M602|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2406|Green|Amachi|2010-07-26|2010-08-05|NaT||||79||1|1|2|2|M|Black||15|Yes|Mother|28215|6|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|Black||50|28078|||Service: Restaurant|28082|0|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|502183217|502183646|31|0|1|501733851|31|0|1|500462588|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294|4952249713946979108|0
M603|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|330|Green||2014-04-11|2014-04-30|2015-03-26|Volunteer: Time constraint|Volunteer: Time constraint||10.8||1|1|1|1|F|Black||14|Yes|Mother|28214|5|One Parent: Female|$35,000 to $39,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Some Other Race||34|28216|Masters Degree|Living w/ Significant Other|Finance: Banking|28216|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018850|503707241|503709207|31|0|2|503767700|41|0|2|500759405|5|2|-2||4|1|500000294|-2||-2|34|2|||7464|9|||1||2437132833506538679|1451515662136476632
M604|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|135|Green|PERL 2014-2016|2015-10-01|2015-10-21|2016-03-04|Child/Family: Moved|Child/Family: Moved||4.4||1|1|2|2|M|Black||14|No|Mother|28212|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|Amachi, PERL 2014-2016|Enrollment|M|White||30|28209|Bachelors Degree|Married|Real Estate: Realtor|28217|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|503863366|503865360|31|0|1|504322037|1|0|1|500843765|5|2|-2||4|1|500000294, 500014681|-2||-2|0|5|||46|2|||1|500014681|3292090474897428830|0
M605|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1174|Yellow||2012-05-11|2012-06-01|2015-08-19|Volunteer: Moved|Volunteer: Moved||38.6||1|1|1|1|F|Black||14|No|Mother|28269|4|One Parent: Female|$20,000 to $24,999||||No||Self|General Community||Match Support|F|White||27|28269|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502896719|502898127|31|0|2|502959645|1|0|2|500614239|10|2|-2||4|2||-2||-2|0|10|||46|2|||1||7679812394383646966|0
M606|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|774|Green|PERL 2014-2016|2015-01-13|2015-01-23|NaT||||25.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||37|28215|Masters Degree|Married|Finance: Banking|28262|15|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|503224764|503226552|31|0|1|504130394|31|0|1|500807724|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||46|2|||1|500014681|6724463016047116758|0
M607|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green|mentor2.0 2016|2016-10-31|2016-11-18|NaT||||3.6||1|1|2|2|M|Hispanic||14|No|Mother|28217|9|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|Hispanic||42|28209|Masters Degree|Married|Finance: Banking|28255|12|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831713|504834215|3|0|1|504380428|3|0|1|500921929|10|1|500014504||2|1|500014505, 500016394|-1|500015184|-1|0|4|||17159|12|||1|500016394|702163000107564368|0
M608|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|987|Green||2014-06-10|2014-06-24|NaT||||32.4||2|2|1|1|F|Black||14|No|Mother|28215|6|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||27|28209|Bachelors Degree|Single|Finance|28202|2|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503318449|503320281|31|0|2|503775488|1|0|2|500766059|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||675142027733303647|6178126991714892144
M609|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2870|Green||2009-04-17|2009-04-28|NaT||||94.3||1|1|1|1|M|White||14|No|Mother|28262|6|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||46|28078|Masters Degree|Single|Retail: Mgt|28207|1|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|501599416|501599736|1|0|1|500188567|1|0|1|500357914|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||4621676786129919860|5529223012138448528
M610|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1713|Green||2012-06-22|2012-06-28|NaT||||56.3||1|1|1|1|M|Black||14|No|Mother|28226|7|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||46|28134|Bachelors Degree|Married|Finance|28105|1|6|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020752|502183053|502183482|31|0|1|503073638|31|0|1|500621039|10|2|-2||2|1||-2|500014681|-2|0|10|||4748|14|633|1|1||4112464363801619560|0
M611|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|136|Green||2016-05-11|2016-06-20|2016-11-03|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.5||1|1|1|1|F|Black||14|No|GrandMother|28105|9|Grandparents|$45,000 to $49,999||||Yes|BBBS National Site|Web Link|General Community||RTBM|F|Black||39|28105|Bachelors Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504631841|504634252|31|0|2|504167347|31|0|2|500892753|7|2|-2||4|1||-2||-2|34|2|||7464|9|||1||2129686509389594346|5605796235524810842
M612|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|740|Green||2015-02-24|2015-02-26|NaT||||24.3||1|1|1|1|M|Black||14|No|Mother|28278|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|Black||29|28209|Bachelors Degree|Single|Finance|20877|0|8|TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504160892|504162947|31|0|1|504171934|31|0|1|500815454|10|2|-2||2|1||-2||-2|0|4|||130|1|||1||8567789404096574827|2876415545463317777
M613|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1694|Green||2012-07-05|2012-07-17|NaT||||55.7||2|2|1|1|F|Black||14|No|Mother|28214|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||49|28215|Bachelors Degree|Married|Business: Mgt, Admin|28277|13|0|Local Print|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502566369|502566823|31|0|2|503065299|1|0|2|500622859|10|2|-2||2|1||-2||-2|0|10|||7439|1|||1||7089569121628268952|0
M614|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||1|1|1|1|M|Hispanic||14|No|Mother|28214|9|Two Parent|$30,000 to $34,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||28|28208|PHD|Single|Tech: Management|28208|5|2|Current/Previous Big|Other Big|Big|General Site|mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504870363|504872882|3|0|1|504719047|1|0|1|500921854|10|1|500014504||2|1|500014505, 500016394|-1|500016394|-1|0|4|||17159|12|||1||702163000107564368|0
M615|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|249|Green||2015-11-04|2015-11-05|2016-07-11|Child: Changed school/site|Child: Changed school/site||8.2||1|1|2|2|M|Black||14|No|Mother|28206|8|One Parent: Male|Unknown||||Yes||Relative|General Site||Match Support|M|Black||63|28216|Some College|Single|Business|28217|1|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504506841|504509136|31|0|1|504024774|31|0|1|500856384|10|1|500009132|2128207319|4|1||-1||-1|0|3|||11247|3|||1||3935539763241716148|0
M616|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1086|Green||2014-02-03|2014-02-05|2017-01-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.7||1|1|1|1|M|Black||14|No|Mother|28262|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Multi-race (Hispanic & White)||33|28226|Some College|Single|Tech: Management|28277|1|7|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503219503|503221284|31|0|1|503589945|35|0|1|500746532|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||3677730851176818072|7044657180546140448
M617|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|771|Green||2015-01-08|2015-01-26|NaT||||25.3||2|2|1|1|F|Black||14|No|Mother|28206|8|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||30|28205|Bachelors Degree|Single|Human Services|28203|1|2|TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503816186|501097065|31|0|2|504090792|1|0|2|500807024|10|2|-2||2|1||-2||-2|0|10|||130|1|||1||932861092942387634|7044657180546140448
M618|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1705|Green||2012-06-19|2012-06-29|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||56||1|1|1|1|F|Black||14|No|Mother|28217|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||31|28211|Bachelors Degree|Single|Real Estate: Realtor|19137|2|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502920377|502921794|31|0|2|502942994|1|0|2|500620441|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||0|0
M619|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|577|Green||2013-10-29|2013-11-18|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19||1|1|1|1|F|Black||14|No|Mother|28205|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||28|28202|||Business|28202|0|0|Duke Energy|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503566749|503568624|31|0|2|503605700|1|0|2|500724784|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M620|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|161|Yellow||2015-07-30|2015-07-30|2016-01-07|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||5.3||1|1|1|1|M|Black||14|No|Mother|28217|6|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||31|28209|Bachelors Degree|Single|Human Services|28203|1|8|Current/Previous Big|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500018851|503063769|503065429|31|0|1|504299841|1|0|1|500834948|10|2|-2||4|2||-2||-2|34|2|||17159|12|||1||7960300212314874874|2141487034287122220
M621|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1325|Green||2013-07-08|2013-07-21|NaT||||43.5||1|1|1|1|M|Black||14|No|Mother|28212|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||28|28273|Bachelors Degree||Business|28217|2|0|Elevation Church|Faith Organization|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503511553|503513424|31|0|1|503504991|1|0|1|500702866|10|2|-2||2|1||-2||-2|0|10|||16414|7|||1||2811191761055817959|0
M622|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3456|Green||2007-09-12|2007-09-20|NaT||||113.5|Y|1|1|1|1|M|Black||14|No|Mother|28210|5|One Parent: Female|$20,000 to $24,999||||No||Self|General Community||Match Support|M|White||54|28207||Married|Business: Sales||0|0|Recruitment Event|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500868942|500869211|31|0|1|500947018|1|0|1|500195082|10|2|-2||2|1||-2||-2|0|10|||7458|9|||1||5473689050106799364|0
M623|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1154|Yellow||2013-03-14|2013-03-27|2016-05-24|Volunteer: Moved|Volunteer: Moved||37.9||1|1|1|1|M|Black||14|No|Mother|28262|5|One Parent: Female|$45,000 to $49,999||||No||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Mgt, Admin|28217|3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503110829|503112489|31|0|1|503130981|1|0|1|500687926|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||0|7674215580094440446
M624|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|225|Red|PERL 2014-2016|2015-04-11|2015-04-21|2015-12-02|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.4||1|1|2|2|M|Black||14|No|Mother|28213|7|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|PERL 2014-2016|RTBM|M|White||32|28202|Masters Degree|Single|Finance: Accountant|28202|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500013781|503917561|503962680|31|0|1|504206321|1|0|1|500822824|7|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|500014681|3677730851176818072|6084148439133243542
M625|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|243|Red||2014-10-20|2014-10-31|2015-07-01|Volunteer: Moved|Volunteer: Moved||8||3|3|1|1|F|Black||14|No|Mother|28269|3|Two Parent|Unknown||||Yes||Relative|General Community||Match Support|F|Black||29|28262||Single|Military|28308|5|0|Local TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502229042|502172965|31|0|2|503849760|31|0|2|500785297|10|2|-2||4|3||-2||-2|0|3|||7438|1|||1||4208486535559819469|0
M626|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|222|Green|PERL 2014-2016|2015-12-02|2015-12-02|2016-07-11|Child: Changed school/site|Child: Changed school/site||7.3||1|1|1|1|M|Black||14|No|Mother|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Site|PERL 2014-2016|Match Support|M|Black||38|28277|Associate Degree|Married|Business|28217|0|6|LPL Financial|Workplace Partner|Big|General Site|PERL 2014-2016|RTBM|0|1|1|0|277|60|598|500000170|500015820|504526211|504528543|31|0|1|504528256|31|0|1|500864681|10|1|500009132|2128207319|4|1|500014681|-1|500014681|-1|0|3|||11247|3|||1|500014681|3935539763241716148|0
M627|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1104|Green|Cabarrus County|2014-02-04|2014-02-27|NaT||||36.3||1|1|1|1|F|White||14|No|Father|28081|9|One Parent: Male|$15,000 to $19,999||||Yes||Self|General Community|Cabarrus County|Match Support|F|White||28|28209|Bachelors Degree|Single|Finance|28217|3|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500013781|503634718|503636659|1|0|2|503595858|1|0|2|500746721|10|2|-2||2|1|500016374|-2|500016374|-2|0|10|||7458|9|||1|500016374|0|1786514887916898235
M628|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|858|Green|PERL 2014-2016, Cabarrus County|2014-10-27|2014-10-31|NaT||||28.2||1|1|1|1|M|White||14|No|Father|28081|8|One Parent: Male|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||28|28277|Bachelors Degree||Finance|28255|0|4|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500013781|503961917|503636659|1|0|1|504052039|1|0|1|500788399|10|2|-2||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|5|||17159|12|||1|500014681, 500016374|5273065343662533495|1786514887916898235
M629|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|106|Green||2016-10-26|2016-11-21|NaT||||3.5||1|1|1|1|M|Multi-race (Hispanic & White)||14|No|Father|28208|9|Two Parent|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||29|28203|Bachelors Degree|Single|Business: Mgt, Admin||7|0|BBBS National Site|Web Link|Big|General Site|mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831449|504833951|35|0|1|504719321|1|0|1|500920204|10|1|500014504||2|1|500014505, 500016394|-1|500016394|-1|0|4|||46|2|||1||702163000107564368|0
M630|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|49|Green||2016-10-31|2017-01-17|NaT||||1.6||1|1|1|1|M|Hispanic||14|No|Father|28202|9|Two Parent|$10,000 to $14,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||24|28202|Bachelors Degree|Single|Business: Marketing||1|0|Community Engagement|Special Event|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504910946|504913466|3|0|1|504687842|1|0|1|500921850|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||18809|8|||1||702163000107564368|0
M631|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2302|Green|Amachi, Cabarrus County|2010-11-11|2010-11-17|NaT||||75.6||1|1|1|1|F|White||14|Yes|Mother|28025|7|Two Parent|Unknown|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||63|28027|High School Graduate|Married|Self-Employed, Entrepreneur|28027|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|501938282|501938680|1|0|2|502356100|1|0|2|500493871|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|500000294, 500016374|7450734758077775903|0
M632|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|580|Green||2013-10-29|2013-11-15|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19.1||4|4|1|1|M|Black||14||Mother|28269|6|One Parent: Female|Unknown||||No||School|General Site||Match Support|M|White||29|28246||Married|Tech: Engineer|28202|3|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|501152789|501153063|31|0|1|503604690|1|0|1|500724447|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M633|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2024|Green|Amachi|2011-08-22|2011-08-22|NaT||||66.5||1|1|1|1|M|Multi-race (Black & Hispanic)||14|No|Mother|28208|7|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||28|28262|High School Graduate|Single|Laborer||0|8|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502245129|502245570|38|0|1|502670839|31|0|1|500551050|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1|500000294|1653226628427425023|0
M634|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|326|Green|PERL 2014-2016|2015-11-03|2015-11-19|2016-10-10|Volunteer: Moved|Volunteer: Moved||10.7||1|1|1|1|M|White||14|No|Mother|28209|7|One Parent: Female|$20,000 to $24,999||||No||Self|General Community|PERL 2014-2016|Enrollment|M|White||27|28278|Masters Degree|Married|Business: Engineer|28278|2|8|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch Training Final Assessment|Match Support|0|1|1|0|277|60|598|500000170|500018851|504298668|504300882|1|0|1|504372921|1|0|1|500855505|5|2|-2||4|1|500014681|-2|500011316|-2|0|10|||17159|12|||1|500014681|4440360203097874486|2656293275676608966
M635|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-27|2016-11-02|NaT||||4.1||1|1|1|1|F|Hispanic||14|No|Mother|28217|9|One Parent: Female|Less than $10,000||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||31|28270|Bachelors Degree|Single|Medical|28277|4|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831525|504834027|3|0|2|504765443|1|0|2|500920670|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M636|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte||N|S|Active|Match Support|125|Green||2016-10-26|2016-11-02|NaT||||4.1||2|2|2|2|F|Black||14|No|Mother|28208|9|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Site|Amachi, mentor2.0, mentor2.0 2016|Match Support|F|Black||45|28217|Bachelors Degree|Divorced|Education: Teacher|28226|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|0|1|277|60|598||0|503492214|503494082|31|0|2|504272278|31|0|2|500920167|10|1|500014504||2|1|500000294, 500014505, 500016394|-1|500015184|-1|0|10|||7462|13|||1||702163000107564368|7044657180546140448
M637|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1130|Yellow||2012-08-30|2012-09-11|2015-10-16|Child/Family: Moved|Child/Family: Moved||37.1||1|1|1|1|F|Black||14|No|Mother|28212|6|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||32|28204|Bachelors Degree|Single|Business: Marketing|29730|0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503021417|501428579|31|0|2|503115600|1|0|2|500631553|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||4048394821927342477|0
M638|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|838|Green||2014-03-27|2014-04-16|2016-08-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||27.5||2|2|1|1|M|Black||14|No|Mother|28215|4|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|Black||32|28209|Masters Degree||Finance|28217|0|9|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|501662021|501090456|31|0|1|503759352|31|0|1|500757152|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1||2417657944362725638|4753237757252407321
M639|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|865|Green|PERL 2014-2016|2014-10-14|2014-10-24|NaT||||28.4||4|4|1|1|M|Black||14||Mother|28206|6|One Parent: Female|Unknown||||No||School|General Community|PERL 2014-2016|Match Support|M|White||29|28205|Bachelors Degree|Single|Finance: Banking|28262|4|0|Man Up Campaign|Web Link|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020910|501091420|501091694|31|0|1|503946168|1|0|1|500783556|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17100|2|||1|500014681|0|0
M640|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|296|Green||2014-11-17|2014-11-25|2015-09-17|Volunteer: Moved|Volunteer: Moved||9.7||2|2|1|1|F|Black||14|No|Mother|28206|7|One Parent: Female|Unknown|||Y|No||Relative|General Community||Enrollment|F|White||27|28278|Bachelors Degree|Single|Education: Teacher|28056|1|9|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|504081573|501091694|31|0|2|503880925|1|0|2|500796131|5|2|-2||4|1||-2||-2|0|3|||17159|12|||1||9134125726462845918|0
M641|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|215|Green||2016-01-13|2016-01-31|2016-09-02|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||7.1||2|2|1|1|F|Black||14|No|Mother|28206|7|One Parent: Female|Unknown|||Y|No||Relative|General Community||Enrollment|F|White||26|28211||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500017777|504081573|501091694|31|0|2|504317495|1|0|2|500871696|5|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|3|||17159|12|||1||9134125726462845918|0
M642|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2389|Green||2010-08-11|2010-08-22|NaT||||78.5||1|1|2|2|M|Black||14|No|Mother|28216|5|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502000252|502000651|31|0|1|502127058|1|0|1|500465318|10|2|-2||2|1||-2||-2|0|10|||130|1|||1||7857548027029642592|0
M643|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1700|Green||2012-06-14|2012-07-11|NaT||||55.9||1|1|1|1|F|Black||14|No|Mother|28208|4|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||30|28203|Bachelors Degree|Single|Business: Marketing|28117|0|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502902247|502903657|31|0|2|502801082|1|0|2|500619356|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||7857548027029642592|0
M644|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|775|Yellow||2013-12-03|2013-12-19|2016-02-02|Volunteer: Time constraint|Volunteer: Time constraint||25.5||1|1|1|1|M|Black||14|No|GrandMother|28206|7|One Parent: Female|Unknown|||Y|Yes||Self|General Site||Enrollment|M|Black||45|28273||Separated|Business|28244|2|6|Recruitment Event|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503515724|503517595|31|0|1|503689721|31|0|1|500736042|5|1|500000295|2128173561|4|2||-1||-1|0|10|||7458|9|||1||7960300212314874874|0
M645|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|728|Green||2013-11-13|2013-11-21|2015-11-19|Volunteer: Time constraint|Volunteer: Time constraint||23.9||2|2|1|1|M|Black||14|No|Mother|28206|5|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||32|28210|Some College||Business||0|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|502008563|502008962|31|0|1|503400112|1|0|1|500730792|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||0|8460600033983851488
M646|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|254|Green||2015-10-16|2015-10-31|2016-07-11|Child: Changed school/site|Child: Changed school/site||8.3||1|1|1|1|F|Black||14|No|Mother|28202|8|Two Parent|Less than $10,000|||Y|Yes||Relative|General Site||Match Support|F|Black||33|28054||Single|Consultant|28217|1|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504416129|504418381|31|0|2|504399706|31|0|2|500848800|10|1|500009132|2128207319|4|1||-1||-1|0|3|||11247|3|||1||3935539763241716148|0
M647|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|737|Green||2012-12-03|2013-01-26|2015-02-02|Volunteer: Time constraint|Volunteer: Time constraint||24.2||2|2|1|1|F|Black||14|No|Mother|28214|4|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||34|28262|Bachelors Degree|Single|Insurance||6|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|501147999|501148273|31|0|2|503112265|31|0|2|500665633|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1||6627885846854295604|3402014428779854546
M648|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-26|2016-11-02|NaT||||4.1||1|1|1|1|M|White||14|Yes|Mother|28208|9|One Parent: Female|Less than $10,000||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||30|28209|Bachelors Degree|Married|Finance|28217|1|6|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504888396|504890916|1|0|1|504767070|1|0|1|500920228|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M649|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1803|Green||2012-03-22|2012-03-30|NaT||||59.2||1|1|1|1|M|Black||14|No|Mother|28217|5|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||36|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502700503|502701348|31|0|1|502931327|1|0|1|500605634|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||0|0
M650|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|241|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-02|2016-05-31|2017-01-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.9||1|1|2|2|M|White||14|No|Mother|28214|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500013781|504231264|504233379|1|0|1|504230177|1|0|1|500891315|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|3|||7462|13|||1|500007920, 500011315, 500011316|9076057728106637014|0
M651|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|350|Green||2014-05-13|2014-05-29|2015-05-14|Volunteer: Time constraint|Volunteer: Time constraint||11.5||1|1|1|1|F|Black||14|No|Mother|28262|6|One Parent: Female|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community||Enrollment|F|White||28|28202|Masters Degree|Single|Finance: Banking|28205|0|1|Other|Service Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503813952|503969639|31|0|2|503829786|1|0|2|500763221|5|2|-2||4|1||-2||-2|34|2|||7452|6|||1||932861092942387634|6619197389800008587
M652|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|96|Yellow||2015-10-16|2015-10-31|2016-02-04|Child/Family: Moved|Child/Family: Moved||3.2||1|1|2|3|M|Black||14|No|Mother|28208|8|Two Parent|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|Black||30|28217|Bachelors Degree|Single|Business|28217|0|9|LPL Financial|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|504416115|504456768|31|0|1|504397175|31|0|2|500848794|10|1|500009132|2128207319|4|2||-1||-2|0|4|||11247|3|||1||3935539763241716148|0
M653|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||1|1|2|2|M|Hispanic||14|No|Mother|28217|9|Two Parent|$20,000 to $24,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||34|28202||Married|Consultant||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504842873|504845375|3|0|1|503969533|1|0|1|500922037|10|1|500014504||2|1|500014505, 500016394|-1|500014506, 500016394|-1|0|4|||7462|13|||1||702163000107564368|1321057499120459151
M654|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1553|Green||2012-11-13|2012-11-28|2017-02-28|Volunteer: Time constraint|Volunteer: Time constraint||51||2|2|1|1|F|Black||14|No|GrandMother|28206|4|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|F|Black||48|28213|Bachelors Degree|Single|Finance: Accountant||8|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501273088|501273365|31|0|2|503079327|31|0|2|500659156|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1||392688197545050058|7044657180546140448
M655|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|867|Green|PERL 2014-2016, Cabarrus County|2014-08-18|2014-10-22|NaT||||28.5||1|1|1|1|F|White||14|No|Father|28025|9|One Parent: Male|$40,000 to $44,999|||Y|No|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||31|28025|Bachelors Degree|Married|Business: Mgt, Admin|28027|4|7|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500022817|503952645|503954653|1|0|2|503942996|31|0|2|500772607|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|34|2|||7464|9|||1|500014681, 500016374|0|6967646101447772925
M656|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|652|Red|PERL 2014-2016|2015-01-07|2015-01-27|2016-11-09|Child: Lost interest|Child: Lost interest||21.4||1|1|4|5|F|White||14|No|Mother|28025|8|One Parent: Female|$35,000 to $39,999||||No||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|0|1|1|0|277|60|598|500000170|500020753|503923436|503925443|1|0|2|501306527|1|0|2|500806777|10|2|-2||4|3|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||7464|9|||1|500014681|6750834084344455219|0
M657|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|296|Green||2015-09-23|2015-10-05|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|1|1|F|Black||14|No|Mother|28208|7|One Parent: Female|$10,000 to $14,999||||Yes||Self|General Site||Match Support|F|White||50|28269||Married|Finance|28208|6|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333795|504336017|31|0|2|504348509|1|0|2|500841761|10|1|500009132|2128207318|4|1||-1||-1|0|10|||12831|3|||1||2611337051335117774|5181319291190669508
M658|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|231|Red||2014-12-18|2015-01-12|2015-08-31|Child/Family: Moved|Child/Family: Moved||7.6||1|1|1|1|F|Multi-race (Black & White)||14|No|Mother|28217|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||49|28210|Masters Degree|Divorced|Education|28211|6|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503535105|503536977|36|0|2|504127300|1|0|2|500805104|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||9134125726462845918|0
M659|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-31|2016-11-02|NaT||||4.1||1|1|2|2|F|Multi-race (Black & White)||14|No|GrandMother|28217|9|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||24|28202||Single|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500022907|504859921|504862440|36|0|2|504353872|1|0|2|500921831|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500015184|-1|0|4|||17159|12|||1||702163000107564368|0
M660|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|255|Green|PERL 2014-2016|2015-10-16|2015-10-30|2016-07-11|Child: Changed school/site|Child: Changed school/site||8.4||1|1|1|1|M|Black||14|No|Mother|28208|8|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|F|White||28|28209|Bachelors Degree|Single|Business: Mgt, Admin|28217|2|0|LPL Financial|Workplace Partner|Big|General Site|PERL 2014-2016|RTBM|0|1|1|0|277|60|598|500000170|500015820|504416012|504418264|31|0|1|504397015|1|0|2|500848797|10|1|500009132|2128207319|4|1|500014681|-1|500014681|-1|0|4|||11247|3|||1|500014681|3935539763241716148|0
M661|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|382|Red||2014-08-20|2014-08-30|2015-09-16|Child/Family: Moved|Child/Family: Moved||12.6||1|1|1|1|M|Black||14|No|Mother|28269|6|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|M|Black||62|28210|Bachelors Degree|Divorced|Business|28202|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503838769|503840748|31|0|1|503948333|31|0|1|500772925|10|2|-2||4|3||-2||-2|0|10|||7671|13|||1||7184048822538031021|6837005360290527271
M662|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-27|2016-11-04|NaT||||4||1|1|1|1|M|Black||14|No|Mother|28208|9|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||28|28206|Bachelors Degree|Single|Finance|28203|4|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504861242|504863761|31|0|1|504786813|1|0|1|500920585|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M663|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3401|Green|Amachi|2007-10-30|2007-11-07|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||111.7||1|1|1|1|M|Black||14|Yes|Mother|28213||One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||66|28075||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|501069450|501048131|31|0|1|500887364|31|0|1|500212043|10|2|-2||4|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294|8461485523552765256|0
M664|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|254|Green||2015-10-16|2015-10-31|2016-07-11|Child: Changed school/site|Child: Changed school/site||8.3||1|1|1|1|M|Black||14|No|Mother|28217|8|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Native Hawaiian or Other Pacific Islander||30|28204|Bachelors Degree|Single|Consultant|28217|0|6|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504416100|504418352|31|0|1|504455617|5|0|1|500848795|10|1|500009132|2128207319|4|1||-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M665|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|495|Red||2015-05-20|2015-05-20|2016-09-26|Child/Family: Moved|Child/Family: Moved||16.3||1|1|1|1|M|Black||14|No|Mother|28269|6|One Parent: Female|$35,000 to $39,999|Yes: Active|No||No||Self|General Community||Match Support|M|White||53|28203|Masters Degree|Married|Business: Sales|17601|0|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503874068|503876064|31|0|1|504196201|1|0|1|500827631|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||1320477920662455183|3501831218874457455
M666|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1260|Green||2013-09-11|2013-09-24|NaT||||41.4||1|1|2|2|M|Multi-race (Black & Hispanic)||14|No|Mother|28273|5|One Parent: Female|$50,000 to $59,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|1|0|0|1|277|60|598|500000170|500008321|503361148|503362993|38|0|1|502459922|1|0|1|500710308|10|2|-2||2|1||-2|500004640|-2|34|2|||7464|9|||1||6202343250032725030|1001458554309997291
M667|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|705|Red|PERL 2014-2016|2015-03-26|2015-03-26|2017-02-28|Volunteer: Moved|Volunteer: Moved||23.2||1|1|1|1|M|Black||14|No|Mother|28262|7|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||32|28262|Bachelors Degree|Single|Customer Service|28262|2|6|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500008321|504045474|504047495|31|0|1|504228594|31|0|1|500820783|10|2|-2||4|3|500014681|-2|500014681|-2|0|10|||46|2|||1|500014681|5441374193599827162|3402014428779854546
M668|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|619|Green|PERL 2014-2016|2014-11-04|2014-11-10|2016-07-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||20.3||1|1|3|3|F|Black||14|No|Mother|28205|7|One Parent: Female|Unknown||||No||School|General Site|PERL 2014-2016|Match Support|F|Black||36|28269||Single|Business|28202|7|5|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|504087114|504089144|31|0|2|503605618|31|0|2|500791543|10|1|500000295|2128173561|4|1|500014681|-1|500014681|-1|0|4|||16705|3|||1|500014681|7960300212314874874|0
M669|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1680|Green||2012-07-05|2012-07-31|NaT||||55.2||1|1|1|1|F|Black||14|No|Mother|28031|4|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Mgt, Admin|28078|1|11|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502863776|502865175|31|0|2|503029273|1|0|2|500622877|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||927920773840777760|1286881276054717070
M670|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3042|Green|Amachi|2008-10-28|2008-11-07|NaT||||99.9||2|2|1|1|F|Black||14|Yes|Mother|28217|9|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||48|28205|Bachelors Degree|Living w/ Significant Other|Human Services: Non-Profit|28205|3|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501014187|500948399|31|0|2|501404007|1|0|2|500306699|10|2|500003586||2|1|500000294|-2||-2|0|10|||7671|13|||1|500000294|702163000107564368|0
M671|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1890|Green|Project Big|2011-04-25|2011-06-27|2016-08-29|Volunteer: Time constraint|Volunteer: Time constraint||62.1||1|1|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community|Project Big|Enrollment|F|Black||33|28215|Bachelors Degree|Single|Human Services: Social Worker|28217|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|1|0|1|0|277|60|598|500000170|500017777|502303088|502303520|31|0|2|502445797|31|0|2|500533193|5|2|-2||4|1|500004640|-2|500000294, 500004640|-2|6854|8|||7464|9|||1|500004640|932861092942387634|0
M672|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2132|Red|Amachi, Project Big, Project Big AND Amachi|2010-11-16|2010-12-30|2016-10-31|Child: Lost interest|Child: Lost interest||70||1|1|1|1|M|Black||14|Yes|Mother|28213|4|One Parent: Female|Unknown||||Yes||School|General Community|Project Big AND Amachi|Match Support|M|White||27|28262||Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|1|0|1|0|277|60|598|500000170|500008321|502335675|502336110|31|0|1|502305990|1|0|1|500495220|10|2|500004772||4|3|500004901|-2|500000294, 500004640|-2|0|4|||7496|10|||1|500000294, 500004640, 500004901|6065435025527210335|0
M673|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|439|Green||2014-09-29|2014-10-15|2015-12-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|Black||32|28202|Bachelors Degree|Single|Consultant|28202|0|9|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503849038|503851023|31|0|1|503930671|31|0|1|500778856|10|2|-2||4|1||-2||-2|0|10|||17101|1|||1||7883015200677941272|2793519126277633342
M674|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1449|Green||2013-03-13|2013-03-19|NaT||||47.6||1|1|1|1|M|Black||14|No|Mother|28214|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||32|29708|Bachelors Degree|Married|Finance||0|9|Local TV|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502858216|502859613|31|0|1|503376842|1|0|1|500687641|10|2|-2||2|1||-2||-2|0|10|||7438|1|||1||9076057728106637014|7044657180546140448
M675|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|126|Green||2016-10-25|2016-11-01|NaT||||4.1||1|1|1|1|M|Black||14|No|Mother|28208|9|One Parent: Female|$30,000 to $34,999||||No||School|General Site|mentor2.0|Match Support|M|White||27|28226|Bachelors Degree|Single|Insurance||0|6|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831574|504834076|31|0|1|504756883|1|0|1|500919677|10|1|500014504||2|1|500014505|-1|500014505, 500016394|-1|0|4|||17159|12|||1||702163000107564368|0
M676|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-27|2016-11-02|NaT||||4.1||1|1|1|1|F|Hispanic||14|No|Father|28217|9|One Parent: Male|Unknown|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||26|28078|Masters Degree|Married|Education|27360|2|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831771|504834273|3|0|2|504784525|1|0|2|500920641|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M677|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|256|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment, PERL 2014-2016|2015-12-07|2015-12-17|2016-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.4||1|1|1|1|M|Black||14|No|Mother|28269|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||RTBM|M|Black||40|28269|Bachelors Degree|Married|Tech: Support, Writing|28269|4|0|Local Radio|Media|Big|General Community|Amachi, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500017777|504245120|504247236|31|0|1|504396885|31|0|1|500865817|7|2|-2||4|1||-2|500000294, 500007920, 500011315, 500011316, 500014681|-2|0|4|||7437|1|||1|500007920, 500011315, 500011316, 500014681|9134125726462845918|1546374315672654438
M678|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3214|Green||2008-04-24|2008-05-19|NaT||||105.6||1|1|1|1|F|White||14|No|Father|28207|1|One Parent: Male|Unknown||||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Finance: Banking|28255|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501213488|501213764|1|0|2|501225276|1|0|2|500262655|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||0|0
M679|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|595|Green||2013-10-11|2013-10-30|2015-06-17|Child/Family: Time constraints|Child/Family: Time constraints||19.5||1|1|1|1|F|Black||14|Yes|Mother|28262||One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Finance|28202|0|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503587461|503587387|31|0|2|503541106|1|0|2|500718377|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||3677730851176818072|5766455966581408090
M680|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1035|Green||2014-04-07|2014-05-07|NaT||||34||3|3|1|1|F|Black||14|No|Mother|28209||One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|White||32|28277|Bachelors Degree|Single|Real Estate: Realtor|28202|1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500021785|502254067|502254499|31|0|2|503590595|1|0|2|500758482|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||0|0
M681|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|127|Green|mentor2.0, mentor2.0 2016|2016-10-31|2016-10-31|NaT||||4.2||3|4|2|2|F|Black||14|No|Mother|28217|7|Two Parent|$15,000 to $19,999|||Y|No||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||31|28203|High School Graduate|Single|Business: Sales|28281|3|3|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|501092822|501093096|31|0|2|503854063|1|0|2|500921966|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||46|2|||1|500014505, 500016394|8567789404096574827|358434295995756137
M682|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|959|Green||2014-06-27|2014-07-22|NaT||||31.5||3|4|2|2|F|Black||14|No|Mother|28217|7|Two Parent|$15,000 to $19,999|||Y|No||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||31|28203|High School Graduate|Single|Business: Sales|28281|3|3|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|1|0|0|1|277|60|598|500000170|500013781|501092822|501093096|31|0|2|503854063|1|0|2|500768017|10|2|-2||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||46|2|||1||8567789404096574827|358434295995756137
M683|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|802|Green||2013-12-11|2014-02-21|2016-05-03|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||26.3||1|1|1|1|F|Black||14|No|Mother|28212|6|One Parent: Female|$20,000 to $24,999|||Y|No||School|General Community||Match Support|F|Black||28|28216|Masters Degree|Single|Consultant|28205|0|0|Recruitment Event|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500021785|503441472|501290021|31|0|2|503551607|31|0|2|500738115|10|2|-2||4|1||-2||-2|0|4|||7458|9|||1||2811191761055817959|7044657180546140448
M684|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|131|Green||2016-09-22|2016-10-27|NaT||||4.3||1|1|1|1|F|Black||14|Yes|Mother|28208|8|Two Parent|$15,000 to $19,999||||Yes||School|General Site||Match Support|F|White||24|28006|Bachelors Degree|Single|Business|28208|1|3|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504855873|504858375|31|0|2|504783357|1|0|2|500909621|10|1|500009132|2128212899|2|1||-1||-1|0|4|||7464|9|||1||8568001799025358453|0
M685|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|612|Green|Amachi, PERL 2014-2016|2014-11-07|2014-11-07|2016-07-11|Child: Changed school/site|Child: Changed school/site||20.1||1|1|2|2|M|Black||14|Yes|Mother|28217|8|One Parent: Female|Unknown||||Yes||School|General Site|Amachi, PERL 2014-2016|Match Support|M|White||31|29707|Bachelors Degree|Married|Customer Service||0|0|LPL Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500015820|502178448|502178877|31|0|1|504024654|1|0|1|500793402|10|1|500009132|2128207319|4|1|500000294, 500014681|-1|500014681|-1|0|4|||11247|3|||1|500000294, 500014681|3935539763241716148|0
M686|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|68|Red||2016-12-01|2016-12-22|2017-02-28|Child/Family: Moved|Child/Family: Moved||2.2||1|1|1|1|M|Black||14|No|Mother|28215|9|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Black||32|28213|Masters Degree|Married|Finance: Auditor|28202|0|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500020753|504851045|504853547|31|0|1|504774982|31|0|1|500932246|10|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316|-2|0|5|||46|2|||1||0|2141487034287122220
M687|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|177|Green||2015-09-17|2015-09-22|2016-03-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||5.8||2|2|1|1|F|Black||14|No|GrandMother|28206|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Native Hawaiian or Other Pacific Islander||39|28211|Masters Degree|Married|Business|28204|8|0|Igniting Breakfast|Special Event|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500017732|502619926|502620542|31|0|2|504288677|5|0|2|500840540|10|2|-2||4|1||-2||-2|0|10|||17266|8|||1||1653226628427425023|0
M688|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1365|Green|Project Big|2011-07-29|2011-08-09|2015-05-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||44.8||2|2|1|1|F|Black||14|No|GrandMother|28206|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||38|28205|Bachelors Degree|Single|Law: Lawyer|28202|2|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502619926|502620542|31|0|2|502642260|1|0|2|500548116|10|2|500004641||4|1||-2||-2|0|10|||7464|9|||1|500004640|1653226628427425023|0
M689|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1642|Green||2010-09-20|2010-10-01|2015-03-31|Child/Family: Moved|Child/Family: Moved||53.9||1|1|1|1|F|Black||14|No|Mother|28208|3|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||37|28277|PHD|Single|Medical: Healthcare Worker||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|502273093|502273525|31|0|2|502252422|31|0|2|500471568|10|2|-2||4|1||-2|500000294|-2|0|4|||7496|10|||1||0|3402014428779854546
M690|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||1|1|1|1|F|Black||14|No|Mother|28216|9|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|Black||32|28210|Bachelors Degree|Single|Finance|28202|0|0|Self|Self|Big|General Site|mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504842845|504845347|31|0|2|504794021|31|0|2|500921980|10|1|500014504||2|1|500014505, 500016394|-1|500016394|-1|0|4|||7464|9|||1||702163000107564368|3402014428779854546
M691|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|228|Green|PERL 2014-2016|2016-06-30|2016-07-22|NaT||||7.5||1|1|2|2|M|Black||14|No|GrandMother|28208|7|One Parent: Female|$20,000 to $24,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||29|28209|Masters Degree|Single|Business|29707|0|8|Community Engagement|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|503711736|503713702|31|0|1|501121735|1|0|1|500898534|10|2|-2||2|1||-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||18809|8|||1|500014681|7581500809034284566|3402014428779854546
M692|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||1|1|3|3|F|Asian||14|No|Father|28208|9|Two Parent|Unknown||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||40|28078|Bachelors Degree|Single|Human Services: Social Worker|28277|0|9|Relative|Relative|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831791|504834293|4|0|2|503529603|1|0|2|500922070|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500015184|-1|0|4|||17161|11|||1||702163000107564368|0
M693|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1570|Yellow|Amachi|2010-09-27|2010-09-28|2015-01-15|Volunteer: Time constraint|Volunteer: Time constraint||51.6||2|2|1|1|M|Multi-race (Black & White)||14|Yes|GrandMother|28215|7|Grandparents|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||58|28226|Masters Degree|Married|Tech: Sales, Mktg|28202|6|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|502183420|502183840|36|0|1|502264770|1|0|1|500473793|10|2|500003586||4|2|500000294|-2||-2|7016|11|||7464|9|||1|500000294|0|4203557099934965158
M694|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|474|Red||2014-08-13|2014-08-22|2015-12-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||15.6||1|1|1|1|F|Black||14|No|Mother|28031|6|Two Parent|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||49|28115|High School Graduate|Single|Customer Service|28115|13|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503937201|503939209|31|0|2|503582646|1|0|2|500772180|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1||3974159976843499574|5113775940557498788
M695|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|49|Green||2017-01-12|2017-01-17|NaT||||1.6||2|2|2|2|M|White||14|No|GrandMother|28031|5|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|White||61|28202|Masters Degree|Married|Retired||0|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503913977|503915984|1|0|1|503898216|1|0|1|500939856|10|2|-2||2|1||-2||-2|0|4|||17101|1|||1||7581500809034284566|0
M696|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|680|Yellow||2014-06-24|2014-06-24|2016-05-04|Child: Family structure changed|Child: Family structure changed||22.3||2|2|2|2|M|White||14|No|GrandMother|28031|5|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|White||61|28202|Masters Degree|Married|Retired||0|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|503913977|503915984|1|0|1|503898216|1|0|1|500767515|10|2|-2||4|2||-2||-2|0|4|||17101|1|||1||7581500809034284566|0
M697|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-27|2016-11-02|NaT||||4.1||1|1|1|1|M|Black||14|No|Mother|28208|9|One Parent: Female|$20,000 to $24,999||||Yes||Relative|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||31|28226|Masters Degree|Married|Finance|28202|0|4|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504867822|504870341|31|0|1|504743932|1|0|1|500920611|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|3|||17159|12|||1||702163000107564368|0
M698|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|123|Green||2016-10-31|2016-11-04|NaT||||4||1|1|1|1|M|White||14|No|Mother|28216|9|Two Parent|$20,000 to $24,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||35|28270|Masters Degree|Married|Business: Engineer|76092|0|5|Self|Self|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504880135|504882655|1|0|1|504738710|1|0|1|500921982|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||7464|9|||1||702163000107564368|0
M699|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1376|Yellow||2013-05-14|2013-05-31|NaT||||45.2||2|2|1|1|F|Hispanic||14|No|Mother|28269|6|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Hispanic||41|28079|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|502829894|502831178|3|0|2|503443998|3|0|2|500696822|10|2|-2||2|2||-2||-2|0|4|||7464|9|||1||5441374193599827162|0
M700|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|137|Green||2016-09-20|2016-10-21|NaT||||4.5||1|1|1|1|M|White||14|No|Mother|28212|7|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|M|White||28|28205|Bachelors Degree|Single|Tech: Sales, Mktg|28202|3|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504574961|504577295|1|0|1|504676344|1|0|1|500908810|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||2811191761055817959|0
M701|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|206|Green||2014-11-06|2014-11-07|2015-06-01|Child: Lost interest|Child: Lost interest||6.8||2|2|2|2|M|Black||14|No|Mother|28208|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|Amachi, Project Big, Project Big AND Amachi|Match Support|M|White||27|29710|Bachelors Degree|Married|Business: Human Resources|28217|3|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|502549830|502550279|31|0|1|504035546|1|0|1|500792594|10|1|500009132|2128207319|4|1|500000294, 500004640, 500004901|-1||-1|0|4|||11247|3|||1||3935539763241716148|0
M702|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2077|Green|Amachi, Project Big, Project Big AND Amachi|2011-05-26|2011-06-30|NaT||||68.2||2|2|1|1|M|Black||14|No|Mother|28208|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|Amachi, Project Big, Project Big AND Amachi|Match Support|M|Black||25|28211||Single|Transport: Driver||0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502549830|502550279|31|0|1|502462453|31|0|1|500538768|10|2|500004772||2|1|500000294, 500004640, 500004901|-1||-2|0|4|||7464|9|||1|500000294, 500004640, 500004901|3935539763241716148|0
M703|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|462|Green||2014-12-18|2015-01-12|2016-04-18|Child: Family structure changed|Child: Family structure changed||15.2||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|White||30|28205|Bachelors Degree|Living w/ Significant Other|Finance: Banking|28217|3|4|Igniting Breakfast|Special Event|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500021785|502107146|502107573|31|0|1|504090344|1|0|1|500804987|10|2|-2||4|1||-2||-2|0|10|||17266|8|||1||4112464363801619560|7151546326379863072
M704|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|380|Yellow|PERL 2014-2016|2015-05-26|2015-06-16|2016-06-30|Child: Lost interest|Child: Lost interest||12.5||1|1|1|1|F|White||14|No|GrandMother|28277|7|Grandparents|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||30|28273|Bachelors Degree|Single|Business: Engineer|28273|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Enrollment|0|1|1|0|277|60|598|500000170|500013781|504221476|504223590|1|0|2|504231286|1|0|2|500828128|10|2|-2||4|2|500014681|-2|500014681|-2|0|5|||17159|12|||1|500014681|0|5605796235524810842
M705|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-27|2016-11-02|NaT||||4.1||1|1|1|1|M|Black||14|No|Mother|28217|9|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site|mentor2.0, mentor2.0 2016|Match Support|M|White||24|28202|Masters Degree|Single|Finance: Accountant|28202|0|9|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500022907|504831698|504834200|31|0|1|504751575|1|0|1|500920622|10|1|500014504||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||17159|12|||1||702163000107564368|0
M706|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|463|Green||2014-02-21|2014-03-12|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||15.2||1|1|3|3|M|Black||14|No|Mother|28206|6|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||29|28202|Masters Degree|Single|Business|28202|5|0|Duke Energy|Workplace Partner|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500016270|503690173|503692138|31|0|1|503604304|1|0|1|500750238|10|1|500009132|2128173561|4|1||-1|500000294|-1|0|4|||16705|3|||1||7960300212314874874|0
M707|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|238|Red||2016-05-04|2016-05-27|2017-01-20|Child: Severity of challenges|Child: Severity of challenges||7.8||1|1|1|1|M|Black||14|No|Mother|28215|7|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|M|White||23|28205|Bachelors Degree|Single|Finance|28210|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500008321|504318423|504320644|31|0|1|504561410|1|0|1|500891770|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||8568001799025358453|2141487034287122220
M708|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2315|Red|Amachi, Project Big, Project Big AND Amachi|2010-10-21|2010-10-28|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||76.1||1|1|1|1|F|Black||14|Yes|Mother|28269|4|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||35|28213|Masters Degree|Married|Business: Clerical||3|6|Radio|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502359051|502359489|31|0|2|502242295|31|0|2|500483954|10|2|500004772||4|3|500000294, 500004640, 500004901|-2||-2|0|10|||131|1|||1|500000294, 500004640, 500004901|540227296891876425|0
M709|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2598|Green|Amachi|2009-12-03|2010-01-25|NaT||||85.4||1|1|1|1|M|Black||14|Yes|Mother|28214|7|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||64|28117||Married|Business: Sales|28031|0|0|Alpha Kappa Alpha|Fraternity/Sorority|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501788776|501789128|31|0|1|501698382|1|0|1|500418170|10|2|500003586||2|1|500000294|-2||-2|0|10|||8697|14|||1|500000294|806697982905023857|0
M710|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1870|Yellow|Amachi|2012-01-04|2012-01-23|NaT||||61.4||1|1|2|2|F|Black||14|Yes|Mother|28273||One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28208|Some College|Single|Education: Teacher|28226|1|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|1|0|0|1|277|60|598|500000170|500008321|502825916|502827199|31|0|2|502367677|31|0|2|500589764|10|2|-2||2|2|500000294|-2|500000294, 500004640|-2|0|10|||7464|9|||1|500000294|6128289346130089489|0
M711|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|489|Red|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2015-04-11|2015-04-28|2016-08-29|Volunteer: Moved|Volunteer: Moved||16.1||1|1|1|1|M|Hispanic||14|No|Mother|28215|8|One Parent: Female|Unknown|||Y|Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Enrollment|M|Hispanic||27|28262|Some College|Single|Finance: Banking|28228|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|0|1|1|0|277|60|598|500000170|500017777|504154297|504156341|3|0|1|504201847|3|0|1|500822827|5|2|-2||4|3|500011312, 500014681|-2|500011312, 500014681|-2|0|10|||17159|12|||1|500011312, 500014681|6724463016047116758|0
M712|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|265|Green|PERL 2014-2016|2014-09-18|2014-09-25|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||1|1|2|3|M|Black||14|No|GrandMother|28269|5|Grandparents|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|Hispanic||34|28205|Masters Degree|Divorced|Tech: Engineer|28202|8|0|Duke Energy|Workplace Partner|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503999208|504001223|31|0|1|503973970|3|0|1|500776594|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-2|0|4|||16705|3|||1|500014681|7960300212314874874|0
M713|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1415|Green||2013-04-08|2013-04-22|NaT||||46.5||2|2|1|1|F|Hispanic||14|No|Mother|28262|9|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||43|28216|Masters Degree|Single|Finance: Accountant|28685|1|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502753873|502751081|3|0|2|503146044|31|0|2|500691867|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||7432163260389731024|0
M714|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|526|Green||2015-08-22|2015-09-28|NaT||||17.3||3|3|1|1|F|Black||14|No|Mother|28216|7|Two Parent|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||43|28269|Masters Degree|Single|Business: Mgt, Admin||0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502186245|501610196|31|0|2|504248899|1|0|2|500836970|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||6381341368426079638|7044657180546140448
M715|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1607|Red||2012-09-19|2012-09-30|2017-02-23|Volunteer: Time constraint|Volunteer: Time constraint||52.8||1|1|1|1|M|Black||14|Yes|Mother|28208|9|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Black||32|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|503016111|503013381|31|0|1|503135600|31|0|1|500636811|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||7496|10|||1||253338316288302752|5553585308107995803
M716|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1349|Green||2013-06-19|2013-06-27|NaT||||44.3||2|2|1|1|F|Black||14|No|Mother|28212|5|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28209|Masters Degree|Single|Medical|28207|0|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502436198|502436641|31|0|2|503255826|1|0|2|500701262|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1||0|6156547733130613405
M717|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|535|Red||2014-04-30|2014-05-09|2015-10-26|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17.6||3|3|2|2|F|Black||14|No|Mother|28227|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||30|28213|Some College|Single|Medical|28209|1|4|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500020990|503643026|503644986|31|0|2|503377601|31|0|2|500761779|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||1421169092898167719|0
M718|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|441|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2015-12-15|2015-12-22|NaT||||14.5||3|3|1|1|F|Black||14|No|Mother|28227|8|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||26|28202||Single|Consultant|28281|1|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|503643026|503644986|31|0|2|504315865|1|0|2|500867875|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|500007920, 500011315, 500011316|1421169092898167719|0
M719|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|435|Green||2014-10-27|2014-11-24|2016-02-02|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.3||2|2|1|1|F|Black||14|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Site||Enrollment|F|Black||25|28205|Some College|Married|Student: College||0|0|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503791020|503792997|31|0|2|503783913|31|0|2|500788555|5|1|500000295|2128173561|4|1||-1||-1|0|4|||7464|9|||1||702163000107564368|4127833823859005557
M720|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|866|Red||2013-02-21|2013-02-28|2015-07-14|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||28.5||1|1|1|1|M|Black||14|No|Mother|28213|K|One Parent: Female|$10,000 to $14,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||50|28269|Associate Degree|Married|Self-Employed, Entrepreneur||12|0|Newspaper|Media|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|501143676|501143950|31|0|1|503315012|31|0|1|500683363|10|2|-2||4|3||-2|500000294|-2|34|2|||129|1|||1||0|0
M721|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|984|Green||2014-06-10|2014-06-27|NaT||||32.3||1|1|1|1|M|Black||14|No|Mother|28227|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|Black||42|28270|Bachelors Degree|Married|Unknown||0|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503803127|503798593|31|0|1|503866013|31|0|1|500766041|10|2|-2||2|1||-2||-2|0|4|||17101|1|||1||7284449467126735125|7044657180546140448
M722|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|312|Green|PERL 2014-2016|2016-04-13|2016-04-29|NaT||||10.3||1|1|1|1|M|Black||14|No|Mother|28212|6|One Parent: Female|$35,000 to $39,999||||Yes|TV|Media|General Community|PERL 2014-2016|Match Support|M|White||35|28215|Some College|Living w/ Significant Other|Tech: Engineer|11735|1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504129013|504131049|31|0|1|504577506|1|0|1|500888874|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|56|1|||7496|10|||1|500014681|2811191761055817959|2197933814735019388
M723|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|48|Yellow|PERL 2014-2016|2015-05-21|2015-05-27|2015-07-14|Volunteer: Time constraint|Volunteer: Time constraint||1.6||2|2|1|1|M|American Indian or Alaska Native||14|No|Mother|28269|7|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||53|28027||Married|Tech: Management|28117|7|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500012459|504150667|504152735|6|0|1|503845717|1|0|1|500827880|10|2|-2||4|2|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681|3677730851176818072|3402014428779854546
M724|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|565|Green||2015-08-13|2015-08-20|NaT||||18.6||2|2|3|3|M|American Indian or Alaska Native||14|No|Mother|28269|7|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Asian||27|28202|Bachelors Degree|Single|Finance|28202|0|1|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500020752|504150667|504152735|6|0|1|504242094|4|0|1|500836074|10|2|-2||2|1|500014681|-2||-1|0|4|||17159|12|||1||3677730851176818072|3402014428779854546
M725|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|503|Green||2013-10-14|2013-11-13|2015-03-31|Child: Lost interest|Child: Lost interest||16.5||1|1|1|1|M|Black||14|No|Mother|28206|6|One Parent: Female|Unknown||||No||School|General Site||Match Support|M|White||39|28036|Masters Degree|Married|Business: Human Resources|28202|8|5|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503217134|503218915|31|0|1|503605778|1|0|1|500718993|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M726|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|268|Green||2014-09-04|2014-09-23|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||2|2|3|3|M|Black||14|No|Mother|28206|6|Two Parent|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||48|28216|Bachelors Degree|Married|Business: Engineer|28262|7|6|Recruitment Event|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503633782|503635723|31|0|1|502441938|31|0|1|500774542|10|1|500009132|2128173561|4|1||-1||-1|0|4|||7446|3|||1||7960300212314874874|0
M727|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|594|Green|PERL 2014-2016|2014-11-13|2014-11-25|2016-07-11|Child: Changed school/site|Child: Changed school/site||19.5||1|1|3|3|F|Multi-race (Black & Hispanic)||14|No|Mother|28217|8|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|Black||34|28273|Bachelors Degree|Single|Business: Mgt, Admin||5|0|LPL Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500015820|504089044|504091074|38|0|2|503255983|31|0|2|500795289|10|1|500009132|2128207319|4|1|500014681|-1|500014681|-1|0|4|||11247|3|||1|500014681|3935539763241716148|0
M728|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|848|Green||2013-09-25|2013-09-30|2016-01-26|Volunteer: Moved|Volunteer: Moved||27.9||1|1|3|3|F|Black||14|No|Mother|28217|7|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Black||34|28273|Bachelors Degree|Single|Retail: Mgt|28217|5|6|AA Task Force|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503524258|503526133|31|0|2|500497043|31|0|2|500713184|5|2|-2||4|1|500000294|-2||-2|34|2|||6247|12|||1||0|8662074432862573840
M729|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|135|Green||2015-09-23|2015-10-07|2016-02-19|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||4.4||1|1|3|3|F|Black||14|No|Aunt|28208|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Enrollment|F|White||28|28203|Bachelors Degree|Single|Finance|28202|0|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333730|504335952|31|0|2|504349844|1|0|2|500841754|5|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|8178900818136675730
M730|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|715|Green||2013-10-29|2013-11-18|2015-11-03|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||23.5||1|1|1|1|F|Black||14|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||30|28202|Bachelors Degree|Single|Business: Marketing|28202|0|2|Duke Energy|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503602213|503604090|31|0|2|503606038|1|0|2|500724439|10|1|500009132|2128173561|4|1||-1||-2|0|4|||16705|3|||1||7960300212314874874|0
M731|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|375|Yellow||2014-09-19|2014-09-26|2015-10-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.3||1|1|2|2|F|Black||14|No|Mother|28227|6|One Parent: Female|$20,000 to $24,999|Yes: Active|No|Y|Yes||Self|General Community||Match Support|F|Black||46|28216|Bachelors Degree|Single|Business: Marketing|28036|0|3|Self|Self|Big|General Community|VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500012459|503544893|503546768|31|0|2|503844843|31|0|2|500777054|10|2|-2||4|2||-2|500007920, 500011312, 500011315, 500011316|-2|0|10|||7464|9|||1||4112464363801619560|5468286809853673926
M732|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|470|Green||2015-01-23|2015-01-26|2016-05-10|Child/Family: Moved|Child/Family: Moved||15.4||1|1|1|1|M|Multi-race (Black & White)||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|M|White||30|28203|Masters Degree|Single|Finance: Banking|28262|4|4|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504054633|504056657|36|0|1|504068503|1|0|1|500809809|10|2|-2||4|1||-2||-2|0|4|||17159|12|||1||1421169092898167719|0
M733|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|423|Green||2014-05-14|2014-05-19|2015-07-16|Child/Family: Moved|Child/Family: Moved||13.9||3|3|2|2|F|Hispanic||14|Yes|Mother|28217|4|One Parent: Female|Unknown||||Yes||School|General Site|Amachi|Match Support|F|White||43|28031|Associate Degree|Single|Finance||4|0|Recruitment Event|BBBS Board/Staff|Big|General Site|Amachi|RTBM|1|0|1|0|277|60|598|500000170|500016847|502776307|502777486|3|0|2|502483716|1|0|2|500763275|10|1|500000295|2128173557|4|1|500000294|-1|500000294|-1|0|4|||7462|13|1204|3|1||8981704271528751143|0
M734|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1778|Green|Amachi|2012-04-10|2012-04-24|NaT||||58.4||2|2|1|1|F|Black||14|Yes|Relative: Other|28227|3|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||35|28277|Masters Degree|Single|Education: Admin||8|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502255156|502255582|31|0|2|502946412|1|0|2|500608992|10|2|500003586||2|1|500000294|-2||-2|0|5|||7462|13|||1|500000294|0|0
M735|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2035|Green|Project Big|2011-08-04|2011-08-11|NaT||||66.9||1|1|2|2|M|Black||14|No|Mother|28216|6|One Parent: Female|$30,000 to $34,999||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||48|28216|Bachelors Degree|Married|Finance: Banking|28255|8|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502529397|502529850|31|0|1|500188946|31|0|1|500548763|10|2|500004641||2|1||-2||-2|6854|8|||7464|9|||1|500004640|806697982905023857|0
M736|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|397|Green|PERL 2014-2016|2014-09-18|2014-09-25|2015-10-27|Volunteer: Time constraint|Volunteer: Time constraint||13||1|1|2|2|F|Hispanic||14|Yes|Mother|28206|7|One Parent: Female|Unknown|||Y|Yes||School|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Enrollment|F|Hispanic||41|28203||Single|Business|28202|2|6|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503999199|504001214|3|0|2|503973076|3|0|2|500776775|5|1|500000295|2128173561|4|1|500011312, 500014681|-2|500014681|-1|0|4|||16705|3|||1|500014681|7960300212314874874|0
M737|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|293|Green||2015-09-28|2015-10-08|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.6||1|1|3|3|M|Black||14|No|Mother|28208|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|M|Asian||27|28202|Bachelors Degree|Single|Finance|28202|0|1|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504348416|504350640|31|0|1|504242094|4|0|1|500842688|10|1|500009132|2128207318|4|1||-1||-1|0|4|||17159|12|||1||2611337051335117774|0
M738|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|621|Green||2014-07-09|2014-07-17|2016-03-29|Volunteer: Moved|Volunteer: Moved||20.4||1|1|1|1|M|Black||14|No|Mother|28212|7|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Enrollment|M|White||28|28270|Bachelors Degree|Married|Real Estate: Realtor|28203|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503479095|503480961|31|0|1|503915425|1|0|1|500768983|5|2|-2||4|1||-2||-2|0|10|||46|2|||1||8202428416367135871|7100264174759976571
M739|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1988|Red||2009-12-14|2009-12-18|2015-05-29|Child: Lost interest|Child: Lost interest||65.3||1|1|2|2|F|Black||14|No|Mother|28216|1|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||37|28078|Bachelors Degree|Single|Business: Human Resources|28226|0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501863951|501864324|31|0|2|501601161|31|0|2|500421259|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||0|0
M740|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|126|Green||2015-01-21|2015-01-21|2015-05-27|Child/Family: Moved|Child/Family: Moved||4.1||2|2|1|1|M|Black||14|No|Mother|28206|6|One Parent: Female|Unknown||||No||School|General Site|PERL 2014-2016|Match Support|F|White||39|28205|Bachelors Degree|Single|Tech: Research/Design|28202|0|5|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504013295|504015310|31|0|1|504146637|1|0|2|500809311|10|1|500009132|2128173561|4|1|500014681|-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M741|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|381|Green|Cabarrus County|2016-02-16|2016-02-20|NaT||||12.5||1|1|2|2|M|Multi-race (Asian & White)||14|No|Mother|28027|9|One Parent: Female|$60,000 to $74,999|||Y|No||Self|General Community|Cabarrus County|Match Support|M|Black||30|28213|Masters Degree|Single|Education|28217|0|7|Recruitment Event|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504545166|504547500|37|0|1|503788318|31|0|1|500879416|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7458|9|||1|500016374|4621676786129919860|6156547733130613405
M742|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1220|Yellow||2012-06-08|2012-06-19|2015-10-22|Volunteer: Moved|Volunteer: Moved||40.1||1|1|1|1|F|Black||14|No|Mother|28270|6|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Multi-Race (None of the above)||28|28215|Some College|Single|Insurance||0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503021552|503023091|31|0|2|502951522|7|0|2|500618601|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1||7284449467126735125|8145184518918286703
M743|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|518|Green||2015-09-22|2015-10-06|NaT||||17||1|1|3|3|M|American Indian or Alaska Native||14|No|Mother|28217|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||29|28202|Masters Degree|Single|Business|28202|5|0|Duke Energy|Workplace Partner|Big|General Site|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500021785|504396237|504398477|6|0|1|503604304|1|0|1|500841339|10|1|500009132|2128212899|2|1||-1|500000294|-1|0|4|||16705|3|||1||7276767778509034039|0
M744|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1265|Green||2013-09-11|2013-09-19|NaT||||41.6||1|1|1|1|F|Black||14|No|Mother|28214|6|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|Black||26|28209|Bachelors Degree|Single|Retail: Sales|28210|0|10|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503497835|503499703|31|0|2|503507978|31|0|2|500710423|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||806697982905023857|186501922587095434
M745|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|148|Green||2016-09-22|2016-10-10|NaT||||4.9||1|1|1|1|F|Black||14|No|Mother|28208|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|Native Hawaiian or Other Pacific Islander||22|28203|Bachelors Degree|Single|Tech: Computer/Programmer|28208|0|3|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504855816|504858318|31|0|2|504839044|5|0|2|500909638|10|1|500009132|2128212899|2|1||-1||-1|0|4|||7464|9|||1||8568001799025358453|0
M746|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|284|Green||2015-09-22|2015-10-01|2016-07-11|Volunteer: Time constraint|Volunteer: Time constraint||9.3||1|1|1|1|F|Black||14|No|Mother|28203|7|One Parent: Female|Unknown|||Y|Yes||School|General Site||Enrollment|F|White||24|28120|Bachelors Degree|Single|Business|28208|2|5|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504410234|504412485|31|0|2|504368847|1|0|2|500841344|5|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M747|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1043|Green||2014-04-17|2014-04-29|NaT||||34.3||1|1|1|1|M|Black||14|No|Mother|28216|4|One Parent: Female|$60,000 to $74,999|Yes: Active|Yes||No|AARTF|Neighbor/Friend|General Community||Match Support|M|White||27|28217|Masters Degree|Single|Finance|28202|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503429736|503431601|31|0|1|503850437|1|0|1|500760086|10|2|-2||2|1||-2||-2|6855|8|||17159|12|||1||2324686837245224089|8110690944529142441
M748|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-31|2016-10-31|NaT||||4.2||2|2|2|2|F|Black||14|No|Mother|28215|5|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|Black||28|28212|Masters Degree|Single|Customer Service|28202|3|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502943644|502945070|31|0|2|503671882|31|0|2|500922104|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||6368218764956286027|7674215580094440446
M749|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|431|Red||2014-08-07|2014-08-25|2015-10-30|Volunteer: Time constraint|Volunteer: Time constraint||14.2||2|2|1|1|F|Black||14|No|Mother|28215|5|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|Black||23|28213||Single|Arts, Entertainment, Sports||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502943644|502945070|31|0|2|503899413|31|0|2|500771637|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||6368218764956286027|7674215580094440446
M750|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|410|Yellow||2014-11-17|2014-11-24|2016-01-08|Child: Lost interest|Child: Lost interest||13.5||2|2|1|1|F|White||14|No|Mother|28031|4|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|F|White||31|28036|Associate Degree|Single|Medical|28202|6|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503166335|503168022|1|0|2|503729353|1|0|2|500796127|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||836952159905822963|4899162720666011799
M751|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|732|Red||2015-02-24|2015-02-26|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||24||2|2|1|1|F|Black||14|No|Mother|28215|3|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||42|28216|Associate Degree|Married|Business: Clerical|28202|8|0|Duke Energy|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502875279|502876679|31|0|2|504151222|31|0|2|500815521|10|2|-2||4|3||-2||-2|0|10|||16705|3|||1||7987165241089060600|0
M752|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|110|Green|PERL 2014-2016|2014-09-18|2014-09-25|2015-01-13|Child/Family: Moved|Child/Family: Moved||3.6||1|1|2|2|F|Black||14|No|Mother|28205||One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|F|Black||39|28025||Divorced|Business|28285|0|6|Duke Energy|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503999194|504001209|31|0|2|503611445|31|0|2|500776592|10|1|500009132|2128173561|4|1|500014681|-1||-1|0|4|||16705|3|||1|500014681|7960300212314874874|0
M753|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1630|Green||2012-08-31|2012-09-19|NaT||||53.6||1|1|1|1|F|Black||14|No|Mother|28214|8|One Parent: Female|$30,000 to $34,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|White||33|28207|Bachelors Degree|Married|Business||0|7|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500021785|503017622|503019155|31|0|2|503095382|1|0|2|500631726|10|2|-2||3|1||-2||-2|34|2|||7464|9|||1||421482027904269589|7992059899544338484
M754|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|434|Green|PERL 2014-2016|2015-03-02|2015-05-14|2016-07-21|Volunteer: Moved|Volunteer: Moved||14.3||1|1|1|1|M|White||14|No|Mother|28206|6|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|M|Black||50|29418|PHD|Separated|Business: Mgt, Admin|27713|0|2|Current/Previous Big|Other Big|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504172774|504174882|1|0|1|504040677|31|0|1|500816352|10|1|500000295|2128173561|4|1|500014681|-1|500014681|-1|0|4|||17159|12|||1|500014681|7960300212314874874|0
M755|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1804|Green||2012-03-12|2012-03-29|NaT||||59.3||1|1|1|1|F|Black||14|No|Mother|28215|8|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||54|28262|Bachelors Degree|Single|Business: Mgt, Admin||0|9|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502945480|502946906|31|0|2|502919780|31|0|2|500603409|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||5441374193599827162|7853254786544686064
M756|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3197|Green|Amachi|2008-05-28|2008-06-05|NaT||||105||1|1|1|1|M|Black||14|Yes|GrandMother|28208|8|One Parent: Female|Less than $10,000||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|M|White||53|28204|Juris Doctorate (JD)|Married|Law: Lawyer|28244|16|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|501142903|501143177|31|0|1|501236825|1|0|1|500268808|10|2|500003586||2|1|500000294|-2|500000294|-2|7294|13|||2238|7|||1|500000294|7276767778509034039|0
M757|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2520|Red|Amachi|2009-07-22|2009-07-24|2016-06-17|Volunteer: Moved|Volunteer: Moved||82.8||2|2|1|1|F|Multi-Race (None of the above)||14|No|Mother|28211|7|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||50|28227|Some College|Single|Human Services: Social Worker||2|5|St. Paul Baptist|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501721579|501721919|7|0|2|501687513|31|0|2|500375006|10|2|500003586||4|3|500000294|-2|500000294|-2|5635|9|||9609|7|||1|500000294|2811191761055817959|0
M758|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1006|Green||2014-05-08|2014-06-05|NaT||||33.1||1|1|2|2|M|Black||14|No|Mother|28206|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||66|28269||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503381531|503383388|31|0|1|500540549|31|0|1|500762593|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||392688197545050058|5081726734274569781
M759|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|268|Green||2014-09-04|2014-09-23|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||2|2|3|3|M|Black||14|No|Mother|28205|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||29|28273|Bachelors Degree|Married|Tech: Computer/Programmer||5|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503690154|503692119|31|0|1|502542324|31|0|1|500774537|10|1|500009132|2128173561|4|1||-1|500014681|-1|0|4|||16705|3|||1||7960300212314874874|0
M760|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-25|2015-10-01|NaT||||17.2||1|1|3|3|F|Black||14|No|Mother|28209|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|Black||36|28269||Single|Business|28202|7|5|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504396225|504398465|31|0|2|503605618|31|0|2|500842435|10|1|500009132|2128212899|2|1||-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M761|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|148|Green||2016-09-20|2016-10-10|NaT||||4.9||2|2|2|2|F|Black||14|No|Mother|28203|8|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||25|28202|Bachelors Degree|Single|Tech: Computer/Programmer|28208|2|1|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504410165|504412416|31|0|2|504445343|1|0|2|500908999|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M762|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|279|Green||2015-09-22|2015-10-06|2016-07-11|Volunteer: Time constraint|Volunteer: Time constraint||9.2||2|2|1|1|F|Black||14|No|Mother|28203|8|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||25|28203|Bachelors Degree|Single|Consultant|28202|2|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504410165|504412416|31|0|2|504403681|1|0|2|500841641|10|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M763|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|223|Green||2015-11-13|2015-12-17|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||7.3||1|1|1|1|M|Black||14|Yes|Mother|28208|6|One Parent: Female|Less than $10,000||||Yes||School|General Site|PERL 2014-2016|Match Support|M|White||26|28027|Masters Degree|Single|Finance: Auditor|28202|0|4|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500016270|504416580|504418832|31|0|1|504504983|1|0|1|500859759|10|1|500009132|2128207318|4|1|500014681|-1|500007920, 500011315, 500011316, 500014681|-1|0|4|||12831|3|||1||2611337051335117774|0
M764|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1350|Green||2013-06-11|2013-06-26|NaT||||44.4||3|3|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||39|28211||Single|Retail: Sales||0|11|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501721762|501722098|31|0|2|503471102|31|0|2|500700196|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||1227369534771287213|0
M765|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1127|Yellow||2012-06-11|2012-06-25|2015-07-27|Volunteer: Time constraint|Volunteer: Time constraint||37||2|2|1|1|M|Black||14|No|Mother|28208|6|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||31|28210|Bachelors Degree|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|501721761|501722098|31|0|1|503023854|1|0|1|500618753|7|2|-2||4|2||-2||-2|0|10|||7464|9|||1||1227369534771287213|0
M766|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1627|Red||2010-08-04|2010-08-17|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||53.5||1|1|1|1|M|Black||14|No|Mother|28212|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||50|28212|Some College|Married|Law: Police Officer||2|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|502236953|502237384|31|0|1|502232559|31|0|1|500464143|10|2|-2||4|3||-2|500000294|-2|0|10|||7464|9|||1||2811191761055817959|0
M767|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|268|Green||2014-09-18|2014-09-23|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|2|2|F|Black||14|No|Father|28208|6|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|F|White||30|28203|Bachelors Degree|Single|Business|28202|1|3|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504013291|504015306|31|0|2|503979108|1|0|2|500776595|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M768|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|359|Green|PERL 2014-2016|2015-04-30|2015-05-19|2016-05-12|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||11.8||1|1|1|1|M|Black||14|No|Mother|28227|6|One Parent: Female|$10,000 to $14,999||||Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Black||33|28215|Associate Degree|Single|Business|28202|0|3|Self|Self|Big|General Community|PERL 2014-2016|Enrollment|0|1|1|0|277|60|598|500000170|500020990|503941174|503943182|31|0|1|503207130|31|0|1|500825477|10|2|-2||4|1|500014681|-2|500014681|-2|0|5|||7464|9|||1|500014681|2728869331911165614|7312235294346727700
M769|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1984|Green||2010-11-10|2010-12-03|2016-05-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||65.2||1|1|1|1|F|Black||14|No|Mother|28208||One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|F|White||35|28210|Bachelors Degree|Living w/ Significant Other|Business: Sales|18034|2|7|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big AND Amachi|Match Support|1|0|1|0|277|60|598|500000170|500021785|502308197|502308629|31|0|2|502325667|1|0|2|500493122|5|2|500003586||4|1|500000294|-2|500000294, 500004901|-2|0|10|||7496|10|||1||0|0
M770|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1585|Yellow||2012-06-15|2012-06-30|2016-11-01|Child: Severity of challenges|Child: Severity of challenges||52.1||1|1|1|1|F|White||14|No|Mother|28210|6|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||33|28277|Bachelors Degree|Single|Consultant|28202|1|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|502506397|502506846|1|0|2|503039829|1|0|2|500619509|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||2272605169937511837|0
M771|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|666|Yellow|PERL 2014-2016|2015-05-11|2015-05-11|NaT||||21.9||2|2|3|3|M|Black||14|No|Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|Black||26|29730|Some High School|Married|Business: Sales|28217|1|6|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504057301|503680204|31|0|1|503796968|31|0|1|500826411|10|1|500000295|2128207319|2|2|500014681|-1||-1|0|4|||46|2|||1|500014681|3935539763241716148|0
M772|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|80|Green|PERL 2014-2016|2014-10-06|2014-11-03|2015-01-22|Child: Changed school/site|Child: Changed school/site||2.6||2|2|3|3|M|Black||14|No|Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|Black||26|29730|Some High School|Married|Business: Sales|28217|1|6|BBBS National Site|Web Link|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|504057301|503680204|31|0|1|503796968|31|0|1|500780724|10|1|500000295|2128207319|4|1|500014681|-1||-1|0|4|||46|2|||1|500014681|3935539763241716148|0
M773|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|156|Red||2015-05-04|2015-05-04|2015-10-07|Child/Family: Moved|Child/Family: Moved||5.1||1|1|1|1|M|Black||14|Yes|Mother|28216|5|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Enrollment|M|Black||37|28213|Some College|Living w/ Significant Other|Self-Employed, Entrepreneur|28206|2|0|Current/Previous Big|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500013781|502821218|502822501|31|0|1|504244628|31|0|1|500825744|5|2|-2||4|3||-2||-2|0|10|||17159|12|||1||7883015200677941272|6971797047831566199
M774|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|707|Green||2015-03-14|2015-03-31|NaT||||23.2||1|1|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Business: Sales|28277|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501843066|501843435|31|0|2|504152982|1|0|2|500818696|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||932861092942387634|0
M775|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|127|Red|PERL 2014-2016|2016-01-15|2016-01-31|2016-06-06|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||4.2||1|1|1|1|M|Black||14|No|Mother|28212|6|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Enrollment|M|White||38|28227|Some College|Single|Business: Sales||3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500013781|504076403|504078432|31|0|1|504415946|1|0|1|500872171|5|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||17159|12|||1|500014681|8758769076374727509|7044657180546140448
M776|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1775|Yellow|2010-2012 OJJDP JJI|2011-09-29|2011-10-13|2016-08-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||58.3||1|1|1|1|M|Black||14|No|Mother|28226|2|One Parent: Female|Less than $10,000||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||71|28277|Bachelors Degree|Married|Retired||0|0||Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502507408|502507857|31|0|1|502673562|31|0|1|500559678|10|2|-2||4|2||-2||-2|34|2|||0|11|||1|500005291|3539543368195872575|0
M777|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|235|Green||2015-01-21|2015-02-12|2015-10-05|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||7.7||1|1|4|4|F|Black||14|Yes|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|F|Multi-race (Black & White)||23|28273|Some College|Single|Student: College|28227|0|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500016270|504170222|504172330|31|0|2|503853917|36|0|2|500809356|5|1|500000295|2128173561|4|1||-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7464|9|||1||7960300212314874874|0
M778|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1803|Green||2012-03-13|2012-03-30|NaT||||59.2||2|2|1|1|F|Black||14|No|Mother|28216|7|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||31|28078|Bachelors Degree||Medical||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501295538|500740560|31|0|2|502897530|1|0|2|500603727|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||9134125726462845918|0
M779|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|654|Green||2014-03-12|2014-03-31|2016-01-14|Child: Lost interest|Child: Lost interest||21.5||1|1|1|1|F|Black||14|No|Mother|28215|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||29|28270||Single|Unemployed||0|0|Self|Self|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500020990|503756716|503758688|31|0|2|503596238|31|0|2|500754325|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||3723482195151978288|7665592423399355114
M780|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|505|Green||2015-02-24|2015-03-16|2016-08-02|Volunteer: Moved|Volunteer: Moved||16.6||1|1|1|1|F|Black||14|No|Mother|28213|6|One Parent: Female|$40,000 to $44,999||||Yes|BBBS National Site|Web Link|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|F|Black||23|28262|Some College|Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504038196|504040273|31|0|2|504062905|31|0|2|500815275|7|2|-2||4|1|500007920, 500011315, 500011316|-2||-2|34|2|||17159|12|||1||932861092942387634|8408514790530965815
M781|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|672|Green||2015-04-22|2015-05-05|NaT||||22.1||1|1|1|1|M|White||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999||||Yes||School|General Community||Match Support|M|White||51|28173|Masters Degree|Married|Self-Employed, Entrepreneur|28173|19|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504235369|504237484|1|0|1|503937954|1|0|1|500824366|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||1421169092898167719|8961132295198487522
M782|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2232|Green||2011-01-07|2011-01-26|NaT||||73.3||1|1|1|1|M|White||14|No|Mother|28277|4|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||67|28277|Bachelors Degree|Divorced|Tech: Sales, Mktg||0|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500017732|502225378|502225809|1|0|1|502245842|1|0|1|500509780|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||3090721985630916616|0
M783|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|169|Red||2015-11-10|2015-12-07|2016-05-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.6||1|1|1|1|M|Black||14|No|Mother|28027|7|One Parent: Female|$25,000 to $29,999||||Yes||School|General Community||Match Support|M|White||24|28262||Single|Medical: Healthcare Worker|28025|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020753|502129820|502130249|31|0|1|504474407|1|0|1|500858150|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||6353565629814722343|2881622112345502539
M784|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|517|Red||2013-08-06|2013-08-22|2015-01-21|Volunteer: Time constraint|Volunteer: Time constraint||17||1|1|1|1|M|Black||14|No|Mother|28211|4|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|Black||41|28216|Bachelors Degree|Single|Customer Service|28262|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503452963|503430105|31|0|1|503489818|31|0|1|500705904|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1||4903779310522421428|3402014428779854546
M785|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Green||2014-05-09|2014-05-16|2016-10-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||29||1|1|1|1|M|Black||14|Yes|Mother|28216|5|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|Black||54|28277|Bachelors Degree|Single|Consultant|28202|7|6|Man Up Campaign|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|1|0|1|0|277|60|598|500000170|500020910|503717073|503719040|31|0|1|503853194|31|0|1|500762798|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|4|||17101|1|||1||4863631750424600365|0
M786|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|680|Green||2013-11-19|2013-11-20|2015-10-01|Child: Graduated|Child: Graduated||22.3||1|1|6|6|F|Black||14|No|Mother|28083||Two Parent|Unknown||||Yes||School|General Site||Match Support|F|Black||38|28269|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500012459|503652810|503654770|31|0|2|500189256|31|0|2|500732404|10|1|500000295|2128212919|4|1||-1|500007920, 500011315, 500011316, 500016374|-1|0|4|||7464|9|1360|3|1||2437132833506538679|0
M787|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1084|Green||2014-03-04|2014-03-19|NaT||||35.6||2|2|1|1|F|Black||14|No|Mother|28216|4|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||35|27713|Associate Degree|Single|Business|28216|0|8|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|502336272|502336707|31|0|2|503743688|31|0|2|500752685|10|2|-2||2|1||-2||-2|6854|8|||7464|9|||1||3664007741235143067|6085623597595523017
M788|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1833|Yellow|Amachi|2010-04-14|2010-04-30|2015-05-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||60.2||2|2|2|3|F|Black||14|Yes|GrandMother|28227||Grandparents|Unknown||||No||Self|General Community|Amachi|Enrollment|F|Black||53|28269|Some College|Married|Business: Sales|28227|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500012459|501222138|501222414|31|0|2|500189173|31|0|2|500447311|5|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294|0|0
M789|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|868|Green||2014-10-03|2014-10-13|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||28.5||1|1|2|2|F|Black||14|Yes|Mother|28278|8|One Parent: Female|$50,000 to $59,999|||Y|No||Self|General Community||Match Support|M|Black||46|28214|Bachelors Degree|Single|Finance: Economist|28217|14|0|Brochure|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503972507|503974518|31|0|2|500189600|31|0|1|500780309|10|2|500003586||4|1||-2||-2|0|10|||127|1|||1||8567789404096574827|5746835512589871315
M790|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|2366|Green||2010-07-26|2010-08-03|2017-01-24|Volunteer: Time constraint|Volunteer: Time constraint||77.7||1|1|1|1|F|Black||14|No|Mother|28216|5|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|F|White||36|28208|Masters Degree|Single|Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|502222545|502222979|31|0|2|502196116|1|0|2|500462566|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1||1653226628427425023|0
M791|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2353|Green||2010-09-14|2010-09-27|NaT||||77.3||1|1|1|1|M|Black||14|No|Mother|28214|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||29|28210|Bachelors Degree|Married|Business: Mgt, Admin|97224|6|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020752|502255210|500910307|31|0|1|502255794|1|0|1|500470233|10|2|-2||2|1||-2|500000294|-2|0|10|||7496|10|||1||6381341368426079638|0
M792|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3080|Green||2008-08-15|2008-09-23|2017-02-28|Volunteer: Moved|Volunteer: Moved||101.2||1|1|1|1|F|Black||14|No|Mother|28230|8|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||34|28205|Masters Degree|Single|Finance: Banking|28217|0|4|Yahoo!|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501254255|501254531|31|0|2|501356688|1|0|2|500282157|10|2|-2||4|1||-2|500000294|-2|0|10|||32|2|||1||4440360203097874486|0
M793|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|665|Green||2014-09-12|2014-09-25|2016-07-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||21.8||1|1|3|3|F|Black||14|Yes|Mother|28206|6|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||36|28209|Masters Degree|Married|Business: Marketing|28202|0|4|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504007361|504009376|31|0|2|503605824|1|0|2|500775716|10|1|500000295|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M794|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|264|Green|PERL 2014-2016|2016-05-27|2016-06-16|NaT||||8.7||1|1|1|1|F|Multi-Race (None of the above)||14|No|Mother|28215|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Black||26|28262|Bachelors Degree|Single|Journalist/Media|28206|2|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504507791|504510086|7|0|2|504650231|31|0|2|500895078|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500014681|3148273126074974335|7044657180546140448
M795|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|130|Red|PERL 2014-2016, Cabarrus County|2016-10-21|2016-10-28|NaT||||4.3||1|1|4|4|F|Black||14|No|Mother|28027|6|Two Parent|$60,000 to $74,999|||Y|No|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Multi-race (Black & White)||23|28273|Some College|Single|Student: College|28227|0|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504655474|504657901|31|0|2|503853917|36|0|2|500918496|10|2|500016307||2|3|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||7464|9|||1|500014681, 500016374|4621676786129919860|7048951337647301192
M796|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1840|Green||2012-02-13|2012-02-22|NaT||||60.5||1|1|1|1|M|Black||14|No|Mother|28212|5|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||30|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502197486|502197915|31|0|1|502870668|1|0|1|500597982|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||7554307376683929204|8113241890313112769
M797|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|879|Green|PERL 2014-2016|2014-09-15|2014-10-10|NaT||||28.9||1|1|1|1|M|Black||14|Yes|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community|Amachi, PERL 2014-2016|Match Support|M|White||28|28209|Bachelors Degree|Single|Tech: Engineer||0|5|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020752|503953654|503955662|31|0|1|503976139|1|0|1|500775808|10|2|-2||2|1|500000294, 500014681|-2|500014681|-2|0|5|||46|2|||1|500014681|0|7044657180546140448
M798|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2400|Green||2010-08-03|2010-08-11|NaT||||78.9||1|1|1|1|F|Hispanic||14|No|Mother|28212|2|One Parent: Female|Unknown|||Y|No|Spanish Radio|Media|General Community||Match Support|F|White||33|28209||Single|Education: Teacher||0|0||High School Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|502255223|502255655|3|0|2|501823103|1|0|2|500463922|10|2|-2||2|1||-2||-2|7068|1|||0|4|||1||0|0
M799|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|88|Green||2015-10-07|2015-11-06|2016-02-02|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||2.9||2|2|1|1|F|Black||14|No|GrandFather|28205|7|One Parent: Female|Unknown||||No||School|General Site||RTBM|F|Black||26|28079|Some College|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|503217214|503218995|31|0|2|504373953|31|0|2|500845329|7|1|500000295|2128173561|4|1||-1||-1|0|4|||7496|10|||1||7960300212314874874|0
M800|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|684|Green||2013-04-16|2013-04-26|2015-03-11|Volunteer: Moved|Volunteer: Moved||22.5||2|2|1|1|F|Black||14|No|GrandFather|28205|7|One Parent: Female|Unknown||||No||School|General Site||RTBM|F|Black||24|28262|Some College|Single|Business|28202|0|5|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503217214|503218995|31|0|2|503350133|31|0|2|500693021|7|1|500000295|2128173561|4|1||-1||-1|0|4|||7464|9|||1||7960300212314874874|0
M801|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|211|Yellow||2014-10-14|2014-10-28|2015-05-27|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||6.9||3|3|1|1|F|Black||14|No|GrandMother|28215|8|Grandparents|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|F|Black||50|28215|Associate Degree|Married|Medical: Nurse||2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502583662|502584168|31|0|2|503943422|31|0|2|500783380|10|2|-2||4|2||-2||-2|0|4|||7464|9|||1||4112464363801619560|3959612471441160400
M802|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|541|Green||2015-08-20|2015-09-13|NaT||||17.8||3|3|1|1|F|Black||14|No|GrandMother|28215|8|Grandparents|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|F|White||23|28202||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502583662|502584168|31|0|2|504286292|1|0|2|500836763|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||4112464363801619560|3959612471441160400
M803|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|589|Yellow||2014-09-15|2014-10-06|2016-05-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.4||2|2|1|1|F|Black||14|No|GrandMother|28215|8|Grandparents|$30,000 to $34,999|||Y|Yes||School|General Community||RTBM|F|White||35|28205|Masters Degree|Single|Education: Teacher|28273|3|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|502583660|502584168|31|0|2|503944507|1|0|2|500775919|7|2|500003586||4|2||-2|500000294|-2|0|4|||46|2|||1||4112464363801619560|3959612471441160400
M804|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|469|Green|PERL 2014-2016|2015-04-07|2015-04-20|2016-08-01|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||15.4||1|1|1|1|M|Black||14|No|Mother|28215|6|One Parent: Female|$15,000 to $19,999||||Yes||Relative|General Community|PERL 2014-2016|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Engineer||0|2|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500020752|503679979|503226552|31|0|1|504191848|1|0|1|500822162|10|2|-2||4|1|500014681|-2|500014681|-2|0|3|||7464|9|||1|500014681|2728869331911165614|0
M805|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|518|Green||2015-10-06|2015-10-06|NaT||||17||1|1|2|2|F|Hispanic||13|No|Mother|28217|8|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|Hispanic||41|28203||Single|Business|28202|2|6|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504410212|504412463|3|0|2|503973076|3|0|2|500844559|10|1|500009132|2128212899|2|1||-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M806|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|260|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-23|2016-06-20|NaT||||8.5||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28213|7|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|Asian||25|28204|Bachelors Degree|Single|Finance|28215|0|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504691840|504694268|36|0|1|504535890|4|0|1|500894068|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1|500007920, 500011315, 500011316|3677730851176818072|8773162532572605235
M807|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1832|Green|Project Big|2012-02-17|2012-03-01|NaT||||60.2||1|1|2|2|M|Black||13|No|Mother|28213|2|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||40|28269||Married|Business: Marketing||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|502278985|502279417|31|0|1|500220237|31|0|1|500599107|10|2|-2||2|1||-2|500000294|-2|6854|8|||2238|7|||1|500004640|6065435025527210335|7044657180546140448
M808|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|837|Green||2014-11-12|2014-11-21|NaT||||27.5||1|1|2|2|M|Black||13|No|Mother|28079|5|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||45|28079|Bachelors Degree|Married|Business||13|6|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500017732|503552606|503554481|31|0|1|501052547|31|0|1|500794702|10|2|-2||2|1||-2|500000294|-2|0|10|||7671|13|||1||4575902950186762737|3402014428779854546
M809|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|106|Green|Cabarrus County|2016-11-18|2016-11-21|NaT||||3.5||1|1|1|1|M|Black||13|No|Mother|28025|7|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|Cabarrus County|Match Support|M|Black||29|28027|Bachelors Degree|Married|Business||0|10|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504732530|504734976|31|0|1|504893030|31|0|1|500929513|10|2|-2||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|5|||7464|9|||1|500016374|6750834084344455219|7044657180546140448
M810|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|434|Yellow||2014-05-21|2014-05-29|2015-08-06|Volunteer: Time constraint|Volunteer: Time constraint||14.3||1|1|1|1|M|Black||13|No|Mother|28227|7|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Enrollment|M|White||55|28031|Bachelors Degree|Separated|Business: Sales|53964|3|3|Local Print|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|503755565|503757537|31|0|1|503814505|1|0|1|500763994|5|2|-2||4|2||-2||-2|0|10|||7439|1|||1||7883015200677941272|2075602243867411528
M811|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|266|Green|PERL 2014-2016|2014-09-18|2014-09-23|2015-06-16|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||2|2|1|1|F|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Community|PERL 2014-2016|Match Support|F|White||28|28202|Bachelors Degree|Single|Business|28202|3|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|504013056|504015071|31|0|2|503976618|1|0|2|500776602|10|1|500009132|2128173561|4|1|500014681|-2|500014681|-1|0|4|||16705|3|||1|500014681|7960300212314874874|0
M812|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|532|Green|PERL 2014-2016|2015-09-13|2015-09-22|NaT||||17.5||2|2|1|1|F|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Community|PERL 2014-2016|Match Support|F|White||26|28202|Bachelors Degree|Single|Finance: Banking|28262|1|7|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|504013056|504015071|31|0|2|504219921|1|0|2|500839610|10|2|-2||2|1|500014681|-2||-2|0|4|||17159|12|||1|500014681|7960300212314874874|0
M813|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1011|Green||2014-05-16|2014-05-31|NaT||||33.2||1|1|1|1|F|Black||13|No|Mother|28269|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||59|28209|Bachelors Degree|Divorced|Medical|28209|1|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503632799|503634738|31|0|2|503567146|1|0|2|500763613|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||3677730851176818072|8242487816501170810
M814|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|531|Green||2013-10-02|2013-10-24|2015-04-08|Volunteer: Moved|Volunteer: Moved||17.4||2|2|1|1|M|Black||13||GrandMother|28213|3|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||42|28212|Bachelors Degree|Married|Arts, Entertainment, Sports|28202|2|11|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|501332660|501332937|31|0|1|503579743|31|0|1|500715179|10|2|-2||4|1|500000294|-2||-2|6854|8|||7464|9|||1||0|0
M815|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|286|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-11|2016-05-25|NaT||||9.4||2|2|1|1|M|Black||13||GrandMother|28213|3|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||26|28205|Bachelors Degree|Married|Real Estate: Realtor|28202|0|2|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|501332660|501332937|31|0|1|504556335|1|0|1|500892769|10|2|-2||2|1|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||17159|12|||1|500007920, 500011315, 500011316|0|0
M816|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1667|Red|Cabarrus County|2012-08-06|2012-08-13|NaT||||54.8||1|1|1|1|M|Hispanic||13|No|Mother|28027|7|One Parent: Female|$25,000 to $29,999||||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||33|28036|Bachelors Degree|Married|Business||2|5|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502605331|502605848|3|0|1|503090281|1|0|1|500627504|10|2|500016307||2|3|500016374|-2|500016374|-2|34|2|||7464|9|||1|500016374|6353565629814722343|3120960401464324192
M817|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|295|Green||2015-09-23|2015-10-07|2016-07-28|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|2|2|M|Black||13|No|Mother|28208|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|White||32|28262|Masters Degree|Married|Business: Mgt, Admin|28202|6|0|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504348425|504350649|31|0|1|503911472|1|0|1|500841772|10|1|500009132|2128207318|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1||2611337051335117774|0
M818|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3024|Green||2008-11-04|2008-11-25|NaT||||99.4||1|1|1|1|M|Black||13|No|Mother|28078||One Parent: Female|Unknown||||No||Relative|General Community||Match Support|M|Black||45|28262|Bachelors Degree|Married|Business: Mgt, Admin||0|6|AA Task Force|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501252806|501253082|31|0|1|501320197|31|0|1|500310204|10|2|-2||2|1||-2||-2|0|3|||6247|12|||1||0|0
M819|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|505|Green||2015-09-22|2015-10-19|NaT||||16.6||1|1|1|1|M|Black||13|No|Mother|28208|8|Two Parent|Unknown|||Y|Yes||School|General Site||Match Support|M|White||33|28278|Masters Degree|Married|Finance: Accountant|28202|1|2|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504416818|504419070|31|0|1|503988229|1|0|1|500841338|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M820|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|772|Green||2013-11-13|2013-11-25|2016-01-06|Child/Family: Moved|Child/Family: Moved||25.4||1|1|1|1|F|Black||13|No|Mother|28217|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||25|28134|Some College|Single|Child/Day Care Worker||0|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503617980|503619857|31|0|2|503573243|1|0|2|500730441|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1||4440360203097874486|634104847858773916
M821|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1251|Green||2013-09-18|2013-09-26|2017-02-28|Child: Family structure changed|Child: Family structure changed||41.1||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28214|4|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|Black||49|28273|Associate Degree|Single|Finance: Accountant|28273|7|0|Agency Sponsored|Special Event|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|503421607|503423471|36|0|2|503520561|31|0|2|500711787|10|2|-2||4|1||-2|500000294|-2|0|10|||16426|8|||1||7857548027029642592|1209912115202285875
M822|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|571|Green||2015-07-22|2015-08-14|NaT||||18.8||1|1|1|1|M|Black||13|No|Mother|28273|6|One Parent: Female|$35,000 to $39,999||||No||Self|General Community||Match Support|M|Black||56|28273|Some College|Married|Govt|28228|0|7|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|504284556|504286757|31|0|1|504260574|31|0|1|500834204|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||8567789404096574827|2392572474128905139
M823|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|789|Green||2014-11-25|2015-01-08|NaT||||25.9||1|1|1|1|M|Multi-race (Black & White)||13|Yes|Aunt|28031|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|Amachi|Match Support|M|White||51|28031|Masters Degree|Married|Real Estate: Realtor|28031|2|0|Local TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503654364|503656324|36|0|1|504076011|1|0|1|500799134|10|2|-2||2|1|500000294|-2||-2|0|4|||7438|1|||1||3974159976843499574|6178126991714892144
M824|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3015|Yellow||2008-11-17|2008-12-04|NaT||||99.1||1|1|1|1|M|Black||13|No|Mother|28217|K|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||39|28134|Bachelors Degree|Single|Business: Mgt, Admin||6|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501314104|501314382|31|0|1|501170940|1|0|1|500315948|10|2|-2||2|2||-2||-2|0|10|||7464|9|||1||0|6156547733130613405
M825|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|294|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-04-13|2016-05-17|NaT||||9.7||1|1|1|1|M|Black||13|No|Mother|28213|8|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|Black||27|28215|Bachelors Degree|Single|Tech: Computer/Programmer|28270|2|1|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500013781|503917550|503962680|31|0|1|504577899|31|0|1|500888953|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|500007920, 500011315, 500011316|5441374193599827162|6084148439133243542
M826|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|267|Green||2014-09-12|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|1|1|M|Black||13|No|Aunt|28205|6|Other Relative|Unknown||||Yes||School|General Site||Match Support|M|White||58|28211|Masters Degree|Married|Business|28202|7|0|Ally Financial|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|504013304|504015319|31|0|1|503910182|1|0|1|500775704|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M827|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-07|2016-10-31|NaT||||4.2||1|1|1|1|M|Black||13|No|Mother|28215|7|One Parent: Female|$40,000 to $44,999||||Yes||Self|General Community||Match Support|M|Multi-race (Hispanic & White)||28|28205|Bachelors Degree|Married|Finance: Banking|28202|1|4|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504564027|504566361|31|0|1|504766711|35|0|1|500913521|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||0|2806833304218536184
M828|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|253|Green||2014-06-26|2014-06-30|2015-03-10|Volunteer: Moved|Volunteer: Moved||8.3||2|2|1|1|F|Black||13|No|Mother|28215|3|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Enrollment|F|White||27|28203|Bachelors Degree|Single|Finance: Banking|28211|2|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500011349|501662033|501090456|31|0|2|503655814|1|0|2|500767861|5|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||0|4753237757252407321
M829|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-31|2016-10-31|NaT||||4.2||2|2|2|2|F|Black||13|No|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||37|28078|Bachelors Degree|Single|Business: Human Resources|28226|0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503977573|503980164|31|0|2|501601161|31|0|2|500922173|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||4440360203097874486|0
M830|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|336|Red|PERL 2014-2016|2014-12-04|2014-12-29|2015-11-30|Volunteer: Moved|Volunteer: Moved||11||2|2|1|1|F|Black||13|No|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||29|28277|Bachelors Degree|Single|Business: Clerical|28202|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500008321|503977573|503980164|31|0|2|504047655|31|0|2|500801295|10|2|-2||4|3||-2|500014681|-2|0|10|||17159|12|||1|500014681|4440360203097874486|0
M831|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1124|Green||2014-01-17|2014-01-31|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||36.9||1|1|1|1|F|Black||13|No|Mother|28216|5|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503662377|503664337|31|0|2|503573326|1|0|2|500743531|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||3664007741235143067|7044657180546140448
M832|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-21|2015-10-01|NaT||||17.2||1|1|2|2|F|Hispanic||13|No|Mother|28203|8|Two Parent|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||30|28203|Bachelors Degree|Single|Business|28202|1|3|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504410257|504412508|3|0|2|503979108|1|0|2|500841081|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M833|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|126|Green||2016-10-18|2016-11-01|NaT||||4.1||2|3|1|1|F|Black||13|No|Mother|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|Native Hawaiian or Other Pacific Islander||22|28209|Bachelors Degree|Single|Tech: Computer/Programmer|28202|0|2|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504401898|504404140|31|0|2|504875613|5|0|2|500917108|10|1|500009132|2128212899|2|1||-2||-1|0|4|||7464|9|||1||7276767778509034039|0
M834|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1619|Green||2012-07-26|2012-09-30|NaT||||53.2||1|1|1|1|F|Hispanic||13|No|Mother|28277|5|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||31|28210|Bachelors Degree|Single|Education: Teacher|29710|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503052850|503027860|3|0|2|503028888|1|0|2|500626321|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||3090721985630916616|8598768071652363430
M835|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|463|Yellow|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2015-11-17|2015-11-30|NaT||||15.2||1|1|2|2|F|Hispanic||13|No|Mother|28205|6|Two Parent|Unknown||||Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504331538|504333760|3|0|2|503843020|3|0|2|500860738|10|2|-2||2|2|500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500011312, 500014681|8758769076374727509|0
M836|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-22|2015-10-01|NaT||||17.2||1|1|1|1|M|Hispanic||13|No|Mother|28210|6|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|PERL 2014-2016|Match Support|M|White||27|28202|Bachelors Degree|Single|Finance|28208|2|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504439764|504442020|3|0|1|504392917|1|0|1|500841644|10|1|500009132|2128212899|2|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M837|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|409|Green||2014-09-11|2014-09-15|2015-10-29|Child/Family: Moved|Child/Family: Moved||13.4||1|1|1|1|F|Black||13|No|Mother|28227|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||26|28207|Masters Degree||Finance: Accountant|28202|0|11|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503959684|503961693|31|0|2|503985328|1|0|2|500775400|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||0|7044657180546140448
M838|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|239|Yellow||2014-09-02|2014-09-17|2015-05-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.9||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28217|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|Black||25|28214|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503535102|503536977|36|0|2|503882165|31|0|2|500774003|5|2|-2||4|2||-2||-2|0|10|||46|2|||1||9134125726462845918|0
M839|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|813|Green|PERL 2014-2016|2014-11-26|2014-12-15|NaT||||26.7||1|1|1|1|M|White||13|No|Mother|28216|6|One Parent: Female|$35,000 to $39,999|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28203|Bachelors Degree|Single|Finance: Banking|28203|7|8|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020753|503989203|503991217|1|0|1|504066226|1|0|1|500799476|10|2|-2||2|1|500014681|-2|500014681|-2|0|5|||17159|12|||1|500014681|3974159976843499574|7314981105541236888
M840|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|965|Red||2012-12-12|2012-12-27|2015-08-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.7||1|1|1|1|F|Black||13|No|Mother|28226|4|One Parent: Female|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||40|28273|Some College|Married|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503268271|503270085|31|0|2|502993922|1|0|2|500669147|5|2|-2||4|3||-2||-2|6854|8|||7496|10|3|3|1||4903779310522421428|7044657180546140448
M841|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1372|Green|Project Big|2012-01-12|2012-01-27|2015-10-30|Volunteer: Moved|Volunteer: Moved||45.1||1|1|1|1|F|Black||13|No|Mother|28206|3|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|F|Black||28|28262|Bachelors Degree|Single|Finance: Banking||0|0|AA Task Force|Special Event|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502868923|502870324|31|0|2|502832013|31|0|2|500591320|10|2|500004641||4|1|500004640|-2||-2|0|4|||11098|8|||1|500004640|7960300212314874874|0
M842|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|24|Green|Cabarrus County|2017-02-02|2017-02-11|NaT||||0.8||1|1|1|1|F|White||13|No|Mother|28025|8|Two Parent|Unknown|||Y|Yes||Therapist/Counselor|General Community|Cabarrus County|Match Support|F|White||31|28025||Separated|Business||0|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504999127|505001687|1|0|2|504999362|1|0|2|500944301|10|2|500016307||2|1|500016374|-2|500016374|-2|0|5|||17159|12|||1|500016374|0|6915279604152465197
M843|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|167|Yellow||2015-07-28|2015-07-28|2016-01-11|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||5.5||1|1|1|1|F|Black||13|No|Mother|28217|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Finance: Banking||2|2|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500018851|504230613|503065429|31|0|2|503995309|1|0|2|500834694|10|2|-2||4|2||-2||-2|0|4|||7464|9|||1||7960300212314874874|2141487034287122220
M844|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|203|Green||2015-09-24|2015-10-13|2016-05-03|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||6.7||1|1|1|1|F|Black||13|No|Mother|28202|6|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Enrollment|F|White||26|28203|Bachelors Degree|Single|Finance|28202|0|5|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333777|504335999|31|0|2|504355120|1|0|2|500842206|5|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|7044657180546140448
M845|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|201|Green|PERL 2014-2016|2014-11-07|2014-11-07|2015-05-27|Child: Changed school/site|Child: Changed school/site||6.6||1|1|4|4|M|Black||13||Mother|28208|6|One Parent: Female|Unknown|||Y|Yes||Self|General Site|PERL 2014-2016|Match Support|M|Black||44|29732|High School Graduate|Married|Business|28217|5|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|501837686|501838054|31|0|1|503754104|31|0|1|500793364|10|1|500009132|2128207319|4|1|500014681|-1||-1|0|10|||11247|3|||1|500014681|3935539763241716148|0
M846|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|280|Green||2016-05-13|2016-05-31|NaT||||9.2||1|1|1|1|M|Black||13|No|Mother|28227|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|Black||27|28205|Some College|Single|Retail: Sales|28210|2|6|Local Radio|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504425160|504427415|31|0|1|504509415|31|0|1|500893007|10|2|-2||2|1||-2||-2|0|4|||7437|1|||1||4112464363801619560|5544164653861671456
M847|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2442|Green||2010-06-14|2010-06-30|NaT||||80.2||2|2|2|2|F|Black||13|No|GrandMother|28269|6|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|501755470|501755813|31|0|2|502038804|31|0|2|500456645|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||6933349951274183958|0
M848|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1117|Green||2013-07-10|2013-07-19|2016-08-09|Volunteer: Moved|Volunteer: Moved||36.7||1|1|1|1|M|Black||13|No|Mother|28213|6|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Enrollment|M|Black||26|28217|Bachelors Degree|Single|Business: Marketing|28217|4|0|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503328946|503330792|31|0|1|503371779|31|0|1|500703253|5|2|-2||4|1||-2||-2|0|10|||7447|3|||1||540227296891876425|514301162572611567
M849|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|120|Green|PERL 2014-2016|2016-10-24|2016-10-31|2017-02-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.9||4|4|1|1|F|Black||13|Yes|Mother|28217|8|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||31|28278|Doctor of Medicine (MD)|Living w/ Significant Other|Medical: Pharmacist||0|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500013781|501319029|500948399|31|0|2|504558901|1|0|2|500918750|5|2|-2||4|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||46|2|||1|500014681|3935539763241716148|0
M850|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1222|Red||2013-01-09|2013-01-31|2016-06-06|Volunteer: Moved|Volunteer: Moved||40.1||4|4|1|1|F|Black||13|Yes|Mother|28217|8|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||28|28212|Bachelors Degree|Married|Child/Day Care Worker||0|3|Local Print|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501319029|500948399|31|0|2|503078205|1|0|2|500673752|5|2|-2||4|3|500014681|-2||-2|0|10|||7439|1|||1||3935539763241716148|0
M851|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|352|Yellow||2014-04-07|2014-04-07|2015-03-25|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||11.6||2|2|1|1|M|Black||13|No|Mother|28027|7|One Parent: Female|Unknown||||Yes||School|General Community|Cabarrus County|RTBM|M|White||50|28025|Associate Degree|Married|Business: Sales|28025|0|7|Current/Previous Big|Other Big|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500012459|503452335|503454201|31|0|1|503845505|1|0|1|500758515|7|1|500000295|2128212924|4|2|500016374|-2||-1|0|4|||17159|12|||1||6750834084344455219|0
M852|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|694|Green||2015-04-13|2015-04-13|NaT||||22.8||1|1|1|1|M|Black||13|No|Mother|28208|6|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||25|28203|Masters Degree|Single|Finance: Accountant|28202|0|3|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504068125|504070152|31|0|1|504241807|1|0|1|500822990|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||932861092942387634|6156547733130613405
M853|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|127|Green||2015-01-15|2015-02-10|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||4.2||1|1|3|3|M|Black||13|No|Mother|28206|6|Two Parent|Unknown|||Y|Yes||School|General Site||Match Support|M|White||29|28202|Bachelors Degree|Single|Business: Engineer|28202|5|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504152757|504154807|31|0|1|503979778|1|0|1|500808239|10|1|500009132|2128173561|4|1||-1|500014681|-1|0|4|||16705|3|||1||7960300212314874874|0
M854|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1442|Green||2013-03-19|2013-03-26|NaT||||47.4||1|1|1|1|M|White||13|No|Mother|28213|6|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||32|28104|Bachelors Degree|Single|Business|20785|0|5|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502866083|502867478|1|0|1|503378884|1|0|1|500688846|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||932861092942387634|0
M855|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1442|Green||2013-03-08|2013-03-26|NaT||||47.4||1|1|1|1|M|White||13|No|Mother|28213|6|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||32|28210|Bachelors Degree|Single|Business: Sales||4|6|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020752|502866079|502867478|1|0|1|503378886|1|0|1|500686789|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||932861092942387634|0
M856|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|143|Green|Cabarrus County|2016-10-05|2016-10-15|NaT||||4.7||1|1|1|1|M|Black||13|No|Mother|28027|7|One Parent: Female|$50,000 to $59,999||||Yes||Self|General Community|Cabarrus County|Match Support|M|White||32|28027|Some College|Married|Business: Sales|28216|5|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504507408|504509703|31|0|1|504651211|1|0|1|500913035|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|500016374|6750834084344455219|4173153455025080196
M857|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|519|Green||2015-09-16|2015-10-05|NaT||||17.1||1|1|1|1|M|Black||13|No|Mother|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|M|Black||27|28262|Bachelors Degree|Single|Finance|28202|0|1|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504401907|504404149|31|0|1|504355133|31|0|1|500840434|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M858|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1725|Green|Amachi|2010-04-29|2010-05-11|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||56.7||2|2|1|1|F|White||13|Yes|GrandMother|28083|6|Grandparents|Unknown||||No||Self|General Community||Enrollment|F|White||40|28027||Single|Customer Service|28027|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|501722052|501227925|1|0|2|502030533|1|0|2|500450450|5|2|-2||4|1||-2||-2|0|10|||7464|9|12|3|1|500000294|675996018716794055|0
M859|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2612|Green||2009-03-26|2009-04-06|2016-05-31|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||85.8||1|1|1|1|M|Black||13||Mother|28227|5|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||54|28262|High School Graduate|Married|Disabled||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501597169|501597489|31|0|1|501563612|31|0|1|500352827|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||2056258660718146620|0
M860|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|296|Green||2015-09-23|2015-10-05|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|1|1|F|Black||13|No|Mother|28208|7|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||32|28269|Bachelors Degree|Married|Business: Mgt, Admin|28202|0|9|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333786|504336008|31|0|2|504359851|1|0|2|500841755|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M861|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|280|Green||2014-04-22|2014-04-29|2015-02-03|Volunteer: Time constraint|Volunteer: Time constraint||9.2||4|4|1|1|F|Black||13|Yes|Mother|28205|7|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||39|28204|Bachelors Degree|Single|Self-Employed, Entrepreneur|28206|6|11|Current/Previous Big|Other Big|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|502763524|502764436|31|0|2|503839682|1|0|2|500760511|10|1|500000295|2128173561|4|1||-2||-1|0|4|||17159|12|||1||7960300212314874874|0
M862|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2016-12-13|2017-01-30|NaT||||1.2||4|4|2|2|F|Black||13|Yes|Mother|28205|7|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||24|28227|Associate Degree|Single|Student: College|28211|1|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|502763524|502764436|31|0|2|504370632|1|0|2|500935268|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||7960300212314874874|0
M863|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|247|Green||2015-11-02|2015-11-24|2016-07-28|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.1||4|4|2|2|F|Black||13|Yes|Mother|28205|7|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||24|28227|Associate Degree|Single|Student: College|28211|1|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500016270|502763524|502764436|31|0|2|504370632|1|0|2|500855054|10|1|500000295|2128173561|4|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||7960300212314874874|0
M864|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|766|Green|PERL 2014-2016|2015-01-21|2015-01-31|NaT||||25.2||1|1|1|1|M|Black||13|No|Mother|28105|6|One Parent: Female|$40,000 to $44,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||28|28105|Bachelors Degree|Single|Business: Human Resources|28204|1|2|Other|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|503413169|503415024|31|0|1|504092153|1|0|1|500809276|10|2|-2||2|1|500014681|-2|500014681|-2|34|2|||7671|13|||1|500014681|2129686509389594346|3714886275549507192
M865|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|897|Green||2012-11-12|2012-11-21|2015-05-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||29.5||1|1|1|1|F|White||13||Mother|28027||Two Parent|Unknown||||No||School|General Site||Match Support|F|White||20|28117|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500002335|503292843|503294667|1|0|2|503233785|1|0|2|500658678|10|1|500000295|2128173571|4|1||-1||-1|0|4|||0|4|||1||1550830965009450729|0
M866|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|132|Green||2016-10-17|2016-10-26|NaT||||4.3||1|1|1|1|F|Hispanic||13|No|Mother|28210|8|Two Parent|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|Hispanic||29|28262|Bachelors Degree|Single|Tech: Computer/Programmer|28208|1|7|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504893713|504896233|3|0|2|504783221|3|0|2|500916377|10|1|500009132|2128212899|2|1|500014681|-1||-1|0|4|||7464|9|||1||7276767778509034039|0
M867|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|169|Green||2014-09-09|2014-09-18|2015-03-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.6||1|1|1|1|M|Black||13|No|Mother|28273|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||54|28226|Masters Degree|Single|Tech: Computer/Programmer|28202|0|3|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|503628199|503630137|31|0|1|503966130|1|0|1|500775002|10|2|-2||4|1|500014681|-2|500000294|-2|0|10|||17159|12|||1||7508998544817094399|1564212873682615975
M868|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|572|Green||2015-08-13|2015-08-13|NaT||||18.8||1|1|1|1|F|Black||13|No|Mother|28214|6|One Parent: Female|$50,000 to $59,999||||Yes||Self|General Community||Match Support|F|White||29|28273|Masters Degree|Married|Finance: Accountant|28210|3|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504328960|504331182|31|0|2|504215323|1|0|2|500836079|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||0|8503368421346667831
M869|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|154|Green||2016-09-22|2016-10-04|NaT||||5.1||1|1|3|3|F|Black||13|No|Mother|28211|8|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||29|28209|Bachelors Degree|Single|Business|28202|6|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504855805|504858307|31|0|2|503605799|1|0|2|500909625|10|1|500009132|2128212899|2|1||-1|500014681|-1|0|4|||16705|3|||1||8568001799025358453|0
M870|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|519|Green||2015-09-22|2015-10-05|NaT||||17.1||1|1|1|1|F|Black||13|No|Mother|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||24|28262|Bachelors Degree|Single|Tech: Support, Writing|28208|0|3|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504401919|504404161|31|0|2|504396776|1|0|2|500841382|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M871|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|284|Green||2015-09-22|2015-10-01|2016-07-11|Volunteer: Time constraint|Volunteer: Time constraint||9.3||2|2|1|1|F|Black||13|No|Mother|28208|8|Two Parent|Less than $10,000||||Yes||School|General Site||Match Support|F|White||27|28034|Bachelors Degree|Married|Business|28208|2|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504416613|504418865|31|0|2|504368299|1|0|2|500841639|10|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M872|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|156|Green||2016-09-22|2016-10-02|NaT||||5.1||2|2|1|1|F|Black||13|No|Mother|28208|8|Two Parent|Less than $10,000||||Yes||School|General Site||Match Support|F|White||23|28209|Bachelors Degree|Single|Finance|28208|1|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504416613|504418865|31|0|2|504776839|1|0|2|500909641|10|1|500009132|2128212899|2|1||-1||-1|0|4|||7464|9|||1||7276767778509034039|0
M873|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|682|Green||2013-04-11|2013-04-16|2015-02-27|Child: Graduated|Child: Graduated||22.4||1|1|1|1|F|Hispanic||13|Yes|Mother|28217|4|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||29|28207|Bachelors Degree|Single|Architect|28210|1|0|TV|Media|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500008321|503462811|503464677|3|0|2|503365326|1|0|2|500692462|10|1|-1||4|1||-1||-1|0|4|||130|1|||1||8568001799025358453|0
M874|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|15|Green||2017-01-24|2017-02-20|NaT||||0.5||1|1|1|1|F|Hispanic||13|No|Mother|28226|7|One Parent: Female|$10,000 to $14,999||||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Hispanic|Mexican|22|28227|Bachelors Degree|Single|Tech: Management|28202|0|4|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504672339|504674766|3|0|2|504870474|3|10|2|500941713|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||384008102559124244|5081726734274569781
M875|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1950|Green||2011-10-14|2011-11-04|NaT||||64.1||1|1|1|1|F|Hispanic||13|No|Mother|28278|3|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|F|White||32|28211||Married|Finance||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500017732|502728289|502729186|3|0|2|502339145|1|0|2|500565493|10|2|-2||3|1||-2|500000294|-2|0|3|||7496|10|||1||3539543368195872575|3151684623133646168
M876|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1973|Green|Amachi, Cabarrus County|2011-10-03|2011-10-12|NaT||||64.8||1|1|1|1|M|White||13|Yes|Mother|28025|5|One Parent: Female|Unknown||||Yes||School|General Community|Cabarrus County|Match Support|M|White||47|28025||Single|Tech: Support, Writing|28026|0|2|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502721278|501938680|1|0|1|502701096|1|0|1|500560499|10|2|500003586||2|1|500016374|-2|500016374|-2|0|4|||7464|9|||1|500000294, 500016374|5173041326630627506|0
M877|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1880|Green||2012-01-03|2012-01-13|NaT||||61.8||1|1|1|1|M|Black||13|No|Mother|28217|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||30|28202|Bachelors Degree|Single|Business: Sales|28212|0|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502700500|502701345|31|0|1|502824634|1|0|1|500589524|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||0|0
M878|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|602|Green||2013-10-07|2013-10-07|2015-06-01|Child: Graduated|Child: Graduated||19.8||2|2|1|1|M|Black||13|No|Mother|28217|2|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||20|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502763379|502764291|31|0|1|503613615|1|0|1|500716288|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M879|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|349|Green||2015-09-22|2015-10-06|2016-09-19|Child: Lost interest|Child: Lost interest||11.5||1|1|3|3|F|Hispanic||13|No|Mother|28210|7|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|F|White||29|28209|Bachelors Degree|Single|Business|28202|6|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504410201|504412452|3|0|2|503605799|1|0|2|500841351|10|1|500009132|2128212899|4|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|7044657180546140448
M880|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1184|Yellow||2011-09-12|2011-10-19|2015-01-15|Volunteer: Moved|Volunteer: Moved||38.9||1|1|2|2|F|Hispanic||13|No|Mother|28269|5|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Enrollment|F|Black||52|30080|Bachelors Degree|Single|Consultant|2451|3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|502551048|502551498|3|0|2|501472128|31|0|2|500554178|5|2|-2||4|2||-2||-2|0|4|||7464|9|||1||4952249713946979108|0
M881|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|368|Red||2014-06-18|2014-06-20|2015-06-23|Volunteer: Time constraint|Volunteer: Time constraint||12.1||3|3|1|1|M|Black||13|No|Mother|28216|6|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||28|28209|Bachelors Degree|Single|Business|28278|2|2|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502912138|502913549|31|0|1|503857059|1|0|1|500767007|5|2|-2||4|3||-2||-2|34|2|||46|2|||1||9134125726462845918|3402014428779854546
M882|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1592|Red||2012-04-05|2012-04-30|2016-09-08|Volunteer: Moved|Volunteer: Moved||52.3||1|1|1|1|M|Black||13|No|Mother|28213|8|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Enrollment|M|White||38|28206|Bachelors Degree|Divorced|Business: Mgt, Admin|28164|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502763968|502764880|31|0|1|502939016|1|0|1|500608284|5|2|-2||4|3||-2||-2|0|10|||7496|10|||1||7284449467126735125|6509979088654253145
M883|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Pending Match|176|Red|PERL 2014-2016|2015-03-26|2015-04-14|2015-10-07|Volunteer: Moved|Volunteer: Moved||5.8||1|2|1|1|F|Multi-race (Hispanic & White)||13|No|Mother|28205|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community||Pending Match|F|White||30|28205|Bachelors Degree|Separated|Business|28205|0|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500013781|504205508|504207619|35|0|2|504157187|1|0|2|500820606|9|2|-2||4|3||-2|500014681|-2|0|5|||17159|12|||1|500014681|8758769076374727509|610388910998118020
M884|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|435|Green||2014-04-10|2014-04-14|2015-06-23|Child: Changed school/site|Child: Changed school/site||14.3||1|1|1|1|M|Black||13|No|Mother|28217|4|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|Black||42|28105|Bachelors Degree|Divorced|Business: Clerical|28210|1|3|BBBS National Site|Web Link|Big|General Site||RTBM|1|0|1|0|277|60|598|500000170|500016847|503870487|503872481|31|0|1|503813685|31|0|1|500759270|10|1|500000295|2128173557|4|1||-1||-1|0|4|||46|2|||1||8981704271528751143|0
M885|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|863|Green|PERL 2014-2016|2014-10-23|2014-10-26|NaT||||28.4||1|1|1|1|M|Black||13|No|Mother|28262|6|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|Multi-race (Asian & White)||36|28203|Masters Degree|Married|Finance: Banking|20815|11|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500018851|503915384|503917391|31|0|1|503995835|37|0|1|500787470|10|2|-2||2|1|500014681|-2|500014681|-2|34|2|||7464|9|||1|500014681|4726905079488957916|8283117761446993531
M886|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|24|Green|Cabarrus County|2017-02-08|2017-02-11|NaT||||0.8||2|2|3|3|M|Multi-race (Black & White)||13|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||||No||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504517520|504519821|36|0|1|501284751|31|0|1|500945238|10|2|-2||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316|-2|0|4|||132|8|||1|500016374|4621676786129919860|0
M887|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|402|Red|PERL 2014-2016, Cabarrus County|2015-11-20|2015-12-07|2017-01-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.2||2|2|1|1|M|Multi-race (Black & White)||13|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||||No||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|Black||26|28262|Bachelors Degree|Single|Business: Sales|28025|0|1|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500022817|504517520|504519821|36|0|1|504355611|31|0|1|500862169|10|2|500016307||4|3|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||17159|12|||1|500014681, 500016374|4621676786129919860|0
M888|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|267|Green||2014-09-04|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|2|2|F|Hispanic||13|No|Mother|28216|3|One Parent: Female|Unknown|||Y|Yes||Self|General Site||Enrollment|F|White||30|28202|High School Graduate|Single|Finance|28202|0|5|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503610365|503612230|3|0|2|503615532|1|0|2|500774531|5|1|500009132|2128173561|4|1||-1||-1|0|10|||16705|3|||1||7960300212314874874|0
M889|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|990|Green||2014-06-12|2014-06-21|NaT||||32.5||1|1|1|1|M|Black||13|No|Mother|28212|6|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28202|Masters Degree|Single|Finance: Banking|28244|0|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503879123|503881119|31|0|1|503889097|1|0|1|500766443|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1||8758769076374727509|5021690776253335384
M890|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1175|Green||2013-12-11|2013-12-18|NaT||||38.6||1|1|1|1|F|Black||13|No|Mother|28214|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||35|28204|Bachelors Degree|Single|Retail: Mgt|28273|1|10|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503688885|503690850|31|0|2|503606993|1|0|2|500738203|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||7089569121628268952|0
M891|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|336|Green||2015-09-22|2015-10-19|2016-09-19|Child: Changed school/site|Child: Changed school/site||11||1|1|1|1|F|Black||13|No|Mother|28215|6|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|F|White||26|28203|Bachelors Degree|Single|Tech: Engineer|28202|2|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504396338|504398578|31|0|2|504353900|1|0|2|500841387|10|1|500009132|2128212899|4|1||-1||-1|0|3|||16705|3|||1||7276767778509034039|0
M892|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|530|Red||2014-08-21|2014-09-17|2016-02-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.4||1|1|1|1|F|Black||13|No|Mother|28214|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||40|28056|Some College|Single|Real Estate: Realtor|28202|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503898651|503891857|31|0|2|503494199|31|0|2|500773073|10|2|-2||4|3||-2||-2|0|10|||46|2|||1||64486389764866818|7044657180546140448
M893|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2205|Green|Amachi|2011-02-09|2011-02-22|NaT||||72.4||1|1|1|1|M|Black||13|Yes|Mother|28134|6|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||29|28273|Some College|Single|Govt: Mgmt/Admin|28208|2|0|Relative|Relative|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020752|501712048|501712386|31|0|1|502405439|1|0|1|500516322|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||17161|11|||1|500000294|7872663507285703533|0
M894|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2297|Green|Amachi, Project Big, Project Big AND Amachi|2010-10-28|2010-11-22|NaT||||75.5||1|1|1|1|F|Black||13|Yes|Mother|28208|4|One Parent: Female|Unknown|||Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||31|29605|Bachelors Degree|Single|Business: Human Resources|29615|1|0|Local TV|Media|Big|General Community|Project Big AND Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|502353937|502354375|31|0|2|501672025|1|0|2|500487322|10|2|500004772||2|1|500000294, 500004640, 500004901|-2|500004901|-2|0|4|||7438|1|||1|500000294, 500004640, 500004901|6458351142431041105|0
M895|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|367|Red||2014-10-01|2014-10-13|2015-10-15|Volunteer: Moved|Volunteer: Moved||12.1||1|1|1|1|M|Black||13|Yes|Mother|28215|6|One Parent: Female|$10,000 to $14,999||||Yes||Self|General Community||Enrollment|M|Black||25|28205|Bachelors Degree|Single|Tech: Research/Design|28202|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503723868|503725860|31|0|1|503940354|31|0|1|500779635|5|2|-2||4|3||-2||-2|0|10|||17159|12|||1||5741767063897867874|8861046674172959830
M896|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|196|Yellow||2014-11-03|2014-12-03|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||6.4||1|1|2|2|F|Black||13|No|Mother|28205|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||28|28203|Bachelors Degree|Single|Tech: Research/Design|28202|0|11|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504100809|504102843|31|0|2|503979771|1|0|2|500791453|10|1|500009132|2128173561|4|2||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M897|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2010|Green||2011-03-08|2011-03-23|2016-09-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||66||1|1|1|1|M|Black||13|No|Mother|28277|5|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||34|28262||Married|Finance|29715|6|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500017732|502249189|502249620|31|0|1|502485458|31|0|1|500523907|10|2|-2||4|1||-2||-2|34|2|||7462|13|||1||0|0
M898|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|793|Yellow||2013-06-05|2013-07-30|2015-10-01|Volunteer: Time constraint|Volunteer: Time constraint||26.1||2|2|2|2|F|White||13|No|Father|28211|8|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||58|28277|High School Graduate|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503405468|503407325|1|0|2|502944301|1|0|2|500699540|10|2|-2||4|2|500014681|-2||-2|0|10|||7464|9|||1||4440360203097874486|5081726734274569781
M899|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|411|Green|PERL 2014-2016|2016-01-04|2016-01-21|NaT||||13.5||2|2|1|1|F|White||13|No|Father|28211|8|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||31|28205|Bachelors Degree|Single|Business: Mgt, Admin|28269|8|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500013781|503405468|503407325|1|0|2|504322859|1|0|2|500870080|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|500014681|4440360203097874486|5081726734274569781
M900|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|284|Green||2015-09-22|2015-10-01|2016-07-11|Volunteer: Time constraint|Volunteer: Time constraint||9.3||1|1|1|1|F|Black||13|No|Mother|28212|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|PERL 2014-2016|Enrollment|F|White||33|28202|Bachelors Degree|Single|Business|28208|0|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504401940|504404182|31|0|2|504368976|1|0|2|500841350|5|1|500009132|2128212899|4|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M901|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|691|Green||2014-07-11|2014-09-10|2016-08-01|Child/Family: Moved|Child/Family: Moved||22.7||1|1|1|1|M|Black||13|No|Mother|28212|7|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Enrollment|M|White||44|28203|Masters Degree|Single|Finance|29715|10|0|Igniting Breakfast|Special Event|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503743876|503261158|31|0|1|503908096|1|0|1|500769242|5|2|-2||4|1||-2||-2|0|10|||17266|8|||1||2811191761055817959|7044657180546140448
M902|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|317|Green|Cabarrus County, mentor2.0 2016|2016-03-28|2016-04-24|NaT||||10.4||1|1|1|1|F|Black||13|No|Mother|28027|7|Two Parent|$60,000 to $74,999||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||30|28269|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|2|Recruitment Event|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504602680|504605091|31|0|2|504579649|1|0|2|500886605|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7462|13|||1|500016374, 500016394|6353565629814722343|993637920138474088
M903|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|155|Green||2016-09-29|2016-10-03|NaT||||5.1||1|1|1|1|M|Black||13|No|GrandMother|28271|8|One Parent: Female|Unknown|||Y|Yes||Self|General Site||Match Support|M|Multi-Race (None of the above)||26|28202|Masters Degree|Married|Tech: Support, Writing|28202|1|1|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504868978|504871497|31|0|1|504855899|7|0|1|500911560|10|1|500009132|2128212899|2|1||-1||-1|0|10|||7464|9|||1||8568001799025358453|0
M904|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|296|Green||2015-09-23|2015-10-05|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|3|3|M|Black||13|Yes|Mother|28208|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||30|28273|Bachelors Degree|Single|Finance|28202|1|8|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504423105|504425358|31|0|1|503911379|1|0|1|500841794|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M905|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|396|Red||2014-09-08|2014-09-29|2015-10-30|Volunteer: Moved|Volunteer: Moved||13||1|1|1|1|M|Black||13|Yes|Mother|28227|5|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||34|28209|Masters Degree|Single|Finance: Accountant|28210|2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|503851354|503853343|31|0|1|503962684|1|0|1|500774775|10|2|-2||4|3||-2|500000294|-2|0|10|||46|2|||1||314687390558932914|7782268353089690742
M906|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|288|Yellow|PERL 2014-2016|2015-05-14|2015-05-31|2016-03-14|Child/Family: Moved|Child/Family: Moved||9.5||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28134|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28273|Bachelors Degree|Single|Architect|28273|0|11|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500008321|504202968|504205079|36|0|1|504285700|1|0|1|500827095|10|2|-2||4|2|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681|3539543368195872575|7165641474360673060
M907|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|111|Green|PERL 2014-2016, Cabarrus County|2016-11-14|2016-11-16|NaT||||3.6||1|1|1|1|M|White||13|No|Foster Parent|28027|6|One Parent: Male|$100,000 to $124,999|||Y|No|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||28|28269|Bachelors Degree|Single|Medical|46250|0|7|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504748250|504750703|1|0|1|504885284|1|0|1|500927298|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||17159|12|||1|500014681, 500016374|0|71389706163855294
M908|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1070|Red||2013-10-14|2013-10-23|2016-09-27|Child: Family structure changed|Child: Family structure changed||35.2||1|1|1|1|M|Black||13|No|Mother|28215|5|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Asian||54|28211|Masters Degree|Married|Self-Employed, Entrepreneur|28211|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503506115|503507986|31|0|1|503552068|4|0|1|500718774|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||0|0
M909|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|372|Green||2014-03-10|2014-03-19|2015-03-26|Child/Family: Moved|Child/Family: Moved||12.2||1|1|1|1|F|Black||13|No|Mother|28134|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||37|28209|Bachelors Degree|Divorced|Medical|28078|5|6|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|502987717|502989174|31|0|2|503559146|1|0|2|500753781|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1||3539543368195872575|6326176198457285184
M910|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|135|Green||2015-09-16|2015-10-07|2016-02-19|Volunteer: Time constraint|Volunteer: Time constraint||4.4||1|1|1|1|M|Black||13|No|Mother|28208|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Enrollment|M|Hispanic||43|28210|Bachelors Degree|Married|Business|28202|2|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504348606|504350830|31|0|1|504368342|3|0|1|500840441|5|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M911|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|736|Green|PERL 2014-2016|2015-02-24|2015-03-02|NaT||||24.2||1|1|1|1|F|Black||13|No|Mother|28216|6|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||33|28205|Bachelors Degree|Single|Tech: Sales, Mktg|28217|7|11|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|504038302|504040320|31|0|2|504099787|1|0|2|500815247|10|2|-2||2|1|500014681|-2|500014681|-2|0|5|||7464|9|||1|500014681|7883015200677941272|0
M912|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|267|Green||2014-09-18|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|1|1|F|Black||13|No|Mother|28205|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||46|29708||Married|Finance: Accountant|28202|5|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504030009|504032027|31|0|2|503910147|1|0|2|500776821|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M913|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|597|Green||2014-02-13|2014-02-25|2015-10-15|Child/Family: Moved|Child/Family: Moved||19.6||1|1|1|1|F|Black||13|No|Mother|28052|5|Two Parent|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||32|28202|Masters Degree|Single|Medical: Doctor, Provider|28204|0|11|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|502939347|502940773|31|0|2|503598887|1|0|2|500748884|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||7508998544817094399|0
M914|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|519|Green||2015-09-22|2015-10-05|NaT||||17.1||1|1|1|1|M|Black||13|No|Mother|28203|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|M|Multi-Race (None of the above)||37|28078|Bachelors Degree|Single|Finance|28202|0|5|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504410173|504412424|31|0|1|504350008|7|0|1|500841395|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|4202495335769973196
M915|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1057|Green||2012-05-08|2012-05-21|2015-04-13|Volunteer: Time constraint|Volunteer: Time constraint||34.7||1|1|1|1|F|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||32|28210|Bachelors Degree|Married|Business: Human Resources|28269|0|5|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|502997224|502998689|31|0|2|502939526|31|0|2|500613729|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1||8758769076374727509|0
M916|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2113|Green||2011-05-05|2011-05-25|NaT||||69.4||1|1|1|1|F|Black||13|No|Mother|28216|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||41|28207|Masters Degree|Married|Business: Marketing|28202|2|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502576641|502577144|31|0|2|502537061|1|0|2|500535114|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||0|0
M917|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1788|Green||2011-09-01|2011-09-09|2016-08-01|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||58.7|Y|1|1|1|1|M|Black||13|Yes|Mother|28212|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||51|28205|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|502471024|502471471|31|0|1|502685747|1|0|1|500552890|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||2811191761055817959|0
M918|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|989|Red||2013-05-10|2013-05-21|2016-02-04|Child/Family: Moved|Child/Family: Moved||32.5||2|2|1|1|F|Black||13|No|Mother|29732|6|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|F|White||31|28226|Bachelors Degree|Single|Medical: Healthcare Worker|28211|0|3|Self|Self|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500013781|502073665|502074089|31|0|2|503245956|1|0|2|500696434|7|2|-2||4|3||-2|500000294|-2|0|10|||7464|9|||1||0|0
M919|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|649|Green|PERL 2014-2016|2015-05-19|2015-05-28|NaT||||21.3||1|1|1|1|M|Multi-race (Black & Hispanic)||13|No|Mother|28208|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||29|28208|Masters Degree|Single|Finance: Accountant|28210|3|6|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503924157|503926164|38|0|1|504277947|1|0|1|500827570|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681|5424205421938369753|7044657180546140448
M920|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|99|Green||2016-11-11|2016-11-28|NaT||||3.3||1|1|1|1|M|White||13|No|Mother|28277|8|One Parent: Female|$60,000 to $74,999||||No||Self|General Community|PERL 2014-2016|Match Support|M|White||26|28207|Masters Degree|Living w/ Significant Other|Tech: Engineer|28203|1|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504808434|504810913|1|0|1|504557160|1|0|1|500926948|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||5994075768656267011|5571803589598086587
M921|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|254|Green|PERL 2014-2016|2015-06-23|2015-06-23|2016-03-03|Child/Family: Moved|Child/Family: Moved||8.3||1|1|1|1|F|Black||13|No|Mother|28134|6|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||30|28277|Bachelors Degree|Single|Business: Clerical|28277|1|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|502205926|502206355|31|0|2|504225335|1|0|2|500831147|10|2|-2||4|1|500014681|-2||-2|0|5|||7464|9|||1|500014681|7872663507285703533|6178126991714892144
M922|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-03|2016-10-20|NaT||||4.5||1|1|3|3|M|Black||13|No|Mother|28269|6|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||30|28202|Bachelors Degree|Single|Finance: Accountant|28202|2|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504875016|504877536|31|0|1|503908898|1|0|1|500911987|10|1|500009132|2128207318|2|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M923|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|354|Green||2015-09-22|2015-10-01|2016-09-19|Child: Changed school/site|Child: Changed school/site||11.6||1|1|2|2|M|Black||13|No|Mother|28203|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|M|White||28|28211|Bachelors Degree|Married|Tech: Computer/Programmer|28202|4|6|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504250982|504253098|31|0|1|504349938|1|0|1|500841347|10|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|7044657180546140448
M924|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-22|2015-10-01|NaT||||17.2||1|1|1|1|F|Black||13|No|Mother|28217|8|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|F|White||49|28117||Married|Law||1|6|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504416684|504418936|31|0|2|504338378|1|0|2|500841380|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M925|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|362|Green|PERL 2014-2016|2016-02-26|2016-03-10|NaT||||11.9||1|1|1|1|M|Black||13|No|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28202|Bachelors Degree|Single|Law|28202|0|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504237243|504239358|31|0|1|504456306|1|0|1|500881682|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|500014681|0|7044657180546140448
M926|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|891|Green||2014-09-18|2014-09-28|NaT||||29.3||1|1|1|1|M|Multi-race (Asian & White)||13|No|Mother|28078|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Married|Unemployed|28031|6|2|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503833936|503835915|37|0|1|502489398|1|0|1|500776719|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||836952159905822963|0
M927|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|819|Green||2014-12-05|2014-12-09|NaT||||26.9||1|1|1|1|F|Black||13|No|Mother|28217|8|One Parent: Female|Unknown|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||28|28105|Masters Degree|Married|Business: Mgt, Admin|28211|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|504139056|504094626|31|0|2|503991266|1|0|2|500801765|10|2|-2||2|1||-2||-2|0|5|||17159|12|||1||8568001799025358453|5021631233330154962
M928|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|775|Yellow||2012-11-07|2012-11-30|2015-01-14|Volunteer: Moved|Volunteer: Moved||25.5||1|1|1|1|F|Black||13|No|Mother|28205|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||34|28202|Associate Degree|Single|Medical: Healthcare Worker||6|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503063881|503065564|31|0|2|503125383|1|0|2|500656877|10|2|-2||4|2||-2||-2|0|10|||46|2|||1||5533634913091743658|7044657180546140448
M929|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|630|Green||2015-05-29|2015-06-16|NaT||||20.7||1|1|1|1|M|Black||13|No|Mother|28216|6|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Business|28217|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504247189|504249305|31|0|1|504228103|1|0|1|500828700|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||2456895876914964961|3402014428779854546
M930|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|642|Green||2013-10-16|2013-10-17|2015-07-21|Volunteer: Moved|Volunteer: Moved||21.1||2|2|1|1|M|Black||13|No|Mother|28215|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503671715|503673676|31|0|1|503576626|1|0|1|500720061|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M931|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|238|Green||2015-10-09|2015-10-15|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.8||2|2|2|2|M|Black||13|No|Mother|28215|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||18|28203|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503671715|503673676|31|0|1|504324165|1|0|1|500846378|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M932|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|296|Green||2015-09-16|2015-10-05|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|3|3|M|Black||13|No|Father|28208|7|Two Parent|$30,000 to $34,999||||Yes||Relative|General Site|PERL 2014-2016|Match Support|M|Black||25|28269|Masters Degree|Single|Finance|28202|0|1|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504423077|504425330|31|0|1|504359606|31|0|1|500840435|10|1|500009132|2128207318|4|1|500014681|-1|500014681|-1|0|3|||12831|3|||1||2611337051335117774|0
M933|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1148|Green||2013-12-02|2014-01-14|NaT||||37.7||1|1|1|1|M|Multi-Race (None of the above)||13|No|Mother|28134|5|Other Relative|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|Hispanic||26|28205|||Student: College||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503594290|503596167|7|0|1|503508074|3|0|1|500735488|10|2|-2||2|1||-2||-2|0|5|||7464|9|||1||3539543368195872575|270895945650648132
M934|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|655|Green||2015-05-22|2015-05-22|NaT||||21.5||1|1|2|2|F|Black||13|No|Mother|28212|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502930499|502931919|31|0|2|502564910|31|0|2|500828045|10|2|-2||2|1||-2||-2|0|10|||17161|11|||1||2811191761055817959|3402014428779854546
M935|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|985|Green||2014-05-06|2014-05-15|2017-01-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||32.4||1|1|1|1|M|White||13|No|Mother|28211|6|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||27|28270|Bachelors Degree|Single|Education: Teacher Asst/Aid|28202|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503770823|503772799|1|0|1|503850589|1|0|1|500762293|10|2|-2||4|1||-2||-2|34|2|||46|2|||1||2762897743412756173|7044657180546140448
M936|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|720|Green||2014-02-25|2014-03-20|2016-03-09|Volunteer: Moved|Volunteer: Moved||23.7||1|1|1|1|F|Black||13|No|Mother|28205|5|One Parent: Female|Unknown|||Y|Yes||Therapist/Counselor|General Community||Enrollment|F|White||33|28210|PHD|Single|Business: Human Resources|28273|0|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503689574|503691539|31|0|2|503577882|1|0|2|500751079|5|2|-2||4|1||-2||-2|0|5|||7464|9|||1||0|7044657180546140448
M937|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|699|Green||2015-03-31|2015-03-31|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||23||1|1|1|1|F|Black||13|No|Mother|28273|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Black||28|28105|Masters Degree|Single|Business: Human Resources|28078|0|5|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|504165911|504167953|31|0|2|504030347|31|0|2|500821362|10|2|-2||4|1||-2||-2|0|4|||46|2|||1||5711791743715234276|5161383151676749743
M938|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|127|Green||2016-02-29|2016-03-23|2016-07-28|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||4.2||1|1|3|3|F|Black||13|No|Mother|28208|5|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|Black||30|28270|Masters Degree|Single|Finance|28202|0|1|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504626085|504628496|31|0|2|504396349|31|0|2|500882057|10|1|500009132|2128207318|4|1||-1||-1|0|4|||16705|3|||1||2611337051335117774|0
M939|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|287|Green||2015-09-23|2015-10-14|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.4||1|1|2|2|F|Black||13|No|Mother|28208|6|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||38|28120|Masters Degree|Divorced|Finance: Accountant|28202|6|4|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333815|504336037|31|0|2|504348456|1|0|2|500841759|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M940|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|47|Green||2015-10-14|2015-10-15|2015-12-01|Child: Changed school/site|Child: Changed school/site||1.5||1|1|3|3|M|Black||13|No|Father|28227|6|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|M|White||24|29708|Bachelors Degree|Single|Finance|28202|0|10|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504431587|504433842|31|0|1|504475369|1|0|1|500847980|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M941|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1813|Green|Amachi|2010-09-13|2010-09-29|2015-09-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||59.6||1|1|1|1|F|Black||13|Yes|Mother|28216|1|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||28|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501859854|501860227|31|0|2|502044100|31|0|2|500469954|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294|1653226628427425023|0
M942|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|321|Green||2016-03-15|2016-04-20|NaT||||10.5||2|2|1|1|M|Black||13|No|GrandMother|28208|6|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|White||45|28205|Bachelors Degree|Married|Business: Mgt, Admin|28244|4|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|503893808|503227914|31|0|1|504546078|1|0|1|500884843|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||8998367770661215127|7044657180546140448
M943|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|312|Red||2014-12-11|2014-12-20|2015-10-28|Volunteer: Moved|Volunteer: Moved||10.3||2|2|1|1|M|Black||13|No|GrandMother|28208|6|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|Asian||27|28203|Bachelors Degree|Single|Finance: Accountant|28202|1|10|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500013745|503893808|503227914|31|0|1|503976460|4|0|1|500803592|10|2|-2||4|3||-2|500014506|-2|0|4|||7462|13|||1||8998367770661215127|7044657180546140448
M944|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1558|Green||2012-11-27|2012-11-30|NaT||||51.2||1|1|1|1|M|Black||13|No|Mother|28269|4|One Parent: Female|$30,000 to $34,999|Yes: Active|No||No||Self|General Community||Match Support|M|Black||32|28217|Masters Degree|Single|Consultant||0|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503163476|503165154|31|0|1|503119713|31|0|1|500663695|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||4356567821563751981|3013910978162986880
M945|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|223|Green||2014-10-04|2014-10-22|2015-06-02|Child: Graduated|Child: Graduated||7.3||4|4|2|2|F|Hispanic||13||Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502335365|502335800|3|0|2|503603503|1|0|2|500780614|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M946|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|179|Red|Cabarrus County|2016-09-02|2016-09-09|NaT||||5.9||1|1|1|1|F|Black||13|No|Mother|28025|7|One Parent: Female|$40,000 to $44,999||||No||Self|General Community|Cabarrus County|Match Support|F|Black||47|28075|Masters Degree|Married|Finance: Banking|28282|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504633835|504636246|31|0|2|504775410|31|0|2|500906055|10|2|500016307||2|3|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7496|10|||1|500016374|0|7410064544211008071
M947|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|358|Green||2016-02-29|2016-03-14|NaT||||11.8||1|1|1|1|F|Black||13|No|Mother|28278|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||39|28134|Bachelors Degree|Single|Business: Marketing|28204|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504161470|504162947|31|0|2|504396335|1|0|2|500882097|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||8567789404096574827|2876415545463317777
M948|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|911|Red||2013-11-18|2013-11-26|2016-05-25|Child: Graduated|Child: Graduated||29.9||1|1|1|1|F|Black||13|No|Mother|28217|4|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||29|28277|Bachelors Degree|Single|Medical|70471|2|0|BBBS National Site|Web Link|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500013781|503718061|503720028|31|0|2|503472779|1|0|2|500731891|10|1|500000295|2128173557|4|3||-1||-1|0|4|||46|2|||1||8981704271528751143|0
M949|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|483|Green||2014-02-03|2014-02-04|2015-06-02|Child: Graduated|Child: Graduated||15.9||4|4|2|2|F|White||13|No|Mother|28211|1|One Parent: Female|Unknown||||No||School|General Site||Match Support|F|White||20|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502375449|502375887|1|0|2|503493703|1|0|2|500746461|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M950|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|637|Yellow||2013-10-14|2013-10-24|2015-07-23|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||20.9||2|2|1|1|F|Some Other Race||13||Mother|28277|2|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||30|29730|Bachelors Degree|Single|Finance: Accountant|28273|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|502969236|502970672|41|0|2|503567563|1|0|2|500718760|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||1078778250813636816|0
M951|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|693|Green||2015-04-13|2015-04-14|NaT||||22.8||1|1|1|1|F|Black||13|No|Mother|28205|5|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|Black||27|28262|Some College|Single|Medical: Healthcare Worker|28210|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504242976|504245092|31|0|2|504198992|31|0|2|500823043|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||314687390558932914|3988279022378749151
M952|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|813|Green|PERL 2014-2016|2014-12-09|2014-12-15|NaT||||26.7||2|2|1|1|M|Black||13|No|Mother|28214|1|One Parent: Female|$50,000 to $59,999||||No|Big|Neighbor/Friend|General Community|PERL 2014-2016|Match Support|M|White||25|28202|Bachelors Degree|Single|Tech: Computer/Programmer|28244|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500013781|502728419|502729316|31|0|1|504011804|1|0|1|500802308|10|2|-2||2|1|500014681|-2|500014681|-2|6854|8|||17159|12|||1|500014681|0|7910650461096015612
M953|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|237|Green||2014-09-25|2014-10-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||7.8||1|1|1|1|F|Black||13|No|Mother|28206|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||31|28273|Bachelors Degree|Single|Tech: Computer/Programmer|28202|3|0|Ally Financial|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|504007349|504009376|31|0|2|503981896|31|0|2|500778209|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M954|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|609|Green||2013-09-30|2013-09-30|2015-06-01|Child: Graduated|Child: Graduated||20||1|1|1|1|F|Black||13|Yes|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28210||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503629812|503646211|31|0|2|503497377|1|0|2|500714475|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M955|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|155|Green||2016-10-03|2016-10-03|NaT||||5.1||1|1|2|2|F|Black||13|No|Mother|28209|7|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||32|28078|Bachelors Degree|Single|Business: Mgt, Admin|28202|1|4|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504450770|504453026|31|0|2|504359867|1|0|2|500911956|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M956|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|462|Red|PERL 2014-2016|2015-06-15|2015-07-17|2016-10-21|Volunteer: Time constraint|Volunteer: Time constraint||15.2||1|1|1|1|F|Black||13|No|Mother|28213|5|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|White||28|28078|Bachelors Degree|Single|Business|28078|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|504218954|504221068|31|0|2|504099424|1|0|2|500830251|10|2|-2||4|3|500014681|-2||-2|0|4|||46|2|||1|500014681|4013586283864837776|6178126991714892144
M957|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|194|Green||2015-05-28|2015-06-18|2015-12-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.4||1|1|1|1|M|Black||13|Yes|Mother|28214|5|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Asian|Indian|49|28203|Bachelors Degree|Married|Tech: Engineer|28204|10|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504217755|504219869|31|0|1|504131744|4|18|1|500828564|10|2|-2||4|1|500000294|-2||-2|34|2|||17159|12|||1||7857548027029642592|7000602719972091240
M958|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2238|Green||2011-01-13|2011-01-20|NaT||||73.5||1|1|1|1|M|Black||13|No|Mother|28269|6|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28031|Bachelors Degree|Single|Business: Engineer|28036|0|8|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|1|0|0|1|277|60|598|500000170|500020910|502097794|502098218|31|0|1|502425119|1|0|1|500510881|10|2|-2||2|1||-2|500000294, 500004640|-2|34|2|||46|2|||1||2798582775385400033|0
M959|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1540|Green||2012-11-12|2012-12-18|NaT||||50.6||2|2|1|1|M|Multi-race (Hispanic & White)||13|No|Mother|28211||One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||28|28210|Bachelors Degree|Single|Business: Marketing|28224|1|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502184849|502185278|35|0|1|503145815|1|0|1|500658541|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||932861092942387634|0
M960|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|629|Red||2013-08-05|2013-08-22|2015-05-13|Volunteer: Time constraint|Volunteer: Time constraint||20.7||3|3|1|1|F|Black||13|Yes|Mother|28208|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||36|28210|Masters Degree|Divorced|Medical|28209|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503071350|503073009|31|0|2|503421602|1|0|2|500705806|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1||932861092942387634|1332839031590943646
M961|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|348|Green||2016-03-15|2016-03-24|NaT||||11.4||3|3|2|2|F|Black||13|Yes|Mother|28208|6|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||35|28206|Bachelors Degree|Single|Business: Marketing|28208|4|2|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|503071350|503073009|31|0|2|500831828|31|0|2|500884742|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||932861092942387634|1332839031590943646
M962|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|225|Green||2014-10-04|2014-10-22|2015-06-04|Child: Graduated|Child: Graduated||7.4||2|2|2|2|M|Black||13|No|Mother|28211|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|White||19|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503281941|503283760|31|0|1|503907559|1|0|1|500780596|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M963|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|164|Green||2016-01-05|2016-02-08|2016-07-21|Volunteer: Time constraint|Volunteer: Time constraint||5.4||1|1|1|1|F|Black||13|No|Mother|28206|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|F|Asian||32|28216|Bachelors Degree|Married|Tech: Management|28244|0|11|Community Engagement|Special Event|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500016270|504517593|504519894|31|0|2|504526149|4|0|2|500870298|10|1|500000295|2128173561|4|1||-1|500007920, 500011315, 500011316|-1|0|4|||18809|8|||1||7960300212314874874|0
M964|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|266|Green|PERL 2014-2016|2014-09-12|2014-09-24|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||1|1|2|2|M|Black||13|No|Mother|28206|5|One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|White||32|28262|Masters Degree|Married|Business: Mgt, Admin|28202|6|0|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503996783|503998751|31|0|1|503911472|1|0|1|500775711|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1|500014681|7960300212314874874|0
M965|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|319|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-04-13|2016-04-22|NaT||||10.5||1|1|2|2|M|Black||13|No|Mother|28269|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|M|White||42|28214|Bachelors Degree|Divorced|Business: Engineer||10|0|Self|Self|Big|General Community|Amachi, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504554067|504556401|31|0|1|503373934|1|0|1|500888917|10|2|-2||3|1||-2|500000294, 500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|500007920, 500011315, 500011316|384008102559124244|1962015587749138391
M966|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|294|Green||2015-09-23|2015-10-07|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|2|2|M|Hispanic||13|No|Mother|28208|6|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|M|White||25|28210|Bachelors Degree|Single|Finance|28210|0|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333747|504335969|3|0|1|504359691|1|0|1|500841771|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M967|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|505|Green||2015-09-22|2015-10-19|NaT||||16.6||3|3|1|1|F|Black||13|No|Mother|28216|7|One Parent: Female|Less than $10,000||||Yes||School|General Site|PERL 2014-2016|Match Support|F|Black||37|28081|Bachelors Degree|Married|Business|28208|0|8|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|501951335|501951733|31|0|2|504368723|31|0|2|500841343|10|1|500009132|2128212899|2|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|7044657180546140448
M968|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2233|Green||2011-01-20|2011-01-25|NaT||||73.4||1|1|1|1|F|Black||13|No|Mother|28214|1|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|F|White||35|28209|Bachelors Degree|Single|Retail: Sales||6|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502261100|502261532|31|0|2|502284382|1|0|2|500512216|10|2|-2||2|1||-2||-2|0|3|||7464|9|||1||1653226628427425023|3151684623133646168
M969|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|294|Green||2015-09-25|2015-10-07|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|2|3|F|Black||13|No|Mother|28208|6|Two Parent|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|F|Black||27|28213|Bachelors Degree|Single|Finance|28202|0|5|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504416740|504418992|31|0|2|503355514|31|0|2|500842439|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M970|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|621|Green||2015-06-11|2015-06-25|NaT||||20.4||3|3|1|1|F|Black||13|No|GrandMother|28227|5|Grandparents|Unknown||||No||Self|General Community||Match Support|F|Black||31|28210|Associate Degree|Single|Finance|28255|0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502252822|502253254|31|0|2|504229640|31|0|2|500829933|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1||6407809237813394802|0
M971|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|682|Green||2013-11-12|2013-11-19|2015-10-02|Child: Graduated|Child: Graduated||22.4||1|1|3|3|M|Black||13|No|Mother|28083||One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||37|28273||Married|Business||0|0|ACN|Workplace Partner|Big|General Site|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500012459|503692165|503694130|31|0|1|503216970|31|0|1|500730232|10|1|500000295|2128212919|4|1||-1|500016374|-1|0|4|||13581|3|||1||2437132833506538679|0
M972|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1860|Green|Cabarrus County|2012-02-01|2012-02-02|NaT||||61.1||1|1|1|1|F|Black||13|No|Mother|28083||One Parent: Female|Unknown||||Yes||Self|General Community|Cabarrus County|Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502083438|502083853|31|0|2|502657267|31|0|2|500595491|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7496|10|||1|500016374|0|0
M973|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1268|Green|Amachi|2012-04-05|2012-04-30|2015-10-20|Child/Family: Moved|Child/Family: Moved||41.7||2|2|1|1|M|Black||13|Yes|Mother|28210||One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||55|28105|Masters Degree|Married|Law: Lawyer||25|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|501853851|501854219|31|0|1|502922901|1|0|1|500608304|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294|0|0
M974|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|515|Green|PERL 2014-2016, Cabarrus County|2015-09-23|2015-10-09|NaT||||16.9||2|3|3|3|F|American Indian or Alaska Native||13|No|Aunt|28027|3|Other Relative|Unknown||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||50|28075|Bachelors Degree|Married|Education: Admin|28083|0|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|503012569|504347632|6|0|2|502949193|1|0|2|500841835|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|4|||7671|13|||1|500014681, 500016374|2437132833506538679|1791051703918408849
M975|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|571|Green|VOL - Mentoring Hispanic Youth|2014-04-06|2014-04-11|2015-11-03|Child: Graduated|Child: Graduated||18.8||1|1|1|1|M|Hispanic||13|No|Mother|28217|4|One Parent: Female|Unknown|||Y|Yes||School|General Site|VOL - Mentoring Hispanic Youth|Match Support|M|Some Other Race||67|28202||Divorced|Retired||0|0|TV|Media|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020753|503756602|503758574|3|0|1|503825615|41|0|1|500758454|10|1|500000295|2128173557|4|1|500011312|-1||-1|0|4|||130|1|||1|500011312|8981704271528751143|0
M976|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|508|Green||2015-04-07|2015-04-27|2016-09-16|Volunteer: Time constraint|Volunteer: Time constraint||16.7||1|1|1|1|F|Black||13|Yes|Mother|28208|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||33|28202|Bachelors Degree|Divorced|Business|28117|4|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|504075185|504048929|31|0|2|504169746|1|0|2|500822245|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1||7777315526213898088|7044657180546140448
M977|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|222|Green||2014-10-04|2014-10-22|2015-06-01|Child: Graduated|Child: Graduated||7.3||3|3|2|2|M|Black||13|No|Mother|28211|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||20|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502335325|502335760|31|0|1|503500437|1|0|1|500780610|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M978|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|519|Green||2015-09-21|2015-10-05|NaT||||17.1||1|1|1|1|F|Hispanic||13|No|Mother|28210|7|One Parent: Female|Unknown||||Yes||Relative|General Site||Match Support|F|White||24|28269|Bachelors Degree|Married|Tech: Computer/Programmer|28208|0|3|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504416703|504418955|3|0|2|504401855|1|0|2|500841076|10|1|500009132|2128212899|2|1||-1||-1|0|3|||16705|3|||1||7276767778509034039|0
M979|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|202|Green|PERL 2014-2016, Cabarrus County|2016-08-16|2016-08-17|NaT||||6.6||1|1|1|1|M|Black||13|Yes|Mother|28025|6|One Parent: Female|$40,000 to $44,999||||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||53|28027|Bachelors Degree|Married|Finance: Banking||11|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|502392338|502392776|31|0|1|504744814|1|0|1|500903717|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7464|9|||1|500014681, 500016374|5629236573169735714|2806833304218536184
M980|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|519|Green||2015-09-16|2015-10-05|NaT||||17.1||1|1|1|1|F|Black||13|Yes|Mother|28203|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||27|28262|Bachelors Degree|Single|Consultant||0|4|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504410188|504412439|31|0|2|504335835|1|0|2|500840433|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M981|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|223|Green||2014-10-17|2014-10-22|2015-06-02|Child: Graduated|Child: Graduated||7.3||3|3|2|2|F|Black||13|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||20|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502385620|502386058|31|0|2|503633995|1|0|2|500784782|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||0|0
M982|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|588|Green||2013-10-15|2013-10-22|2015-06-02|Child: Graduated|Child: Graduated||19.3||2|2|1|1|F|Black||13|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28210|Some High School|Single|Student: High School|28226|0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502335383|502335818|31|0|2|503493859|1|0|2|500719615|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M983|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-22|2015-10-01|NaT||||17.2||1|1|2|2|M|Black||13|No|Mother|28208|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Site||Match Support|M|White||34|28202|Masters Degree|Single|Business: Engineer|28202|4|5|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|502262109|504229491|31|0|1|503605726|1|0|1|500841373|10|1|500009132|2128212899|2|1||-1||-1|0|10|||16705|3|||1||7276767778509034039|2692660633362571702
M984|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|294|Green||2015-09-23|2015-10-07|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|2|2|M|Black||13|No|Mother|28208|6|Two Parent|$20,000 to $24,999|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|White||50|28134||Single|Tech: Research/Design|28202|0|0|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504348774|504335952|31|0|1|503911351|1|0|1|500841769|10|1|500009132|2128207318|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1||2611337051335117774|8178900818136675730
M985|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1728|Green||2012-05-17|2012-06-13|NaT||||56.8||1|1|1|1|F|Black||13|No|Mother|28206|6|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||27|28208|Bachelors Degree|Single|Business: Mgt, Admin|28213|1|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|502882034|501390617|31|0|2|502983700|31|0|2|500615277|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1||4863631750424600365|5161383151676749743
M986|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1028|Green||2014-04-30|2014-05-14|NaT||||33.8||1|1|1|1|M|Black||13|No|Mother|28213|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|Black||27|28216|Some College|Single|Retail: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503584428|503586305|31|0|1|503839843|31|0|1|500761714|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||4863631750424600365|0
M987|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|569|Green||2014-03-10|2014-03-12|2015-10-02|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||18.7||2|2|1|1|F|Multi-race (Black & White)||13|No|Mother|28083||Two Parent|Unknown||||No||Self|General Site||Match Support|F|White||20|28027|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500002335|502786012|502787193|36|0|2|503553020|1|0|2|500753731|10|1|500000296|2128173571|4|1||-1||-1|0|10|||0|4|||1||5208542183136337346|0
M988|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|1149|Green||2013-04-09|2013-04-15|2016-06-07|Child: Changed school/site|Child: Changed school/site||37.7||1|1|1|1|M|Hispanic||13||Mother|28031|5|One Parent: Female|Unknown||||No||School|General Site||Match Support|M|Hispanic||23|28035|Some College|Single|Student: College||0|0|Kappa Alpha Psi|Fraternity/Sorority|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|502813481|502814758|3|0|1|503009633|3|0|1|500691991|10|1|500000295|2128173570|4|1||-1||-1|0|4|||8693|14|||1||8034889377453131101|0
M989|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|267|Yellow||2014-09-15|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|1|1|M|Black||13|Yes|Father|28206|5|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|Asian||47|28105|Masters Degree|Married|Tech: Management|28202|3|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504025425|504027443|31|0|1|503948833|4|0|1|500776018|10|1|500009132|2128173561|4|2||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M990|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|333|Green|PERL 2014-2016|2015-03-26|2015-03-26|2016-02-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.9||1|1|1|1|M|Black||13|No|Mother|28215|5|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||26|28204|Bachelors Degree|Single|Consultant|28244|1|6|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500018851|502722096|502722991|31|0|1|504213418|1|0|1|500820735|10|2|-2||4|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681|5741767063897867874|8136849793711030748
M991|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|227|Red|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2015-02-20|2015-02-28|2015-10-13|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||7.5||3|3|1|1|M|Hispanic||13|No|Mother|28206|6|One Parent: Female|Unknown||||Yes|Spanish Radio|Media|General Community|PERL 2014-2016|Match Support|M|Hispanic||35|28205|Some College|Single|Business: Mgt, Admin||7|7|Current/Previous Big|Other Big|Big|General Community|VOL - Mentoring Hispanic Youth|Enrollment|0|1|1|0|277|60|598|500000170|500017777|503575828|503577713|3|0|1|504188100|3|0|1|500814809|10|2|-2||4|3|500014681|-2|500011312|-2|7068|1|||17159|12|||1|500011312, 500014681|932861092942387634|0
M992|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|151|Green||2016-09-21|2016-10-07|NaT||||5||3|3|1|1|M|Hispanic||13|No|Mother|28206|6|One Parent: Female|Unknown||||Yes|Spanish Radio|Media|General Community|PERL 2014-2016|Match Support|M|Multi-Race (None of the above)||30|28202|Bachelors Degree|Single|Business|28025|1|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|503575828|503577713|3|0|1|504686759|7|0|1|500909330|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|7068|1|||7464|9|||1||932861092942387634|0
M993|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|239|Green||2014-10-04|2014-10-06|2015-06-02|Child: Graduated|Child: Graduated||7.9||2|2|2|2|F|Hispanic||13|No|Mother|28227|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||23|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503241922|503243719|3|0|2|503507368|1|0|2|500780587|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M994|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|293|Green||2015-09-28|2015-10-08|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.6||1|1|1|1|F|Black||13|No|Mother|28208|6|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|Black||25|28273|Bachelors Degree|Single|Finance|28202|0|1|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504416720|504418972|31|0|2|504438102|31|0|2|500842591|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M995|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|266|Green||2014-09-18|2014-09-23|2015-06-16|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||1|1|1|1|M|Black||13|No|Mother|28205|4|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|White||37|28105|Bachelors Degree|Married|Finance|28202|3|2|Ally Financial|Workplace Partner|Big|General Site||RTBM|1|0|1|0|277|60|598|500000170|500016270|504030013|504032031|31|0|1|503910089|1|0|1|500776838|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M996|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|91|Green||2014-10-04|2014-10-22|2015-01-21|Child/Family: Moved|Child/Family: Moved||3||3|3|3|3|F|Black||13|No|Mother|28211|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502416642|502417080|31|0|2|503500482|1|0|2|500780615|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M997|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|357|Red||2014-05-06|2014-05-22|2015-05-14|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||11.7||2|2|1|1|M|Black||13|Yes|Mother|28204||One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Insurance|28277|5|3|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503663975|503665933|31|0|1|503854225|31|0|1|500762272|10|2|-2||4|3|500000294|-2||-2|0|10|||17159|12|||1||4440360203097874486|0
M998|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|435|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2015-12-17|2015-12-28|NaT||||14.3||2|2|1|1|M|Black||13|Yes|Mother|28204||One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||24|28202|Bachelors Degree|Single|Finance: Banking|28202|0|5|Other|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|503663975|503665933|31|0|1|504468271|1|0|1|500868596|10|2|-2||2|1|500000294|-2|500007920, 500011315, 500011316|-2|0|10|||18267|3|||1|500007920, 500011315, 500011316|4440360203097874486|0
M999|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1284|Green||2011-08-01|2011-08-16|2015-02-20|Child/Family: Moved|Child/Family: Moved||42.2||1|1|1|1|F|Black||13|No|Mother|28212|2|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|F|Black||42|28210|Masters Degree|Single|Business: Clerical|28036|3|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|502634923|502635617|31|0|2|501197016|31|0|2|500548227|10|2|-2||4|1||-2||-2|0|3|||46|2|||1||3038247238543299436|0
M1000|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|111|Red|PERL 2014-2016|2015-08-06|2015-08-11|2015-11-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.6||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28212|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community|PERL 2014-2016|Enrollment|F|White||47|28270|Some College|Married|Homemaker|29020|18|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|504280484|504282684|36|0|2|504226821|1|0|2|500835375|5|2|-2||4|3|500014681|-2||-2|0|3|||7464|9|||1|500014681|2811191761055817959|4694273237201497095
M1001|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|12|Green||2017-02-08|2017-02-23|NaT||||0.4||1|1|1|1|M|Black||13|Yes|GrandMother|28214|7|Grandparents|$75,000 to $99,999|||Y|Yes||Self|General Community||Match Support|M|White||31|28078|Bachelors Degree|Single|Business: Sales|28202|4|9|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504910266|504912793|31|0|1|504829494|1|0|1|500945213|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1||806697982905023857|5163136606149365864
M1002|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|817|Green|PERL 2014-2016, Cabarrus County|2014-12-05|2014-12-11|NaT||||26.8||1|1|1|1|M|Black||13|No|Mother|28025|7|One Parent: Female|$75,000 to $99,999||||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|Black||35|28027|Bachelors Degree|Married|Finance|28217|1|9|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500022817|503666549|503668509|31|0|1|504106972|31|0|1|500801599|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||46|2|||1|500014681, 500016374|1834158761762606452|0
M1003|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|817|Green|PERL 2014-2016, Cabarrus County|2014-12-05|2014-12-11|NaT||||26.8||2|2|2|2|F|Black||13|Yes|Mother|28025|7|One Parent: Female|$75,000 to $99,999||||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||29|28027|Associate Degree|Single|Education||5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500022817|503666553|503668509|31|0|2|500991324|1|0|2|500801722|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||2238|7|||1|500014681, 500016374|1834158761762606452|0
M1004|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-03|2016-10-20|NaT||||4.5||1|1|1|1|M|Black||13|No|Aunt|28208|6|Two Parent|$15,000 to $19,999|||Y|Yes||School|General Site||Match Support|M|White||23|28207|Bachelors Degree|Single|Finance|28202|1|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504869056|504871576|31|0|1|504788305|1|0|1|500911985|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1005|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1131|Green||2014-01-23|2014-01-31|NaT||||37.2||1|1|1|1|M|Black||13|No|Mother|28226|5|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|Black||39|28210|Some College|Single|Arts, Entertainment, Sports|28202|7|2|Recruitment Event|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503034769|503036365|31|0|1|503650997|31|0|1|500744436|10|2|-2||2|1||-2||-2|0|10|||7458|9|||1||6095563712459522926|4319555889117084469
M1006|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|214|Green|PERL 2014-2016|2014-12-01|2015-01-09|2015-08-11|Child/Family: Moved|Child/Family: Moved||7||1|1|1|1|F|Black||13|Yes|Mother|28206|5|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Enrollment|F|Black||24|28216|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Site|PERL 2014-2016|RTBM|0|1|1|0|277|60|598|500000170|500016270|504100841|504102875|31|0|2|503964951|31|0|2|500799926|5|1|500000295|2128173561|4|1|500014681|-1|500014681|-1|0|4|||46|2|||1|500014681|7960300212314874874|0
M1007|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|238|Green||2014-09-15|2014-10-22|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||7.8||1|1|1|1|F|Asian||13|No|Father|28206|5|Two Parent|Unknown||||Yes||School|General Community||Enrollment|F|Black||26|28273|Bachelors Degree|Single|Finance|28202|0|9|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504016980|504018995|4|0|2|503931457|31|0|2|500775987|5|1|500009132|2128173561|4|1||-2||-1|0|4|||12831|3|||1||7960300212314874874|0
M1008|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|596|Red||2013-06-10|2013-06-24|2015-02-10|Volunteer: Time constraint|Volunteer: Time constraint||19.6||2|2|1|1|M|White||13||GrandMother|28210|4|One Parent: Female|Unknown|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||35|28217||Married|Finance||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503469072|503470938|1|0|1|503478672|1|0|1|500700143|10|2|-2||4|3|500014681|-2||-2|0|10|||7464|9|||1||6898335769881586649|7044657180546140448
M1009|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|658|Green|PERL 2014-2016|2015-05-08|2015-05-19|NaT||||21.6||2|2|1|1|M|White||13||GrandMother|28210|4|One Parent: Female|Unknown|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||29|28217|Some College|Single|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|503469072|503470938|1|0|1|504202910|1|0|1|500826264|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||46|2|||1|500014681|6898335769881586649|7044657180546140448
M1010|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|538|Green|PERL 2014-2016|2015-09-10|2015-09-16|NaT||||17.7||1|1|1|1|M|Some Other Race||13|No|Mother|28217|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||38|28205|Masters Degree|Married|Human Services: Social Worker|28204|5|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504155180|501093096|41|0|1|502462446|1|0|1|500839295|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||7464|9|||1|500014681|8981704271528751143|358434295995756137
M1011|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|211|Green||2015-09-24|2015-10-05|2016-05-03|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||6.9||1|1|1|1|F|Some Other Race||13|No|Father|28208|6|Two Parent|Less than $10,000||||Yes||School|General Site||Enrollment|F|White||29|28208|Bachelors Degree|Single|Finance: Auditor|28202|0|3|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504431606|504433861|41|0|2|504355024|1|0|2|500842209|5|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1012|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1657|Green||2012-06-15|2012-07-12|2017-01-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||54.4||1|1|1|1|M|Black||13|No|Mother|28262|5|One Parent: Female|$50,000 to $59,999||||Yes||School|General Community||Match Support|M|Black||34|28269|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|502637766|502638462|31|0|1|503016558|31|0|1|500619500|10|2|-2||4|1||-2||-2|0|4|||7462|13|||1||7102230088759381237|4588361775303425846
M1013|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|217|Green||2014-10-04|2014-10-29|2015-06-03|Child: Graduated|Child: Graduated||7.1||3|3|2|2|M|Multi-race (Black & White)||13|No|Mother|28211|1|One Parent: Female|Unknown||||No||School|General Site||Match Support|M|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502375441|502375879|36|0|1|503507295|1|0|1|500780595|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1014|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|981|Green||2014-06-12|2014-06-30|NaT||||32.2||1|1|1|1|M|Black||13|No|Mother|28215|3|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|M|Black||30|28215|Some College|Single|Transport: Driver|28269|2|4|Local Radio|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|502582366|502582874|31|0|1|503858870|31|0|1|500766366|10|2|-2||2|1||-2||-2|0|10|||7437|1|||1||5741767063897867874|386356889061704511
M1015|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|992|Green||2014-06-13|2014-06-19|NaT||||32.6||1|1|1|1|M|Black||13|No|Mother|28202|4|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Finance: Accountant|28226|0|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503710095|503712061|31|0|1|503872736|1|0|1|500766579|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1||6368218764956286027|5056473444237941296
M1016|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|522|Red||2013-12-17|2014-01-13|2015-06-19|Volunteer: Time constraint|Volunteer: Time constraint||17.1||1|1|1|1|M|Black||13|No|Mother|28034|5|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||25|28217|Bachelors Degree|Single|Tech: Engineer|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|503496815|503773736|31|0|1|503673962|31|0|1|500739342|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1||0|0
M1017|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|46|Green||2017-01-10|2017-01-20|NaT||||1.5||2|3|1|1|M|Black||13|No|Mother|28031|6|Other/Unknown|Unknown||||Yes||School|General Community||Match Support|M|White||27|28031|Masters Degree|Married|Business: Sales|28210|2|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|503250358|503252163|31|0|1|504861106|1|0|1|500939332|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||3974159976843499574|0
M1018|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|189|Green||2016-08-22|2016-08-30|NaT||||6.2||1|1|1|1|F|Multi-race (Black & White)||13|No|Foster Parent|28214|6|Two Parent|$60,000 to $74,999||||No||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||34|28209|Doctor of Medicine (MD)||Medical|28202|0|4|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504338170|504340392|36|0|2|504465810|31|0|2|500904260|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|5|||17159|12|||1||0|2806833304218536184
M1019|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1422|Red||2011-10-17|2011-11-17|2015-10-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||46.7||1|1|1|1|F|Multi-Race (None of the above)||13|No|Mother|28229|2|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Enrollment|F|Black||34|28226|Bachelors Degree|Single|Business: Clerical|28208|0|6|Self|Self|Big|General Community|Project Big|Enrollment|1|0|1|0|277|60|598|500000170|500017777|502747706|502748616|7|0|2|502618438|31|0|2|500566066|5|2|-2||4|3||-2|500004640|-2|0|10|||7464|9|||1||7807202941877299922|6908726775633097392
M1020|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|348|Green||2016-03-14|2016-03-24|NaT||||11.4||1|1|1|1|F|Black||13|No|Mother|28213|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||38|28205|Bachelors Degree|Divorced|Business|28209|6|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504399552|504401793|31|0|2|504544485|1|0|2|500884475|10|2|-2||3|1||-2|500007920, 500011315, 500011316|-2|0|5|||7464|9|||1||6065435025527210335|458259588635328527
M1021|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|154|Green||2016-09-22|2016-10-04|NaT||||5.1||1|1|3|3|F|Black||13|Yes|Mother|28203|7|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||36|28209|Masters Degree|Married|Business: Marketing|28202|0|4|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504853140|504855642|31|0|2|503605824|1|0|2|500909630|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||8568001799025358453|0
M1022|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|377|Green||2014-09-12|2014-09-23|2015-10-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.4||2|3|1|1|M|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||42|28078||Married|Tech: Management||0|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503610226|503612103|31|0|1|503935226|1|0|1|500775736|10|1|500009132|2128173561|4|1||-2||-1|0|4|||12831|3|||1||7960300212314874874|0
M1023|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|407|Green|PERL 2014-2016|2014-09-12|2014-09-29|2015-11-10|Child: Changed school/site|Child: Changed school/site||13.4||1|1|1|1|M|Black||13|Yes|Mother|28206|6|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|M|White||32|28210|Bachelors Degree|Married|Finance: Banking|28202|4|5|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Enrollment|1|0|1|0|277|60|598|500000170|500016270|504013021|504015036|31|0|1|503910269|1|0|1|500775707|10|1|500000295|2128173561|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1|500014681|7960300212314874874|0
M1024|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|115|Green|Cabarrus County|2016-10-17|2016-11-12|NaT||||3.8||1|1|1|1|F|Black||13|No|Mother|28025|7|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community|Cabarrus County|Match Support|F|White||41|28027|Masters Degree|Married|Homemaker||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504792692|504795152|31|0|2|504760167|1|0|2|500916273|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|500016374|6750834084344455219|3918615128866826495
M1025|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|296|Green||2015-09-23|2015-10-05|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|1|1|F|Black||13|Yes|Mother|28208|6|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||28|28226|Bachelors Degree|Married|Business: Mgt, Admin|28202|1|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504416788|504419040|31|0|2|504353866|1|0|2|500841757|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|3337539259677656630
M1026|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1625|Yellow||2012-02-24|2012-03-21|2016-09-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||53.4||1|1|1|1|F|Black||13|No|Mother|28206|2|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||40|28216|Masters Degree|Single|Finance||6|0|Charlotte Cares|Service Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502873189|502874592|31|0|2|502882530|31|0|2|500600322|10|2|-2||4|2||-2||-2|0|4|||11246|6|||1||4208486535559819469|0
M1027|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|790|Green||2014-04-01|2014-04-09|2016-06-07|Child: Changed school/site|Child: Changed school/site||26||1|1|1|1|F|Black||12|No|Father|28031|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||43|28031|Bachelors Degree|Single|Real Estate: Realtor|28031|4|0|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017786|503720575|503722547|31|0|2|503714604|1|0|2|500757766|10|1|500009132|2128207319|4|1||-1||-1|0|4|||7464|9|||1||8034889377453131101|0
M1028|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|58|Green||2017-01-08|2017-01-08|NaT||||1.9||1|1|3|3|M|Black||12|No|Father|28208|7|Two Parent: Not Married|Unknown||||Yes||School|General Site||Match Support|M|White||30|29707|Bachelors Degree|Married|Business: Engineer|28202|6|2|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504976117|504978668|31|0|1|503605644|1|0|1|500938918|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M1029|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1323|Green||2013-07-15|2013-07-23|NaT||||43.5||2|2|1|1|F|Black||12|No|Mother|28216|1|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||38|28273|Bachelors Degree|Separated|Customer Service|28134|1|2|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502207223|502207652|31|0|2|503251424|1|0|2|500703587|10|2|-2||2|1||-2||-2|6854|8|||7464|9|||1||7869308672550505300|0
M1030|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|607|Green||2013-10-04|2013-10-04|2015-06-03|Child: Graduated|Child: Graduated||19.9||3|3|1|1|F|Hispanic||12|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502355228|502355666|3|0|2|503507223|1|0|2|500716170|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1031|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|366|Green||2015-02-02|2015-02-23|2016-02-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12||2|2|1|1|F|White||12|No|Mother|28212||Two Parent|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Enrollment|F|White||27|28209|Bachelors Degree|Single|Business: Sales|28262|0|10|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|503869451|503871445|1|0|2|504135282|1|0|2|500811559|5|2|-2||4|1||-2||-2|0|5|||46|2|||1||540227296891876425|0
M1032|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1132|Green||2014-01-27|2014-01-30|NaT||||37.2||1|1|1|1|F|Black||12|No|Mother|28216|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||29|28210|Bachelors Degree|Single|Business: Marketing|28277|1|5|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503552498|503554371|31|0|2|503538554|1|0|2|500744965|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1||4863631750424600365|1698789781793629886
M1033|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|156|Green||2016-09-22|2016-10-02|NaT||||5.1||1|1|1|1|F|Black||12|No|Mother|28217|7|Two Parent|$15,000 to $19,999||||Yes||School|General Site||Match Support|F|White||22|28204|Bachelors Degree|Single|Business|28208|0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504855744|504858246|31|0|2|504783146|1|0|2|500909640|10|1|500009132|2128212899|2|1||-1||-1|0|4|||7464|9|||1||8568001799025358453|0
M1034|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1019|Green||2014-05-12|2014-05-23|NaT||||33.5||1|1|1|1|F|Multi-race (Black & Hispanic)||12|No|Mother|28215|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||60|28211|Bachelors Degree|Divorced|Tech: Management|28202|2|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503774057|503776034|38|0|2|503665969|1|0|2|500762915|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||4575902950186762737|0
M1035|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|474|Yellow||2014-03-10|2014-03-21|2015-07-08|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||15.6||2|2|2|2|M|White||12|No|Mother|28025|4|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||58|28075|Masters Degree|Married|Business|32824|0|6|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500012459|503532014|503533889|1|0|1|503694720|1|0|1|500753716|10|2|-2||4|2|500000294, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7464|9|||1||4085045877112350207|1786514887916898235
M1036|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|475|Green|Cabarrus County|2015-10-28|2015-11-18|NaT||||15.6||2|2|1|1|M|White||12|No|Mother|28025|4|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||56|28269|Doctor of Medicine (MD)|Married|Medical: Doctor, Provider|28025|28|0|Agency Sponsored|Special Event|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|503532014|503533889|1|0|1|504408440|1|0|1|500853427|10|2|500016307||2|1|500000294, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||16426|8|||1|500016374|4085045877112350207|1786514887916898235
M1037|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|127|Green||2016-03-02|2016-03-23|2016-07-28|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||4.2||1|1|2|2|F|Black||12|Yes|Mother|28205|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|F|White||35|28226|Bachelors Degree|Married|Finance|28202|0|1|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500016270|504626128|504628539|31|0|2|504632567|1|0|2|500882619|10|1|500009132|2128207318|4|1|500014681|-1|500007920, 500011315, 500011316, 500014681|-1|0|4|||12831|3|||1||2611337051335117774|0
M1038|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1061|Green||2014-04-01|2014-04-11|NaT||||34.9||1|1|1|1|M|Multi-race (Black & Hispanic)||12|No|Mother|28270|5|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||54|28110|Some College|Married|Self-Employed, Entrepreneur|28110|11|6|Relative|Relative|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|1|0|0|1|277|60|598|500000170|500017777|503207102|503208876|38|0|1|503688236|1|0|1|500757797|10|2|-2||3|1||-2|500011312|-2|0|10|||17161|11|||1||4726905079488957916|1161486385597736500
M1039|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-09-21|2016-10-31|NaT||||4.2||1|1|1|1|M|White||12|No|Mother|28031|6|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||28|28031|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|7|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504417121|504419373|1|0|1|504579745|1|0|1|500909172|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||3974159976843499574|458920933571351085
M1040|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|215|Green||2014-12-10|2014-12-18|2015-07-21|Child: Graduated|Child: Graduated||7.1||1|1|2|2|M|Black||12|No|Mother|28212|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||19|28213||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504143296|504145339|31|0|1|503540922|31|0|1|500803218|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1041|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|519|Green||2015-09-24|2015-10-05|NaT||||17.1||1|1|1|1|F|Black||12|No|Mother|28215|6|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Multi-Race (None of the above)||27|28269|Bachelors Degree|Single|Transport: Flight Attendant|28208|1|5|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504358312|504320644|31|0|2|504048355|7|0|2|500842174|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||8202428416367135871|2141487034287122220
M1042|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|93|Green|Cabarrus County|2016-11-22|2016-12-04|NaT||||3.1||1|1|1|1|F|Black||12|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||24|28262|Masters Degree|Single|Human Services: Social Worker|28027|0|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504937152|504939686|31|0|2|504797758|31|0|2|500930335|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|7061088365951887132|0
M1043|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|265|Green||2015-10-20|2015-10-20|2016-07-11|Volunteer: Time constraint|Volunteer: Time constraint||8.7||2|2|1|1|M|Black||12|No|Mother|28209|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||27|28208|Bachelors Degree|Single|Tech: Engineer|28202|3|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504474573|504476847|31|0|1|504349165|1|0|1|500849467|10|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M1044|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|96|Green||2016-09-23|2016-10-02|2017-01-06|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||3.2||2|2|2|2|M|Black||12|No|Mother|28209|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||23|28202|Bachelors Degree|Single|Business|28202|0|9|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504474573|504476847|31|0|1|504685043|1|0|1|500909932|10|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M1045|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2770|Green|Amachi|2009-07-27|2009-08-06|NaT||||91||1|1|1|1|M|Black||12|Yes|GrandMother|28273|4|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|Black||40|28273|No High School|Single|Business: Human Resources||2|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501806165|501806520|31|0|1|501706064|31|0|1|500375643|10|2|-2||2|1|500000294|-2||-2|0|10|||7446|3|||1|500000294|0|0
M1046|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|294|Green||2015-09-23|2015-10-07|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|2|2|M|Black||12|No|Mother|28208|7|One Parent: Female|$10,000 to $14,999||||Yes||School|General Community||RTBM|M|Black||44|28105|Masters Degree|Married|Business: Mgt, Admin|28202|3|6|Ally Financial|Workplace Partner|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500016270|504416598|504784888|31|0|1|502432606|31|0|1|500841768|7|1|500009132|2128207318|4|1||-2||-1|0|4|||12831|3|1209, 635|1|1||2611337051335117774|7044657180546140448
M1047|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|301|Green|PERL 2014-2016|2016-05-02|2016-05-10|NaT||||9.9||1|1|3|3|M|Multi-race (Black & White)||12|Yes|Mother|28215|6|One Parent: Female|$35,000 to $39,999||||No||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||57|28269|Bachelors Degree|Married|Finance: Accountant|28202|34|2|Omega Psi Phi|Fraternity/Sorority|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|502183411|502183840|36|0|1|500189229|31|0|1|500891295|10|2|-2||2|1|500000294, 500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||8694|14|||1|500014681|0|4203557099934965158
M1048|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1350|Yellow||2013-06-19|2013-06-26|NaT||||44.4||1|1|1|1|M|Black||12|No|Mother|28227|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||32|28262|Some College|Single|Business||0|5|United Way|Service Organization|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502787404|502788587|31|0|1|503485414|31|0|1|500701279|10|2|-2||2|2||-2||-2|0|10|||16263|6|||1||8452412398369747552|7044657180546140448
M1049|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|135|Green||2015-09-23|2015-10-07|2016-02-19|Child/Family: Moved|Child/Family: Moved||4.4||1|1|3|3|F|Black||12|No|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|Black||30|28270|Masters Degree|Single|Finance|28202|0|1|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504416752|504419004|31|0|2|504396349|31|0|2|500841764|10|1|500009132|2128207318|4|1||-1||-1|0|4|||16705|3|||1||2611337051335117774|0
M1050|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|217|Green|PERL 2014-2016|2014-09-15|2014-09-23|2015-04-28|Child: Changed school/site|Child: Changed school/site||7.1||1|1|2|2|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28206|5|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|M|White||50|28134||Single|Tech: Research/Design|28202|0|0|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|504025428|504027446|38|0|1|503911351|1|0|1|500776020|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1|500014681|7960300212314874874|0
M1051|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|287|Green||2015-09-23|2015-10-14|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.4||1|1|3|3|M|Multi-race (Black & Hispanic)||12|No|Mother|28208|6|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Site||Match Support|M|White||30|28202|Bachelors Degree|Single|Finance: Accountant|28202|2|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333764|504335986|38|0|1|503908898|1|0|1|500841780|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|2369272735379862405
M1052|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|236|Green||2015-12-01|2015-12-04|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||7.8||1|1|3|3|M|Black||12|No|Mother|28208|6|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||24|29708|Bachelors Degree|Single|Finance|28202|0|10|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504517710|504520011|31|0|1|504475369|1|0|1|500864201|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1053|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|127|Green||2016-02-29|2016-03-23|2016-07-28|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||4.2||1|1|3|3|F|Black||12|No|Mother|28208|6|One Parent: Female|Unknown||||No||School|General Site||Match Support|F|White||28|28203|Bachelors Degree|Single|Finance|28202|0|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504626092|504628503|31|0|2|504349844|1|0|2|500882091|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1054|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|284|Green||2015-10-01|2015-10-01|2016-07-11|Child: Changed school/site|Child: Changed school/site||9.3||1|1|2|2|F|Black||12|No|Mother|28213|6|Two Parent|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||25|28202|Bachelors Degree|Single|Tech: Computer/Programmer|28208|2|1|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504410223|504412474|31|0|2|504445343|1|0|2|500843871|10|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M1055|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|598|Green||2013-10-07|2013-10-11|2015-06-01|Child: Graduated|Child: Graduated||19.6||1|1|1|1|M|Black||12|No|Mother|28212|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||20|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503637786|503639746|31|0|1|503577771|1|0|1|500716450|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1056|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|615|Red|PERL 2014-2016|2015-06-17|2015-06-24|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.2||1|1|1|1|M|Black||12|Yes|Mother|28208|4|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi, PERL 2014-2016|Match Support|M|White||30|28202|Masters Degree|Single|Finance: Accountant|28202|0|6|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|504054004|504056028|31|0|1|504265163|1|0|1|500830573|10|2|-2||4|3|500000294, 500014681|-2||-2|34|2|||17159|12|||1|500014681|6407809237813394802|3402014428779854546
M1057|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|247|Green||2014-09-29|2014-09-30|2015-06-04|Child: Graduated|Child: Graduated||8.1||4|4|2|2|F|Black||12||Mother|28212||One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502097375|502097799|31|0|2|503901690|1|0|2|500778745|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1058|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|349|Green||2015-09-22|2015-10-06|2016-09-19|Child: Changed school/site|Child: Changed school/site||11.5||1|1|2|2|F|Black||12|No|Mother|28203|6|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Site||Match Support|F|White||32|28078|Bachelors Degree|Single|Business: Mgt, Admin|28202|1|4|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504410217|504412468|31|0|2|504359867|1|0|2|500841637|10|1|500009132|2128212899|4|1||-1||-1|0|3|||16705|3|||1||7276767778509034039|0
M1059|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|138|Green||2016-09-16|2016-10-20|NaT||||4.5||1|1|1|1|M|Black||12|No|GrandMother|28212|6|One Parent: Female|$10,000 to $14,999|||Y|No||School|General Community||Match Support|M|White||26|28210|Bachelors Degree|Married|Business: Sales|28277|0|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504592666|504595050|31|0|1|504625671|1|0|1|500908174|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||0|0
M1060|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|757|Green||2015-01-16|2015-02-09|NaT||||24.9||1|1|1|1|M|Black||12|No|Mother|28208|7|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||52|28211||Married|Unknown||0|0|United Way|Service Organization|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504176462|504178571|31|0|1|504109704|1|0|1|500808567|10|1|500000295|2128207319|2|1||-1||-1|0|4|||16263|6|||1||3935539763241716148|0
M1061|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|602|Green||2013-10-07|2013-10-08|2015-06-02|Child: Graduated|Child: Graduated||19.8||1|1|1|1|F|Hispanic||12|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|Match Support|F|White||20|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503418316|503420158|3|0|2|503493771|1|0|2|500716279|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1062|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2017-01-17|2017-01-30|NaT||||1.2||1|1|1|1|M|Black||12|No|Mother|28217|6|One Parent: Female|$25,000 to $29,999|||Y|No|BBBS National Site|Web Link|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|M|White||37|28203|Masters Degree|Single|Business: Mgt, Admin|28226|0|1|Radio|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504736266|504738712|31|0|1|504634630|1|0|1|500940290|10|2|-2||2|1|500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|34|2|||131|1|||1||194235582162093094|2876415545463317777
M1063|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|569|Green||2013-11-11|2013-11-12|2015-06-04|Volunteer: Moved|Volunteer: Moved||18.7||2|2|1|1|F|White||12|No|Mother|28211|3|Two Parent|Unknown||||No||School|General Site||Match Support|F|Asian||20|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503704203|503706168|1|0|2|503493888|4|0|2|500729897|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1064|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|226|Green||2015-10-09|2015-10-27|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.4||2|2|2|2|F|White||12|No|Mother|28211|3|Two Parent|Unknown||||No||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503704203|503706168|1|0|2|504297059|1|0|2|500846357|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1065|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|311|Red|PERL 2014-2016|2014-10-30|2014-11-24|2015-10-01|Volunteer: Time constraint|Volunteer: Time constraint||10.2||1|1|1|1|F|Black||12|No|Mother|28206|5|Two Parent|$10,000 to $14,999|||Y|Yes||Relative|General Community|PERL 2014-2016|Match Support|F|Black||44|28269||Single|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500013781|503995803|503997818|31|0|2|503963125|31|0|2|500790223|10|2|-2||4|3|500014681|-2|500014681|-2|0|3|||17159|12|||1|500014681|7960300212314874874|7044657180546140448
M1066|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|267|Green||2014-09-12|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|2|2|F|Black||12|No|Aunt|28205|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||39|28134|Masters Degree|Separated|Business: Human Resources|28202|1|0|Self|Self|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|504013115|504015130|31|0|2|503675532|1|0|2|500775709|10|1|500009132|2128173561|4|1||-1||-1|0|4|||7464|9|||1||7960300212314874874|0
M1067|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|560|Green||2014-01-14|2014-01-23|2015-08-06|Child/Family: Moved|Child/Family: Moved||18.4||1|1|1|1|M|Black||12|No|Mother|28212|4|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28277|Bachelors Degree|Divorced|Business|28273|4|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503547661|503549536|31|0|1|503731665|1|0|1|500742652|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1||7554307376683929204|4568161510412752900
M1068|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|613|Red||2015-02-18|2015-02-26|2016-10-31|Child/Family: Moved|Child/Family: Moved||20.1||1|1|1|1|M|Black||12|No|Mother|28269|5|One Parent: Female|$20,000 to $24,999|Yes: Active|No||No||Self|General Community||Match Support|M|White||34|28078|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28078|1|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503884921|503876064|31|0|1|504160910|1|0|1|500814243|10|2|-2||4|3||-2||-2|0|10|||46|2|||1||5367149751093883357|3501831218874457455
M1069|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|335|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-03-30|2016-04-06|NaT||||11||1|1|1|1|M|Black||12|No|Mother|28208|5|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Community||Match Support|M|White||32|28203|Juris Doctorate (JD)|Single|Law: Lawyer|28277|1|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|503952082|503954090|31|0|1|504546069|1|0|1|500887070|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|3|||46|2|||1|500007920, 500011315, 500011316|4208486535559819469|0
M1070|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|572|Green||2013-10-15|2013-11-08|2015-06-03|Child: Graduated|Child: Graduated||18.8||1|1|1|1|F|Hispanic||12|No|Mother|28211|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503629807|503631746|3|0|2|503603514|1|0|2|500719608|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1071|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|742|Green|PERL 2014-2016|2015-02-12|2015-02-24|NaT||||24.4||1|1|1|1|M|Black||12|No|Mother|28216|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||50|28211|Juris Doctorate (JD)|Married|Law: Lawyer|28211|17|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500017732|503533041|503534897|31|0|1|504183712|1|0|1|500813495|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||7496|10|||1|500014681|3935539763241716148|1786514887916898235
M1072|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2095|Green|Project Big|2011-06-02|2011-06-12|NaT||||68.8||1|1|1|1|F|Black||12|No|GrandMother|28208|1|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|Project Big|Match Support|F|White||28|28209|Bachelors Degree|Single|Business: Sales|28277|0|9|Self|Self|Big|General Community|Amachi, Project Big|Match Support|1|0|0|1|277|60|598|500000170|500020910|502552445|502552891|31|0|2|502545537|1|0|2|500539524|10|2|500004641||2|1|500004640|-2|500000294, 500004640|-2|0|4|||7464|9|||1|500004640|7869308672550505300|0
M1073|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|603|Green||2013-10-07|2013-10-07|2015-06-02|Child: Graduated|Child: Graduated||19.8||3|3|1|1|F|Hispanic||12|No|Mother|28212||One Parent: Female|Unknown||||No||School|General Site||Match Support|F|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502395420|502395858|3|0|2|503497477|1|0|2|500716286|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1074|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|721|Green|PERL 2014-2016|2015-03-16|2015-03-17|NaT||||23.7||1|1|1|1|M|Black||12|No|Aunt|28216|7|One Parent: Female|$40,000 to $44,999||||Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||33|28208|Masters Degree|Married|Finance|28202|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|503946469|503948477|31|0|1|504188283|31|0|1|500818848|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681|9134125726462845918|529594392811859839
M1075|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|518|Green||2015-09-22|2015-10-06|NaT||||17||1|1|1|1|F|Black||12|No|Mother|28208|7|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|PERL 2014-2016|Match Support|F|White||24|28107|Bachelors Degree|Single|Tech: Computer/Programmer|28208|0|7|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504410249|504412500|31|0|2|504369534|1|0|2|500841376|10|1|500009132|2128212899|2|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M1076|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|155|Green||2016-09-29|2016-10-03|NaT||||5.1||1|1|2|2|M|Black||12|No|GrandMother|28217|7|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|M|White||28|28211|Bachelors Degree|Married|Tech: Computer/Programmer|28202|4|6|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504869115|504871634|31|0|1|504349938|1|0|1|500911559|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||8568001799025358453|0
M1077|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|130|Green||2016-10-28|2016-10-28|NaT||||4.3||1|1|1|1|M|White||12|No|Mother|28226|6|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|M|White||31|28205|Bachelors Degree|Single|Real Estate: Realtor|28202|1|6|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504436181|504438437|1|0|1|504741299|1|0|1|500921121|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||0|6694016660882153370
M1078|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|476|Green|PERL 2014-2016, Cabarrus County|2015-11-10|2015-11-17|NaT||||15.6||1|1|1|1|M|White||12|Yes|Mother|28025|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||32|28025|Bachelors Degree||Business: Sales||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|503821686|503823656|1|0|1|504460050|1|0|1|500858397|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7496|10|||1|500014681, 500016374|5064856656261650513|7044657180546140448
M1079|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|225|Green||2014-10-04|2014-10-22|2015-06-04|Child: Graduated|Child: Graduated||7.4||2|2|2|2|F|Hispanic||12|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503229410|503231198|3|0|2|503493684|1|0|2|500780613|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1080|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|519|Green||2015-09-22|2015-10-05|NaT||||17.1||1|1|3|3|M|Black||12|No|Mother|28217|7|Two Parent|$10,000 to $14,999|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|Black||29|28273|Bachelors Degree|Married|Tech: Computer/Programmer||5|0|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504396333|504045278|31|0|1|502542324|31|0|1|500841349|10|1|500009132|2128212899|2|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||8568001799025358453|0
M1081|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2286|Green||2010-11-15|2010-12-03|NaT||||75.1||1|1|1|1|F|Black||12|No|Mother|28213|1|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||40|28269|Bachelors Degree|Married|Tech: Management|28255|1|9|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|502278991|502279417|31|0|2|502263116|31|0|2|500494784|10|2|-2||2|1||-2|500000294|-2|6854|8|||6247|12|||1||0|7044657180546140448
M1082|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|600|Green||2013-10-08|2013-10-09|2015-06-01|Child: Graduated|Child: Graduated||19.7||3|3|1|1|M|Hispanic||12|Yes|Mother|28270|1|One Parent: Female|Unknown||||Yes||School|General Site|Amachi|Match Support|M|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502335396|502335831|3|0|1|503507119|1|0|1|500717197|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1083|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|633|Green||2013-11-10|2013-11-12|2015-08-07|Volunteer: Moved|Volunteer: Moved||20.8||2|2|1|1|F|Hispanic||12|Yes|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||20|28211||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503704276|503706241|3|0|2|503507098|1|0|2|500729563|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1084|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|231|Green||2015-10-09|2015-10-22|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.6||2|2|2|2|F|Hispanic||12|Yes|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503704276|503706241|3|0|2|504306171|1|0|2|500846366|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1085|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|225|Green|PERL 2014-2016|2016-07-08|2016-07-25|NaT||||7.4||1|1|1|1|F|Black||12|No|Mother|28216|6|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||29|28269|Some College|Single|Business: Sales|28262|1|0|Community Engagement|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504628514|504630931|31|0|2|504599441|31|0|2|500899221|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||18809|8|||1|500014681|806697982905023857|7044657180546140448
M1086|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|296|Green||2015-09-23|2015-10-05|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|2|2|F|Hispanic||12|No|Mother|28208|6|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||33|28209|Bachelors Degree|Single|Finance|28202|4|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504333802|504336025|3|0|2|504354941|1|0|2|500841763|10|1|500009132|2128207318|4|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1087|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|12|Green||2017-02-23|2017-02-23|NaT||||0.4||1|1|1|1|M|Black||12|No|Foster Parent|28215|6|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|M|Black||25|28223|Bachelors Degree|Single|Business|28202|1|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500013781|504463138|504465396|31|0|1|504819424|31|0|1|500947979|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||1421169092898167719|7044657180546140448
M1088|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|190|Green||2015-01-21|2015-01-29|2015-08-07|Child: Graduated|Child: Graduated||6.2||1|1|3|3|F|Black||12|No|Mother|28211|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504176233|504178342|31|0|2|503500482|1|0|2|500809250|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1089|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|250|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-06-16|2016-06-30|NaT||||8.2||1|1|1|1|F|Black||12|No|Mother|28211|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||27|28205|Some College||Medical|28269|0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504471617|504473895|31|0|2|504458762|31|0|2|500897003|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1|500007920, 500011315, 500011316|8758769076374727509|1545381051186164660
M1090|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|421|Green|PERL 2014-2016|2015-11-04|2015-11-23|2017-01-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.8||1|1|1|1|M|Black||12|No|GrandMother|28215|6|Grandparents|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI, PERL 2014-2016|Enrollment|M|Black||30|28262|Some College|Married|Architect|28207|0|6|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment|Match Support|0|1|1|0|277|60|598|500000170|500021785|502458458|502458905|31|0|1|504387453|31|0|1|500855881|5|2|-2||4|1|500005291, 500014681|-2|500011316, 500014681|-2|0|5|||46|2|||1|500014681|5441374193599827162|3274057295643004474
M1091|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1461|Red||2013-02-14|2013-02-28|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||48||1|1|1|1|M|Black||12|No|Mother|28211|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||31|28210|Bachelors Degree|Single|Business: Engineer||5|0|Relative|Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502979757|502981210|31|0|1|503161988|1|0|1|500682191|10|2|-2||4|3||-2||-2|0|10|||17161|11|||1||421482027904269589|8247408236389589972
M1092|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|501|Green|PERL 2014-2016, Cabarrus County|2015-09-29|2015-10-23|NaT||||16.5||3|3|1|1|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28083|2|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|M|White||39|28027|Masters Degree|Married|Business|28269|9|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|502234905|502777258|38|0|1|504334608|1|0|1|500843097|10|2|500016307||2|1|500000294, 500014681, 500016374|-2|500014681, 500016374|-2|0|10|||17159|12|||1|500014681, 500016374|370020301266015142|0
M1093|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1359|Green|Amachi|2011-11-30|2011-12-05|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||44.6||3|3|1|1|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28083|2|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|M|White||36|28097|Masters Degree|Divorced|Finance|28026|7|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|502234905|502777258|38|0|1|502799047|1|0|1|500583119|10|2|-2||4|1|500000294, 500014681, 500016374|-2||-2|0|10|||7671|13|||1|500000294|370020301266015142|0
M1094|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|469|Green||2015-11-13|2015-11-24|NaT||||15.4||1|1|1|1|M|Black||12|No|Mother|28211|5|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||48|28105||Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504227502|504229617|31|0|1|504460839|31|0|1|500859784|10|2|-2||2|1|500000294|-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1||976372749760822282|2077565980961547475
M1095|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|361|Green||2014-10-23|2014-11-21|2015-11-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.9||4|4|1|1|F|Hispanic||12|No|Mother|28027|4|Other/Unknown|Unknown||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||40|28027||Single|Business|28027|2|0|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500012459|503270485|503272299|3|0|2|504039802|31|0|2|500787379|10|1|500000295|2128212924|4|1|500014681, 500016374|-2||-1|0|4|||7464|9|||1||3232906304025417619|0
M1096|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|381|Green|PERL 2014-2016, Cabarrus County|2016-02-19|2016-02-20|NaT||||12.5||4|4|1|1|F|Hispanic||12|No|Mother|28027|4|Other/Unknown|Unknown||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||28|28075|Bachelors Degree|Single|Education: Teacher|28025|2|6|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|503270485|503272299|3|0|2|504574450|1|0|2|500880422|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||46|2|||1|500014681, 500016374|3232906304025417619|0
M1097|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|370|Red|PERL 2014-2016|2016-01-11|2016-02-09|2017-02-13|Volunteer: Moved|Volunteer: Moved||12.2||1|1|1|1|M|White||12|No|Mother|28214|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community|PERL 2014-2016|Match Support|M|White||56|28012|Some College|Married|Business: Mgt, Admin|33401|4|7|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500013781|504231267|504233379|1|0|1|504379684|1|0|1|500871125|10|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|3|||46|2|||1|500014681|9076057728106637014|0
M1098|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|813|Green|PERL 2014-2016|2014-11-21|2014-12-15|NaT||||26.7||1|1|1|1|F|Black||12|No|Mother|28208|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||37|28227|Associate Degree|Single|Student: College|28223|1|0|Web in a Box, v1|Web Link|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500008321|503978153|503980164|31|0|2|504039547|31|0|2|500798168|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||15467|2|||1|500014681|6368218764956286027|0
M1099|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|160|Green|PERL 2014-2016|2016-09-13|2016-09-28|NaT||||5.3||1|1|1|1|F|Black||12|No|Mother|28269||One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||28|28203|Bachelors Degree|Single|Finance: Banking|28203|0|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504489376|504491661|31|0|2|504604779|1|0|2|500907166|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||7464|9|||1|500014681|8568001799025358453|7341607196510895077
M1100|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1698|Green||2012-07-09|2012-07-13|NaT||||55.8||2|2|1|1|M|Black||12|No|Mother|28206|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Site||Match Support|M|White||37|28209|Bachelors Degree|Married|Unemployed|22202|9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502933371|502934793|31|0|1|503080292|1|0|1|500623322|10|2|-2||2|1||-1||-2|0|10|||7496|10|||1||7960300212314874874|0
M1101|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|267|Green||2014-09-15|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||2|2|3|3|M|Black||12|No|Mother|28206|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Site||Match Support|M|White||30|28273|Bachelors Degree|Single|Finance|28202|1|8|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|502933371|502934793|31|0|1|503911379|1|0|1|500776006|10|1|500009132|2128173561|4|1||-1||-1|0|10|||12831|3|||1||7960300212314874874|0
M1102|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|93|Red||2016-11-11|2016-12-04|NaT||||3.1||1|1|1|1|M|White||12|No|Mother|29715|6|One Parent: Female|$30,000 to $34,999||||No||Self|General Site||Match Support|M|White||31|28277|Bachelors Degree|Married|Finance: Accountant|29715|1|6|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504886657|504889177|1|0|1|504807149|1|0|1|500927129|10|1|500009132|2128233620|2|3||-1||-1|0|10|||7464|9|||1||1174067921639243853|4314330004570465916
M1103|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|509|Green||2015-03-16|2015-03-20|2016-08-10|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||16.7||1|1|1|1|F|Black||12|No|Father|28205|6|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|F|White||33|28227|Associate Degree|Divorced|Medical: Healthcare Worker|28213|1|4|Local TV|Media|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504200641|504202752|31|0|2|504222624|1|0|2|500818777|10|1|500000295|2128173561|4|1||-1||-1|0|4|||7438|1|||1||7960300212314874874|0
M1104|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|862|Red|PERL 2014-2016|2014-10-17|2014-10-20|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||28.3||3|3|1|1|F|Black||12|Yes|Mother|28211|4|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|F|Black||58|28269|Bachelors Degree|Married|Self-Employed, Entrepreneur|28269|26|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500008321|502173768|503800801|31|0|2|503831898|31|0|2|500784859|10|2|-2||4|3|500000294, 500014681|-2|500014681|-2|0|4|||7464|9|||1|500014681|7807202941877299922|0
M1105|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|426|Green||2014-03-18|2014-03-28|2015-05-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14||1|1|3|3|F|Black||12|Yes|Mother|28203|4|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|Match Support|F|White||36|28104|Bachelors Degree|Married|Business: Sales||2|4|Self|Self|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|503807556|503809533|31|0|2|502105224|1|0|2|500755253|10|1|-1||4|1|500000294|-1|500000294|-1|0|4|||7464|9|||1||8981704271528751143|0
M1106|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|862|Green|PERL 2014-2016|2014-09-25|2014-10-27|NaT||||28.3||1|1|1|1|M|Black||12|No|Mother|28215|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28205|Bachelors Degree|Single|Finance: Accountant|28202|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500013781|503636487|503665377|31|0|1|503899296|1|0|1|500778337|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681|6724463016047116758|0
M1107|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|763|Red||2014-08-07|2014-08-27|2016-09-28|Volunteer: Time constraint|Volunteer: Time constraint||25.1||1|1|1|1|M|Hispanic||12|No|Mother|28277|5|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|Some Other Race||31|28270|Bachelors Degree|Married|Real Estate: Realtor|28110|0|5|Man Up Campaign|Media|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|1|0|1|0|277|60|598|500000170|500008321|503590328|503592205|3|0|1|503874645|41|0|1|500771736|10|2|-2||4|3||-2|500011312|-2|0|10|||17101|1|||1||3090721985630916616|2156718237896110088
M1108|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1964|Green||2011-10-04|2011-10-21|NaT||||64.5||2|2|1|1|F|Black||12|No|Mother|28216|3|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Mgt, Admin|28204|0|9|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|502223076|502223507|31|0|2|502694717|1|0|2|500560829|10|2|-2||2|1|500004640|-2||-2|0|10|||7464|9|||1||7869308672550505300|0
M1109|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|383|Yellow||2014-07-02|2014-08-28|2015-09-15|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12.6||2|2|1|1|F|Black||12|No|Mother|28273|6|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||34|28214|Some College|Single|Transport: Driver|28273|9|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503895740|503897736|31|0|2|503765053|31|0|2|500768490|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||194235582162093094|3184471850140890355
M1110|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|286|Green||2015-12-15|2016-01-06|2016-10-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||9.4||2|2|1|1|F|Black||12|No|Mother|28273|6|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||30|28210|Bachelors Degree|Single|Business|28211|4|6|Community Engagement|Special Event|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500020910|503895740|503897736|31|0|2|504364485|1|0|2|500867759|10|2|-2||4|1||-2||-2|0|10|||18809|8|||1||194235582162093094|3184471850140890355
M1111|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|742|Green|PERL 2014-2016|2015-02-18|2015-02-24|NaT||||24.4||1|1|1|1|F|Black||12|Yes|Mother|28217|6|One Parent: Female|$20,000 to $24,999||||No|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||28|28205|Bachelors Degree|Single|Journalist/Media|28202|4|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504171035|504173143|31|0|2|504150234|1|0|2|500814425|10|2|-2||2|1|500014681|-2|500014681|-2|34|2|||46|2|||1|500014681|3974159976843499574|7044657180546140448
M1112|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1348|Green|Cabarrus County|2013-06-05|2013-06-28|NaT||||44.3||1|1|2|2|M|Black||12|No|Mother|28083|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||60|28027|Bachelors Degree|Separated|Insurance|28262|24|0|Local Radio|Media|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502761742|502762654|31|0|1|503041890|1|0|1|500699565|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7437|1|||1|500016374|643003066716863548|4058276550489173605
M1113|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|265|Green||2014-09-12|2014-09-25|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||1|1|1|1|F|Black||12|No|Mother|28206|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||26|28202|Masters Degree|Single|Tech: Research/Design|28202|0|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504013104|504015119|31|0|2|503933411|1|0|2|500775718|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M1114|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|232|Green||2015-11-02|2015-12-08|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||7.6||1|1|1|1|M|Black||12|No|Mother|28208|6|One Parent: Female|$15,000 to $19,999||||Yes||Relative|General Site||Match Support|M|Black||50|28216|Bachelors Degree|Married|Tech: Management|28202|0|7|Ally Financial|Workplace Partner|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500016270|504333758|504335980|31|0|1|504484385|31|0|1|500855108|10|1|500009132|2128207318|4|1||-1|500007920, 500011315, 500011316|-1|0|3|||12831|3|||1||2611337051335117774|2710650624457676912
M1115|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|505|Green||2015-09-22|2015-10-19|NaT||||16.6||1|1|1|1|F|Black||12|Yes|Mother|28203|7|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||29|28023|Masters Degree|Married|Finance: Accountant|28202|1|4|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504437000|504429531|31|0|2|503979153|1|0|2|500841337|10|1|500009132|2128212899|2|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M1116|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-22|2015-10-01|NaT||||17.2||1|1|1|1|F|Black||12|Yes|Mother|28203|7|One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|F|Black||26|28269|Masters Degree|Single|Tech: Computer/Programmer|28202|0|3|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504427276|504429531|31|0|2|504354996|31|0|2|500841643|10|1|500009132|2128212899|2|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M1117|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|853|Green||2014-06-16|2014-07-11|2016-11-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28||1|1|1|1|M|Black||12|No|Mother|28211|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|M|White||27|28226|Bachelors Degree|Single|Tech: Research/Design|28269|0|8|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503512877|503514748|31|0|1|503893014|1|0|1|500766726|5|2|-2||4|1||-2||-2|0|10|||17101|1|||1||5533634913091743658|0
M1118|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|237|Green|PERL 2014-2016|2014-09-25|2014-10-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||7.8||1|1|1|1|F|Black||12|No|Mother|28206|5|Two Parent|Unknown||||No||School|General Site|PERL 2014-2016|Match Support|F|Black||35|28202|Bachelors Degree|Single|Tech: Computer/Programmer|28202|10|0|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|504039826|504041844|31|0|2|503980178|31|0|2|500778282|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1|500014681|7960300212314874874|0
M1119|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|189|Green||2016-08-03|2016-08-30|NaT||||6.2||1|1|3|3|M|Black||12|No|Mother|28262|6|One Parent: Female|$20,000 to $24,999||||Yes||School|General Community||Match Support|M|Black||25|28269|Masters Degree|Single|Finance|28202|0|1|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|504275306|504277506|31|0|1|504359606|31|0|1|500901552|10|2|-2||2|1||-2|500014681|-1|0|4|||12831|3|||1||0|7674215580094440446
M1120|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|812|Green||2014-12-02|2014-12-16|NaT||||26.7||1|1|1|1|F|Black||12|No|Mother|28216|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||25|28209|Bachelors Degree|Single|Finance|28202|1|3|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020752|504038458|504040320|31|0|2|503971368|1|0|2|500800323|10|2|-2||2|1||-2|500000294|-2|0|10|||17159|12|||1||7883015200677941272|0
M1121|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|418|Green|PERL 2014-2016|2015-03-02|2015-03-12|2016-05-03|Volunteer: Time constraint|Volunteer: Time constraint||13.7||1|1|2|2|F|Black||12|No|Mother|28206|6|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Enrollment|F|White||55|28277|Associate Degree|Single|Law: Paralegal|28217|0|8|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500016270|504200631|504202742|31|0|2|503404737|1|0|2|500816351|5|1|500000295|2128173561|4|1|500014681|-1|500000294|-2|0|4|||7464|9|||1|500014681|7960300212314874874|0
M1122|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|294|Green||2015-09-21|2015-10-07|2016-07-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.7||1|1|2|2|F|Black||12|No|Mother|28206|6|One Parent: Female|Unknown||||Yes||Relative|General Site|PERL 2014-2016|Match Support|F|Black||31|28277|Associate Degree|Single|Finance: Auditor|28202|0|3|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504416771|504419023|31|0|2|504349862|31|0|2|500841103|10|1|500009132|2128207318|4|1|500014681|-1|500014681|-1|0|3|||12831|3|||1||2611337051335117774|0
M1123|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1801|Red||2010-07-12|2010-08-25|2015-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||59.2||1|1|1|1|M|Black||12|No|Mother|28210||One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||45|28211|Masters Degree|Married|Finance: Banking||11|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501314348|501314626|31|0|1|502205797|1|0|1|500460633|10|2|-2||4|3||-2||-2|0|10|||2230|7|||1||0|7151546326379863072
M1124|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|523|Green||2015-09-23|2015-10-01|NaT||||17.2||1|1|2|2|F|Black||12|No|Mother|28217|7|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|F|White||29|28031|Masters Degree|Married|Tech: Support, Writing|28202|2|5|Duke Energy|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504396318|504398558|31|0|2|503605621|1|0|2|500841724|10|1|500009132|2128212899|2|1|500014681|-1|500014681|-1|0|4|||16705|3|||1||7276767778509034039|0
M1125|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|111|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-01-14|2016-01-30|2016-05-20|Volunteer: Moved|Volunteer: Moved||3.6||2|2|1|1|F|Black||12|No|Mother|28214|5|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||32|28208|Bachelors Degree|Single|Journalist/Media||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503976557|503978568|31|0|2|504365048|1|0|2|500871811|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|500007920, 500011315, 500011316|0|3198188609986797983
M1126|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|250|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-06-16|2016-06-30|NaT||||8.2||2|2|1|1|F|Black||12|No|Mother|28214|5|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||26|28203|Bachelors Degree|Married|Business: Mgt, Admin|29707|0|4|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|503976557|503978568|31|0|2|504538747|1|0|2|500896984|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||18809|8|||1|500007920, 500011315, 500011316|0|3198188609986797983
M1127|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|686|Green|PERL 2014-2016|2015-02-23|2015-02-26|2017-01-12|Volunteer: Time constraint|Volunteer: Time constraint||22.5||1|1|1|1|F|Black||12|No|Mother|28213|5|One Parent: Female|$45,000 to $49,999||||Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Enrollment|F|Black||21|28269|Some College|Single|Business: Sales|28269|0|5|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500017732|504038255|504040273|31|0|2|504034443|31|0|2|500814943|5|2|-2||4|1|500014681|-2|500014681|-2|34|2|||46|2|||1|500014681|7679812394383646966|8408514790530965815
M1128|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|487|Green||2014-01-21|2014-01-31|2015-06-02|Child: Graduated|Child: Graduated||16||2|2|2|2|F|Black||12|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||20|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503254146|503255951|31|0|2|503509874|1|0|2|500744048|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1129|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|602|Green||2014-10-07|2014-10-09|2016-06-02|Child: Changed school/site|Child: Changed school/site||19.8||1|1|1|1|M|Black||12|No|Mother|28212|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020908|504049432|504044051|31|0|1|503908413|31|0|1|500781517|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1130|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|354|Green||2015-10-01|2015-10-01|2016-09-19|Child: Changed school/site|Child: Changed school/site||11.6||1|1|2|3|F|Black||12|No|Mother|28210|6|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||49|28278|Masters Degree|Single|Business|28202|12|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504410241|504412492|31|0|2|503605964|1|0|2|500843880|10|1|500009132|2128212899|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M1131|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|997|Green||2013-11-15|2013-11-25|2016-08-18|Volunteer: Time constraint|Volunteer: Time constraint||32.8||1|1|1|1|F|Black||12|Yes|Mother|28269|4|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|White||53|28227|Some College|Married|Customer Service|28105|30|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|503701025|501153063|31|0|2|503576358|1|0|2|500731543|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1||7960300212314874874|0
M1132|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|204|Green||2014-10-21|2014-11-25|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||6.7||1|1|1|1|M|Black||12|No|Mother|28206|4|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||31|28120|Masters Degree|Married|Finance|28202|0|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504040012|504042030|31|0|1|503935151|1|0|1|500785775|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M1133|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|112|Red||2015-11-10|2015-11-19|2016-03-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.7||4|4|1|1|F|Black||12|No|Mother|28081|5|One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|White||31|28081|Masters Degree|Married|Education|28223|1|10|Current/Previous Big|Other Big|Big|General Community|Amachi, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020753|502789637|502790820|31|0|2|504034331|1|0|2|500858188|10|2|-2||4|3|500016374|-2|500000294, 500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||2362631343152316267|7044657180546140448
M1134|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|701|Yellow||2013-09-03|2013-09-23|2015-08-25|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||23||4|4|2|2|F|Black||12|No|Mother|28081|5|One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|Black||30|28027|Masters Degree|Married|Unemployed|28027|2|5|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500012459|502789637|502790820|31|0|2|503542037|31|0|2|500708902|10|2|-2||4|2|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||7464|9|||1||2362631343152316267|7044657180546140448
M1135|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|270|Green|Cabarrus County|2016-05-24|2016-06-10|NaT||||8.9||4|4|1|1|F|Black||12|No|Mother|28081|5|One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|Black||25|28025|Bachelors Degree|Single|Insurance|28213|1|10|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|502789637|502790820|31|0|2|504703410|31|0|2|500894186|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|2362631343152316267|7044657180546140448
M1136|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1102|Green||2013-04-02|2013-04-26|2016-05-02|Volunteer: Time constraint|Volunteer: Time constraint||36.2||1|1|1|1|F|Black||12|Yes|Mother|28212|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||36|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28202|5|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|503355095|503356940|31|0|2|503373533|31|0|2|500691042|10|2|-2||4|1|500000294|-2||-2|0|10|||7496|10|||1||0|1407725786000053166
M1137|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1077|Yellow||2014-03-04|2014-03-26|NaT||||35.4||1|1|1|1|M|Black||12|No|Mother|28105|2|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||31|28226|Bachelors Degree|Single|Finance: Accountant|28217|4|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503401214|503403071|31|0|1|503758808|1|0|1|500752693|10|2|-2||2|2||-2||-2|0|10|||7496|10|||1||7134583514356134698|3714886275549507192
M1138|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|491|Yellow||2015-01-05|2015-01-12|2016-05-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.1||1|1|1|1|M|Black||12|No|GrandMother|28217|4|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|M|Black||31|28273|Bachelors Degree|Single|Finance|28209|0|3|Man Up Campaign|Media|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500013781|504133883|504135920|31|0|1|503868128|31|0|1|500806524|10|1|500000295|2128173557|4|2||-1||-1|0|3|||17101|1|||1||8981704271528751143|0
M1139|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|389|Green||2014-01-07|2014-01-23|2015-02-16|Volunteer: Time constraint|Volunteer: Time constraint||12.8||1|1|1|1|F|Hispanic||12|No|Mother|28217|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||51|29707|Juris Doctorate (JD)|Widowed|Law: Lawyer|28273|15|0|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016847|503756537|503758509|3|0|2|503403281|1|0|2|500741577|10|1|500000295|2128173557|4|1||-1||-1|0|4|||7464|9|||1||8981704271528751143|0
M1140|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|601|Green||2013-10-07|2013-10-08|2015-06-01|Child: Graduated|Child: Graduated||19.7||1|1|1|1|M|Black||12|Yes|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|Match Support|M|White||20|28205|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503281891|503263744|31|0|1|503507494|1|0|1|500716280|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1141|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Inactive|Match Support|517|Green||2015-09-23|2015-10-07|NaT||||17||2|2|1|1|F|Black||12|No|Mother|28208|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|Project Big|Match Support|F|Black||36|28213|Masters Degree|Married|Finance|28202|3|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500008321|502234486|502234907|31|0|2|504359670|31|0|2|500841766|10|1|-1||3|1|500004640|-1||-1|0|4|||12831|3|||1||2611337051335117774|5656517387001249169
M1142|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|620|Green||2013-12-31|2014-01-17|2015-09-29|Child: Graduated|Child: Graduated||20.4||3|3|2|2|F|Black||12||Mother|28031|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||70|28031||Divorced|Consultant||0|0|Self|Self|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017786|502813499|502814776|31|0|2|503633204|1|0|2|500740854|10|1|500000295|2128173570|4|1||-1|500000294|-1|0|4|||7464|9|||1||8034889377453131101|0
M1143|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|263|Green||2015-01-05|2015-01-30|2015-10-20|Child/Family: Moved|Child/Family: Moved||8.6||1|1|1|1|M|Hispanic||12|No|Mother|28217|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Hispanic||60|28104|Bachelors Degree|Widowed|Retired||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500020753|504133877|504135914|3|0|1|503908101|3|0|1|500806523|10|1|500000295|2128173557|4|1||-1||-1|0|4|||7496|10|||1||8981704271528751143|0
M1144|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|173|Green|PERL 2014-2016|2016-09-01|2016-09-15|NaT||||5.7||1|1|2|2|M|Black||12|No|Mother|28215|5|One Parent: Female|$40,000 to $44,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|Black||54|28262|Bachelors Degree|Married|Business||7|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504310625|504312843|31|0|1|503442370|31|0|1|500905889|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||7464|9|||1|500014681|7284449467126735125|7399582438680751686
M1145|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|456|Green||2015-09-22|2015-10-05|2017-01-03|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||15||1|1|3|3|M|Hispanic||12|No|Father|28217|7|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|M|White||30|29707|Bachelors Degree|Married|Business: Engineer|28202|6|2|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504439749|504442005|3|0|1|503605644|1|0|1|500841647|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7276767778509034039|0
M1146|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-17|2016-12-02|NaT||||3.1||1|1|4|4|M|Black||12|Yes|Mother|29715|6|Two Parent|$50,000 to $59,999||||No||Self|General Site||Match Support|M|Black||44|29732|High School Graduate|Married|Business|28217|5|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504886640|504889160|31|0|1|503754104|31|0|1|500929268|10|1|500009132|2128233620|2|1||-1||-1|0|10|||11247|3|||1||1174067921639243853|386356889061704511
M1147|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|438|Yellow||2015-02-09|2015-02-09|2016-04-22|Child: Changed school/site|Child: Changed school/site||14.4||1|1|3|3|M|Multi-Race (None of the above)||12|No|Mother|28208|6|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|Black||26|29730|Some High School|Married|Business: Sales|28217|1|6|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504205445|504207556|7|0|1|503796968|31|0|1|500812652|10|1|500000295|2128207319|4|2||-1||-1|0|4|||46|2|||1||3935539763241716148|0
M1148|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|264|Green||2014-09-22|2014-09-25|2015-06-16|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||1|1|1|1|M|Black||12|No|Mother|28205|4|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||40|28209|Bachelors Degree|Married|Business|28202|5|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504030001|504032019|31|0|1|503935202|1|0|1|500777116|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M1149|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2133|Green|Amachi|2011-04-21|2011-05-05|NaT||||70.1||1|1|1|1|M|Black||12|Yes|Mother|28216|1|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||32|28104|Bachelors Degree|Single|Business|28216|5|3|Relative|Relative|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502245343|502245774|31|0|1|502526001|1|0|1|500532810|10|2|500003586||2|1|500000294|-2||-2|0|10|||17161|11|||1|500000294|0|9181709468273956350
M1150|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|547|Green||2015-04-20|2015-05-01|2016-10-29|Child: Graduated|Child: Graduated||18||1|1|1|1|F|Hispanic||12|No|Mother|28217|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||31|28277|Bachelors Degree|Divorced|Business: Mgt, Admin|28277|1|5|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500013781|504133872|504135909|3|0|2|504225360|1|0|2|500824003|10|1|500000295|2128173557|4|1||-1||-1|0|4|||17159|12|||1||8981704271528751143|0
M1151|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|369|Green||2014-10-04|2014-10-09|2015-10-13|Volunteer: Time constraint|Volunteer: Time constraint||12.1||2|2|1|1|M|Hispanic||12|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504041825|504043821|3|0|1|503907538|1|0|1|500780593|10|1|500000296|2128173564|4|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1152|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|240|Green||2015-10-13|2015-10-13|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.9||2|2|2|2|M|Hispanic||12|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|M|White||18|28277|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504041825|504043821|3|0|1|504303741|1|0|1|500847619|10|1|500000296|2128173564|4|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1153|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-21|2016-10-31|NaT||||4.2||1|1|1|1|M|Multi-race (Black & White)||12|No|Mother|28078|5|One Parent: Female|$40,000 to $44,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||31|28078|Some College|Married|Business: Sales|28078|0|5|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504416044|504418296|36|0|1|504623074|1|0|1|500918304|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||927920773840777760|7269080898586176194
M1154|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1148|Red||2013-06-10|2013-06-17|2016-08-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||37.7||1|1|1|1|M|Black||12||Mother|28217|2|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||48|28273|Some College|Divorced|Transport: Driver|29730|3|0|TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503472232|503474098|31|0|1|503444888|31|0|1|500700046|10|2|-2||4|3||-2||-2|34|2|||130|1|||1||5386346637278076349|7044657180546140448
M1155|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|1|1|F|Hispanic||12|No|Father|28208|6|One Parent: Female|Less than $10,000||||Yes||School|General Site|PERL 2014-2016|Match Support|F|White||26|28203|Bachelors Degree|Single|Business|28202|0|3|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861201|504863720|3|0|2|504804012|1|0|2|500911904|10|1|500009132|2128207318|2|1|500014681|-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1156|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|619|Green|Cabarrus County|2015-06-15|2015-06-27|NaT||||20.3||1|1|1|1|M|Multi-race (Black & Asian)||12|No|Mother|28025|7|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Asian||32|28025|Bachelors Degree|Married|Tech: Sales, Mktg|28202|8|9|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi, Cabarrus County, mentor2.0|Match Support|0|1|0|1|277|60|598|500000170|500022817|504051660|504053684|39|0|1|504277513|4|0|1|500830267|10|2|500016307||2|1|500016374|-2|500000294, 500014505, 500016374|-2|0|10|||7462|13|||1|500016374|0|887254134148570071
M1157|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|602|Green||2014-10-04|2014-10-09|2016-06-02|Child: Changed school/site|Child: Changed school/site||19.8||1|1|1|1|M|Black||12|No|Mother|28211|4|One Parent: Female|Unknown||||Yes||School|General Site|Amachi|Match Support|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020909|504049365|504051389|31|0|1|503908435|1|0|1|500780584|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1158|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|661|Green||2013-10-08|2013-10-15|2015-08-07|Volunteer: Moved|Volunteer: Moved||21.7||2|2|1|1|F|Hispanic||12|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503629858|504178353|3|0|2|503507250|1|0|2|500717193|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1159|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|247|Green||2015-10-06|2015-10-06|2016-06-09|Child: Changed school/site|Child: Changed school/site||8.1||2|2|2|2|F|Hispanic||12|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503629858|504178353|3|0|2|504303791|1|0|2|500844553|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1160|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1511|Yellow|Amachi|2011-12-20|2011-12-20|2016-02-08|Volunteer: Moved|Volunteer: Moved||49.6||3|3|2|2|F|Black||12|Yes|Mother|28227|6|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Some Other Race||75|28213|Some College|Widowed|Human Services||20|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020990|502347820|502348258|31|0|2|502419409|41|0|2|500588112|10|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294|8758769076374727509|0
M1161|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|112|Green||2016-11-07|2016-11-15|NaT||||3.7||3|3|1|1|F|Black||12|Yes|Mother|28227|6|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||24|28209|Bachelors Degree|Single|Business: Sales|28208|0|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|502347820|502348258|31|0|2|504547241|1|0|2|500925514|10|2|-2||2|1|500000294|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||8758769076374727509|0
M1162|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|650|Red||2013-12-18|2014-01-08|2015-10-20|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||21.4||1|1|1|1|F|Black||12|No|Mother|28208|3|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|Black||46|28227|Masters Degree|Married|Finance|28202|8|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503689205|503691170|31|0|2|503689218|31|0|2|500739856|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||7089569121628268952|0
M1163|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|441|Green|PERL 2014-2016, Cabarrus County|2015-12-04|2015-12-22|NaT||||14.5||1|1|2|2|M|White||12|No|Mother|28027|5|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||58|28075|Masters Degree|Married|Business|32824|0|6|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504530586|504532918|1|0|1|503694720|1|0|1|500865400|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|3|||7464|9|||1|500014681, 500016374|3232906304025417619|0
M1164|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|1|1|M|Black||12|No|Mother|28216|6|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|M|Black||39|28278||Married|Business|28202|1|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861229|504863748|31|0|1|504798600|31|0|1|500911906|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1165|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|393|Green||2014-01-15|2014-01-30|2015-02-27|Child: Graduated|Child: Graduated||12.9||1|1|1|1|F|Black||12|No|Mother|28203|3|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|Match Support|F|White||52|28211||Married|Homemaker||0|0|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500008321|503770372|503772348|31|0|2|503594093|1|0|2|500742898|10|1|-1||4|1|500000294|-1||-1|0|4|||7464|9|||1||8568001799025358453|0
M1166|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2017-01-30|2017-01-30|NaT||||1.2||1|1|4|4|M|Black||12|No|Mother|28134|5|One Parent: Female|$50,000 to $59,999|||Y|Yes||Self|General Community||Match Support|M|Black||43|28173|Masters Degree|Married|Finance: Banking|28281|7|0|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504675071|504677498|31|0|1|500353496|31|0|1|500942748|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1||3539543368195872575|3894730386800788938
M1167|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1392|Green|Cabarrus County|2013-04-01|2013-05-15|NaT||||45.7||2|2|1|1|F|Black||12|Yes|Mother|28052|7|One Parent: Female|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|White||40|28052|Bachelors Degree|Single|Transport: Pilot||1|1|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502391396|502391834|31|0|2|503228398|1|0|2|500690843|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|7581500809034284566|0
M1168|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|199|Green|PERL 2014-2016|2015-02-05|2015-02-17|2015-09-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.5||1|1|1|1|M|Black||12|No|Mother|28216|4|One Parent: Female|$45,000 to $49,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||28|28214|Some College|Single|Transport: Driver||0|1|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500017732|504065282|504067309|31|0|1|504168627|31|0|1|500812249|10|2|-2||4|1|500014681|-2|500014681|-2|0|4|||46|2|||1|500014681|7659437100141520816|139697663694671798
M1169|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green||2016-11-11|2016-11-28|NaT||||3.3||1|1|1|1|F|White||12|No|Mother|29715|6|One Parent: Female|$50,000 to $59,999||||No||Self|General Site||Match Support|F|White||45|28079|Masters Degree|Single|Business||0|0|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504886567|504889087|1|0|2|504799615|1|0|2|500927136|10|1|500009132|2128233620|2|1||-1||-1|0|10|||18809|8|||1||1174067921639243853|5215706220873550392
M1170|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|1|1|F|Black||12|No|Mother|28208|6|Two Parent|$20,000 to $24,999||||Yes||Relative|General Site||Match Support|F|White||26|28202|Bachelors Degree|Single|Business|28202|0|3|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861191|504863710|31|0|2|504783413|1|0|2|500911907|10|1|500009132|2128207318|2|1||-1||-1|0|3|||7464|9|||1||2611337051335117774|0
M1171|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|562|Green||2014-11-11|2014-11-18|2016-06-02|Child: Changed school/site|Child: Changed school/site||18.5||1|1|1|1|F|Black||12|No|Mother|28212|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020908|504103367|504105401|31|0|2|503907299|1|0|2|500794438|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1172|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|93|Green||2016-11-21|2016-12-04|NaT||||3.1||1|1|2|2|M|Multi-race (Black & Hispanic)||12|No|Mother|29715|6|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|M|White||31|29707|Bachelors Degree|Married|Customer Service||0|0|LPL Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504908795|504911315|38|0|1|504024654|1|0|1|500929984|10|1|500009132|2128233620|2|1||-1|500014681|-1|0|4|||11247|3|||1||1174067921639243853|0
M1173|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green||2016-11-11|2016-11-28|NaT||||3.3||1|1|1|1|F|White||12|No|Father|29715|6|One Parent: Male|$50,000 to $59,999||||No||School|General Site||Match Support|F|White||39|28204|Bachelors Degree|Single|Business|29715|2|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504890014|504892534|1|0|2|504807342|1|0|2|500927125|10|1|500009132|2128233620|2|1||-1||-1|0|4|||7464|9|||1||1174067921639243853|539886077940116151
M1174|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|266|Green|PERL 2014-2016|2014-09-12|2014-09-23|2015-06-16|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||1|1|1|1|M|Black||12||Mother|28205|4|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|M|White||31|28031||Married|Finance|28202|2|5|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|504016998|504019013|31|0|1|503931397|1|0|1|500775710|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1|500014681|7960300212314874874|0
M1175|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|554|Green||2013-11-18|2013-11-20|2015-05-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.2||1|1|1|1|M|Black||12|No|Mother|28203|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Multi-race (Black & White)||28|28262|Bachelors Degree|Living w/ Significant Other|Personal Trainer/Coach|28205|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500008321|503718040|503720007|31|0|1|503449923|36|0|1|500732241|10|1|-1||4|1||-1||-1|0|4|||7496|10|||1||8568001799025358453|0
M1176|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|726|Yellow||2013-09-18|2013-10-24|2015-10-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||23.9||1|1|1|1|F|Black||12|No|Mother|28208|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||27|28205|Bachelors Degree|Single|Business: Clerical|28277|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503492220|503494082|31|0|2|503521240|1|0|2|500711792|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||976372749760822282|7044657180546140448
M1177|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|168|Green||2016-08-23|2016-09-20|NaT||||5.5||1|1|1|1|M|Black||12|No|Mother|28212|4|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|White||28|28205|Bachelors Degree|Married|Business: Sales|28209|0|10|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504260159|504262304|31|0|1|504639152|1|0|1|500904577|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||0|4802885652788112046
M1178|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1182|Red|Cabarrus County|2013-07-26|2013-08-13|2016-11-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||38.8||1|1|2|2|F|Black||12|No|Mother|28025|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|RTBM|F|Black||43|28027|Masters Degree||Education: Teacher|28027|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500022817|503530345|501204816|31|0|2|502460114|31|0|2|500704946|7|2|500016307||4|3|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|2362631343152316267|0
M1179|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|373|Green||2015-03-05|2015-03-16|2016-03-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.3||1|1|1|1|M|Black||12|No|Mother|28211|4|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|Black||27|28215|High School Graduate|Single|Transport: Driver|28202|3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|503312337|503314167|31|0|1|504201470|31|0|1|500817147|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1||2762897743412756173|4253272603994307857
M1180|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|556|Green||2014-11-17|2014-11-24|2016-06-02|Child: Changed school/site|Child: Changed school/site||18.3||1|1|1|1|F|Black||12|No|Mother|28211|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020908|504112178|504114212|31|0|2|503916397|1|0|2|500796522|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1181|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|225|Green||2014-11-03|2014-11-05|2015-06-18|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||7.4||1|1|2|2|M|Black||12|No|Mother|28205|6|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|White||28|28211|Bachelors Degree|Single|Finance: Accountant|28202|2|0|Duke Energy|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|504085860|504087890|31|0|1|503605925|1|0|1|500791101|10|1|500009132|2128173561|4|1||-1||-1|0|4|||16705|3|||1||7960300212314874874|0
M1182|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|1|1|M|Black||12|No|Father|28208|6|Two Parent|Unknown||||Yes||Relative|General Site||Match Support|M|White||27|28203|Juris Doctorate (JD)|Single|Finance|28202|0|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504870329|504872848|31|0|1|504814162|1|0|1|500911913|10|1|500009132|2128207318|2|1||-1||-1|0|3|||12831|3|||1||2611337051335117774|0
M1183|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1091|Green||2014-03-05|2014-03-12|NaT||||35.8||1|1|1|1|M|White||12|No|Mother|28226|5|One Parent: Female|$200,000 or more||||No||Self|General Community||Match Support|M|White||59|28104|Bachelors Degree|Married|Finance||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503703048|503705013|1|0|1|503354824|1|0|1|500753007|10|2|500009594||2|1||-2||-2|0|10|1562|2|7671|13|1561|2|1||7987165241089060600|6156547733130613405
M1184|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|477|Green|PERL 2014-2016|2015-11-05|2015-11-16|NaT||||15.7||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28216|Bachelors Degree|Married|Business|28202|0|10|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504378557|1|0|1|500856483|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|500014681|4952249713946979108|3402014428779854546
M1185|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|86|Red|PERL 2014-2016|2015-06-16|2015-06-29|2015-09-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||2.8||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28031||Single|Service: Restaurant|28078|0|2|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504186384|1|0|1|500830331|10|2|-2||4|3|500014681|-2|500000294, 500014681|-2|0|4|||7464|9|||1|500014681|4952249713946979108|3402014428779854546
M1186|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1003|Red||2012-10-23|2012-10-31|2015-07-31|Volunteer: Time constraint|Volunteer: Time constraint||33||1|1|1|1|M|Black||12|No|Mother|28215|1|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Asian||39|28262|PHD|Married|Business: Mgt, Admin|28202|4|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502875668|502877071|31|0|1|503114677|4|0|1|500649397|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||314687390558932914|8166272525880133677
M1187|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|319|Green||2016-03-29|2016-04-22|NaT||||10.5||1|1|1|1|F|Black||12|No|Mother|28217|4|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||35|28210|Masters Degree|Married|Finance||5|9|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504268884|504271081|31|0|2|504240747|1|0|2|500886770|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1||7987165241089060600|20998188998147742
M1188|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|76|Green||2016-12-01|2016-12-21|NaT||||2.5||1|1|1|1|M|Black||12|No|Mother|28210|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|M|Black||30|28210|Bachelors Degree|Married|Military||1|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504565095|504567429|31|0|1|504860995|31|0|1|500932205|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||421482027904269589|6156547733130613405
M1189|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-04|2016-10-20|NaT||||4.5||1|1|1|1|F|Black||12|No|Mother|28208|6|Two Parent|Less than $10,000||||Yes||School|General Site||Match Support|F|White||22|28202|Bachelors Degree|Single|Finance|28202|0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504878306|504880826|31|0|2|504775341|1|0|2|500912546|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1190|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|536|Green||2014-01-21|2014-01-31|2015-07-21|Volunteer: Moved|Volunteer: Moved||17.6||2|2|2|2|M|Hispanic||12|No|Father|28212||One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|M|Asian||20|28210||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503777913|503779890|3|0|1|503572872|4|0|1|500744046|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1191|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|237|Green||2015-10-09|2015-10-09|2016-06-02|Child: Changed school/site|Child: Changed school/site||7.8||2|2|2|2|M|Hispanic||12|No|Father|28212||One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503777913|503779890|3|0|1|503907463|1|0|1|500846229|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1192|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|394|Yellow||2015-10-04|2015-10-20|2016-11-17|Volunteer: Moved|Volunteer: Moved||12.9||1|1|1|1|M|Black||12|No|Mother|28273|7|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||RTBM|M|Black||29|28273|High School Graduate|Married|Military|28078|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|504290756|504292957|31|0|1|504315689|31|0|1|500844152|7|2|-2||4|2||-2||-2|0|10|||46|2|||1||194235582162093094|2763237020791144915
M1193|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|389|Green||2014-01-14|2014-02-03|2015-02-27|Child: Graduated|Child: Graduated||12.8||2|2|1|1|F|Black||12|No|Mother|28203|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||59|28211|Bachelors Degree|Married|Retired||0|0|Self|Self|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|502559020|502559473|31|0|2|503590913|1|0|2|500742839|10|1|500000295|2128173558|4|1||-1|500000294|-1|0|4|||7464|9|||1||8568001799025358453|0
M1194|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|945|Green||2013-12-05|2014-01-08|2016-08-10|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||31||1|1|1|1|F|Black||12|No|Mother|28213|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||40|28210|PHD|Single|Medical: Doctor, Provider||0|0|Self|Self|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500016270|503602276|503604153|31|0|2|503381037|31|0|2|500736642|10|1|500000295|2128173561|4|1||-1|500000294|-1|0|4|||7464|9|||1||7960300212314874874|0
M1195|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-10-18|2016-11-17|NaT||||3.6||1|1|2|2|M|Asian||12|No|Mother|28214|6|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site||Match Support|M|Black||48|28205|Masters Degree|Single|Finance|28202|3|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504899975|504902495|4|0|1|504359583|31|0|1|500917107|10|1|500009132|2128207318|2|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1196|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|125|Green||2016-10-19|2016-11-02|NaT||||4.1||1|1|1|1|F|Black||12|Yes|Mother|28208|6|One Parent: Female|Less than $10,000||||Yes||School|General Site|PERL 2014-2016|Match Support|F|White||29|28203|Bachelors Degree|Married|Business|28202|0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861210|504863729|31|0|2|504890087|1|0|2|500917505|10|1|500009132|2128207318|2|1|500014681|-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1197|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|42|Green||2017-01-17|2017-01-24|NaT||||1.4||1|1|2|2|F|Hispanic||12|No|Mother|28212|5|Two Parent|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504998006|505000557|3|0|2|504303308|1|0|2|500940366|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1198|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|161|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-09-27|2016-09-27|NaT||||5.3||2|2|1|1|M|Black||12|No|Mother|28216|3|One Parent: Female|$45,000 to $49,999||||No||Relative|General Community||Match Support|M|Black||37|28269|Bachelors Degree|Single|Business: Engineer||0|9|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|503885975|503887971|31|0|1|504620475|31|0|1|500910396|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|3|||4748|14|||1|500007920, 500011315, 500011316|7702821268191715138|6774573001421433148
M1199|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|444|Red||2014-07-10|2014-08-01|2015-10-19|Volunteer: Moved|Volunteer: Moved||14.6||2|2|1|1|M|Black||12|No|Mother|28216|3|One Parent: Female|$45,000 to $49,999||||No||Relative|General Community||Match Support|M|White||28|28262|Associate Degree|Single|Finance: Banking|28081|1|1|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503885975|503887971|31|0|1|503885544|1|0|1|500769090|10|2|-2||4|3||-2||-2|0|3|||17101|1|||1||7702821268191715138|6774573001421433148
M1200|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|267|Green||2014-09-12|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|1|1|F|Black||12|No|Mother|28269|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Enrollment|F|White||49|28117|Masters Degree|Married|Finance: Banking|28202|5|0|Ally Financial|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|504019066|504021081|31|0|2|503931438|1|0|2|500775724|5|1|500009132|2128173561|4|1||-2||-1|0|4|||12831|3|||1||4952249713946979108|7044657180546140448
M1201|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|324|Red|PERL 2014-2016|2015-02-13|2015-03-09|2016-01-27|Child/Family: Moved|Child/Family: Moved||10.6||1|1|1|1|M|Black||12|No|Mother|29301|5|Two Parent|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28203|Bachelors Degree|Single|Business|28208|0|1|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500013781|504152161|504154211|31|0|1|504180963|1|0|1|500813750|10|2|-2||4|3|500014681|-2|500014681|-2|0|4|||46|2|||1|500014681|0|0
M1202|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|104|Green||2016-11-11|2016-11-23|NaT||||3.4||1|1|3|3|F|Multi-race (Black & White)||12|No|Father|29715|6|Two Parent|$50,000 to $59,999||||No||Self|General Site||Match Support|F|Black||34|28273|Bachelors Degree|Single|Business: Mgt, Admin||5|0|LPL Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504886516|504889036|36|0|2|503255983|31|0|2|500927135|10|1|500009132|2128233620|2|1||-1|500014681|-1|0|10|||11247|3|||1||1174067921639243853|0
M1203|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|454|Yellow||2014-04-10|2014-04-25|2015-07-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.9||2|2|1|1|M|Some Other Race||12||Mother|28277|4|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|White||29|28209|Bachelors Degree|Single|Business|28281|0|1|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|502969243|502970672|41|0|1|503837125|1|0|1|500759182|10|2|-2||4|2||-2||-2|0|10|||132|8|||1||1078778250813636816|0
M1204|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|978|Green||2014-06-25|2014-07-03|NaT||||32.1||1|1|1|1|F|Black||12|No|Mother|28208|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Insurance|28277|0|10|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503739899|503702247|31|0|2|503802084|1|0|2|500767689|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||2611337051335117774|7044657180546140448
M1205|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|298|Green||2014-12-05|2014-12-08|2015-10-02|Child/Family: Moved|Child/Family: Moved||9.8||2|2|1|1|F|Black||12|No|Mother|28083||Other/Unknown|Unknown||||Yes||School|General Site||Match Support|F|Black||37|28025|Associate Degree|Single|Business|28025|12|0|Self|Self|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500012459|503652763|503654723|31|0|2|503985312|31|0|2|500801756|10|1|500000295|2128212919|4|1||-1||-1|0|4|||7464|9|||1||2437132833506538679|0
M1206|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|187|Green||2016-08-30|2016-09-01|NaT||||6.1||1|1|1|1|M|Black||12|No|Mother|28215|4|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28203|Bachelors Degree|Single|Business: Sales|28202|0|3|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504280334|504282534|31|0|1|504556921|1|0|1|500905599|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||18809|8|||1||8998367770661215127|5081726734274569781
M1207|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|676|Green||2013-09-30|2013-09-30|2015-08-07|Volunteer: Moved|Volunteer: Moved||22.2||2|2|1|1|F|Black||12|No|Mother|28211|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503637810|503639770|31|0|2|503603518|1|0|2|500714462|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1208|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|233|Green||2015-10-09|2015-10-13|2016-06-02|Child: Changed school/site|Child: Changed school/site||7.7||2|2|2|2|F|Black||12|No|Mother|28211|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503637810|503639770|31|0|2|503901690|1|0|2|500846292|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1209|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|401|Yellow||2014-04-04|2014-04-22|2015-05-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.2||2|2|1|1|M|Black||12|No|Mother|28212|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||48|28269|Masters Degree|Married|Finance: Banking|28262|9|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503565188|503567063|31|0|1|503814392|31|0|1|500758306|10|2|-2||4|2||-2||-2|0|10|||46|2|||1||0|0
M1210|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|581|Green||2015-06-30|2015-08-04|NaT||||19.1||2|2|1|1|M|Black||12|No|Mother|28212|6|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||27|28211|Bachelors Degree|Married|Finance: Banking|28211|0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503565188|503567063|31|0|1|504265907|1|0|1|500831744|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||0|0
M1211|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|1|1|F|Black||12|No|Mother|28208|6|Two Parent|$25,000 to $29,999||||Yes||School|General Site||Match Support|F|White||27|28202|Bachelors Degree|Single|Finance|28202|0|3|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861159|504863678|31|0|2|504801626|1|0|2|500911905|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1212|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1811|Green||2012-03-09|2012-03-22|NaT||||59.5||2|2|1|1|M|White||12|No|Mother|28277|5|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|White||32|28210|Bachelors Degree|Single|Business: Mgt, Admin|28226|1|5|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502629201|502629856|1|0|1|502893231|1|0|1|500603253|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||3090721985630916616|0
M1213|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-02|2016-10-20|NaT||||4.5||1|1|2|2|F|Black||12|No|Mother|28202|6|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||38|28120|Masters Degree|Divorced|Finance: Accountant|28202|6|4|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504870336|504872855|31|0|2|504348456|1|0|2|500911919|10|1|500009132|2128207318|2|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|241873092051491969
M1214|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1042|Green||2013-07-15|2013-07-19|2016-05-26|Child/Family: Moved|Child/Family: Moved||34.2||1|1|1|1|F|Black||12||Mother|28208|2|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|Black||30|28173|Masters Degree|Single|Education|28262|0|5|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503424337|503426202|31|0|2|503446943|31|0|2|500703604|10|2|-2||4|1||-2||-2|0|5|||7464|9|||1||7581500809034284566|7044657180546140448
M1215|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|289|Green||2014-10-04|2014-10-22|2015-08-07|Volunteer: Moved|Volunteer: Moved||9.5||3|3|2|2|M|White||12|No|Mother|28211|2|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Site||Match Support|M|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503195998|503197751|1|0|1|503507195|1|0|1|500780609|10|1|500000296|2128173564|4|1||-1||-1|6855|8|||0|4|||1||2762897743412756173|0
M1216|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|212|Green||2015-11-03|2015-11-03|2016-06-02|Child: Changed school/site|Child: Changed school/site||7||3|3|3|3|M|White||12|No|Mother|28211|2|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Site||Match Support|M|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503195998|503197751|1|0|1|503905482|1|0|1|500855725|10|1|500000296|2128173564|4|1||-1||-1|6855|8|||0|4|||1||2762897743412756173|0
M1217|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-04|2016-10-20|NaT||||4.5||1|1|2|2|M|Asian||12|No|Mother|28208|6|Two Parent|$15,000 to $19,999||||Yes||School|General Site||Match Support|M|White||25|28210|Bachelors Degree|Single|Finance|28210|0|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504869078|504871597|4|0|1|504359691|1|0|1|500912226|10|1|500009132|2128207318|2|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1218|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1314|Red||2012-02-07|2012-02-10|2015-09-16|Child/Family: Moved|Child/Family: Moved||43.2||1|1|1|1|M|Black||12|No|Mother|28227||One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Multi-race (Hispanic & White)||33|28204|PHD||Medical: Doctor, Provider||0|5|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502290468|502290900|31|0|1|502873884|35|0|1|500596681|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1||0|0
M1219|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|91|Green||2016-11-11|2016-12-06|NaT||||3||1|1|1|1|M|Black||12|No|Mother|28213|5|One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||33|28203|Bachelors Degree|Married|Business|32207|9|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|502383218|502383656|31|0|1|504867282|1|0|1|500926962|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|6854|8|||46|2|||1||0|20998188998147742
M1220|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|650|Green||2013-10-08|2013-10-09|2015-07-21|Volunteer: Moved|Volunteer: Moved||21.4||2|2|1|1|M|Black||12|No|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||20|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503629852|503631791|31|0|1|503613527|31|0|1|500717198|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1221|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|244|Green||2015-10-09|2015-10-13|2016-06-13|Child: Changed school/site|Child: Changed school/site||8||2|2|2|2|M|Black||12|No|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503629852|503631791|31|0|1|503907559|1|0|1|500846287|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1222|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|3|3|M|Black||12|Yes|Mother|28208|6|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|M|Asian||27|28202|Bachelors Degree|Single|Finance|28202|0|1|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861120|504863639|31|0|1|504242094|4|0|1|500911914|10|1|500009132|2128207318|2|1||-1||-1|0|4|||17159|12|||1||2611337051335117774|0
M1223|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2387|Green||2010-08-13|2010-08-24|NaT||||78.4||1|1|1|1|M|Black||12|No|Mother|28216|3|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|White||40|28211|Bachelors Degree|Married|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020753|502222548|502222979|31|0|1|502214317|1|0|1|500465659|10|2|-2||2|1||-2|500000294|-2|0|4|||7496|10|||1||2324686837245224089|0
M1224|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1622|Yellow|Amachi|2011-08-04|2011-08-18|2016-01-26|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||53.3||1|1|1|1|M|Black||12|Yes|Mother|28208|4|One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||42|28212|Masters Degree|Married|Retail: Mgt||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|502367953|502368391|31|0|1|502658210|31|0|1|500548740|10|2|500003586||4|2|500000294|-2||-2|6854|8|||46|2|||1|500000294|4208486535559819469|0
M1225|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|105|Green||2016-11-18|2016-11-22|NaT||||3.4||1|1|2|2|M|Black||12|No|Mother|28212|5|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|White||18|28211||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504932757|504935308|31|0|1|504311367|1|0|1|500929297|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1226|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|103|Green||2016-11-21|2016-11-24|NaT||||3.4||1|1|2|2|M|Hispanic||12|No|Mother|29715|6|Two Parent|$15,000 to $19,999||||No||School|General Site||Match Support|M|White||33|28216|Bachelors Degree|Single|Customer Service||2|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504908812|504911332|3|0|1|504024992|1|0|1|500929993|10|1|500009132|2128233620|2|1||-1||-1|0|4|||11247|3|||1||1174067921639243853|0
M1227|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|135|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-10-16|2016-10-23|NaT||||4.4||1|1|1|1|F|White||12|No|Non-Relative: Other|28205|5|Two Parent|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||25|28207|Bachelors Degree|Single|Tech: Computer/Programmer|28202|1|5|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500021785|504536121|504538455|1|0|2|504562411|1|0|2|500916158|10|2|-2||2|1||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|500007920, 500011315, 500011316|4875067736105190023|2082620892288628337
M1228|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|97|Green||2016-11-09|2016-11-30|NaT||||3.2||1|1|1|1|F|White||12|Yes|Non-Relative: Other|28205|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||28|28202|Bachelors Degree|Single|Finance|28202|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504539986|504538455|1|0|2|504793129|1|0|2|500926111|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||4875067736105190023|2082620892288628337
M1229|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green||2016-11-18|2016-11-28|NaT||||3.3||1|1|1|1|F|Multi-race (Hispanic & White)||12|No|Mother|29715|6|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|Black||50|29708|Bachelors Degree|Widowed|Business||0|5|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504908748|504911268|35|0|2|504821304|31|0|2|500929458|10|1|500009132|2128233620|2|1||-1||-1|0|4|||7464|9|||1||1174067921639243853|3696246430573106858
M1230|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|563|Green||2014-11-11|2014-11-17|2016-06-02|Child: Changed school/site|Child: Changed school/site||18.5||1|1|1|1|F|White||12|No|Mother|28211|4|One Parent: Female|Unknown|||Y|No||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020908|504103364|504105398|1|0|2|503907420|1|0|2|500794450|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1231|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|244|Green||2015-10-13|2015-10-13|2016-06-13|Child: Changed school/site|Child: Changed school/site||8||3|3|2|2|F|Black||12|No|Mother|28211|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28209||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|502776261|502777441|31|0|2|503995722|1|0|2|500847382|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1232|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|655|Green||2013-10-04|2013-10-04|2015-07-21|Volunteer: Moved|Volunteer: Moved||21.5||3|3|1|1|F|Black||12|No|Mother|28211|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28278||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502776261|502777441|31|0|2|503540978|1|0|2|500716168|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1233|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|924|Green|Cabarrus County|2014-08-11|2014-08-26|NaT||||30.4||1|1|1|1|M|White||12|No|Mother|28269|5|One Parent: Female|$60,000 to $74,999||||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|White||35|28075|Masters Degree|Single|Finance: Accountant|28202|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502068488|502068912|1|0|1|503953186|1|0|1|500771917|10|2|500016307||2|1|500016374|-2|500016374|-2|6854|8|||7464|9|||1|500016374|3325175628848876741|5384292856609783094
M1234|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1223|Green||2013-10-31|2013-10-31|NaT||||40.2||1|1|1|1|M|Black||12|No|Mother|28270|2|One Parent: Female|$30,000 to $34,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||32|28210|Bachelors Degree|Single|Tech: Research/Design|28273|0|9|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|503486227|503186577|31|0|1|503555261|31|0|1|500725969|10|2|-2||2|1||-2|500000294|-2|34|2|||46|2|||1||4726905079488957916|663674543177263727
M1235|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|950|Green||2014-07-11|2014-07-31|NaT||||31.2||1|1|1|1|M|Black||12|No|Mother|28214|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||63|28078|Bachelors Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|0|1|277|60|598|500000170|500017732|503810996|503812973|31|0|1|503799211|31|0|1|500769226|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7671|13|||1||7089569121628268952|2763237020791144915
M1236|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-10-02|2016-11-17|NaT||||3.6||1|1|1|1|M|Asian||12|No|Mother|28208|6|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|M|White||47|28216|PHD|Married|Business||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861100|504863619|4|0|1|504798309|1|0|1|500911903|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1237|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|269|Green|Amachi|2015-07-24|2015-08-22|2016-05-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.8||1|1|1|1|F|Black||12|No|Mother|28214|4|One Parent: Female|Unknown|||Y|Yes||School|General Community|Amachi|Match Support|F|Asian||33|28205|Bachelors Degree|Single|Consultant|60654|2|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|504166613|504168697|31|0|2|503823941|4|0|2|500834370|10|2|-2||4|1|500000294|-2||-2|0|4|||7464|9|||1|500000294|7089569121628268952|0
M1238|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|246|Green||2015-01-26|2015-01-29|2015-10-02|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||8.1||1|1|1|1|F|Black||12|Yes|GrandMother|28081|3|Grandparents|Unknown||||Yes||School|General Site||Match Support|F|White||19|28117|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500002335|504106278|504108312|31|0|2|504043172|1|0|2|500810108|10|1|500000296|2128173571|4|1||-1||-1|0|4|||0|4|||1||0|0
M1239|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-11|2016-12-02|NaT||||3.1||1|1|3|3|M|Black||12|Yes|GrandMother|29715|6|Two Parent|Unknown||||No||School|General Site||Match Support|M|Black||31|29710|Bachelors Degree|Married|Consultant|28217|3|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504890029|504892549|31|0|1|504060437|31|0|1|500927118|10|1|500009132|2128233620|2|1||-1||-1|0|4|||11247|3|||1||1174067921639243853|0
M1240|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|300|Green||2014-09-21|2014-09-23|2015-07-20|Volunteer: Moved|Volunteer: Moved||9.9||4|4|2|2|F|White||12|No|Mother|28211|1|Two Parent|Unknown||||No||School|General Site||Match Support|F|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502763403|502764315|1|0|2|503603510|1|0|2|500777105|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1241|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|248|Green||2015-10-09|2015-10-09|2016-06-13|Child: Changed school/site|Child: Changed school/site||8.1||4|4|2|2|F|White||12|No|Mother|28211|1|Two Parent|Unknown||||No||School|General Site||Match Support|F|White||18|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|502763403|502764315|1|0|2|503905493|1|0|2|500846254|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1242|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|981|Green||2014-06-20|2014-06-30|NaT||||32.2||1|1|1|1|M|Black||12|No|GrandMother|28216|3|Grandparents|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||45|28269|Bachelors Degree|Married|Finance: Banking|28273|1|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503866348|503838583|31|0|1|503862591|1|0|1|500767276|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1||7679812394383646966|9060571453147419923
M1243|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1076|Green||2014-03-21|2014-03-27|NaT||||35.4||2|2|1|1|M|Black||12|Yes|Mother|28205||One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||27|28202|Bachelors Degree|Single|Business|28217|0|8|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502162237|503458866|31|0|1|503151333|1|0|1|500756070|10|2|-2||2|1|500000294|-2||-2|6854|8|||7464|9|||1||0|4899444095790462270
M1244|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|613|Green||2013-11-10|2013-11-14|2015-07-20|Volunteer: Moved|Volunteer: Moved||20.1||2|2|1|1|F|Black||12|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503707963|503709929|31|0|2|503507325|1|0|2|500729570|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1245|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|232|Green||2015-10-09|2015-10-21|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.6||2|2|2|2|F|Black||12|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||18|28227|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503707963|503709929|31|0|2|504302535|31|0|2|500846355|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1246|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|393|Green||2014-01-15|2014-01-30|2015-02-27|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||12.9||1|1|1|1|F|Black||12|No|Father|28202|3|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|F|White||83|28226|Masters Degree|Widowed|Retired||0|0|Self|Self|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|503770356|503772332|31|0|2|503479599|1|0|2|500742899|10|1|-1||4|1||-1|500000294|-1|0|4|||7464|9|||1||8568001799025358453|0
M1247|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|281|Green||2014-10-17|2014-10-30|2015-08-07|Volunteer: Moved|Volunteer: Moved||9.2||1|1|2|2|M|Hispanic||12|No|Mother|28212|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|M|Asian||19|28211|Some High School|Single|Student: College||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504070362|504072390|3|0|1|503507276|4|0|1|500784776|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1248|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|346|Red||2015-03-09|2015-03-30|2016-03-10|Child/Family: Moved|Child/Family: Moved||11.4||1|1|1|1|M|Hispanic||12|No|Mother|28217||One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Hispanic||32|28203|Bachelors Degree|Single|Business: Sales|28203|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500020753|504234460|504236575|3|0|1|503812408|3|0|1|500817510|10|1|500000295|2128173557|4|3||-1||-1|0|4|||7496|10|||1||8981704271528751143|0
M1249|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|3|3|M|Hispanic||12|No|Mother|28208|6|Two Parent|$20,000 to $24,999||||Yes||School|General Site||Match Support|M|White||24|29708|Bachelors Degree|Single|Finance|28202|0|10|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504875023|504877543|3|0|1|504475369|1|0|1|500911912|10|1|500009132|2128207318|2|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1250|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|382|Red|PERL 2014-2016, Cabarrus County|2016-02-02|2016-02-19|NaT||||12.6||1|1|2|2|F|Black||12|No|Mother|28083|5|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||41|28025|Some College|Single|Business|28217|4|0|LPL Financial|Workplace Partner|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504540553|504805582|31|0|2|503680923|31|0|2|500877015|10|2|500016307||2|3|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||11247|3|||1|500014681, 500016374|2437132833506538679|0
M1251|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|640|Green||2013-11-01|2013-11-05|2015-08-07|Volunteer: Moved|Volunteer: Moved||21||2|2|2|2|F|Black||12|Yes|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503670769|503672730|31|0|2|503493268|1|0|2|500726477|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1252|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|244|Green||2015-10-09|2015-10-13|2016-06-13|Child: Changed school/site|Child: Changed school/site||8||2|2|2|2|F|Black||12|Yes|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503670769|503672730|31|0|2|503905510|1|0|2|500846278|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1253|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|589|Green||2015-07-16|2015-07-27|NaT||||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|||Y|Yes||Relative|General Community||Match Support|F|White||29|28209|Bachelors Degree|Single|Retail: Mgt|28217|3|3|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504312629|504314787|31|0|2|504262612|1|0|2|500833665|10|2|-2||2|1||-2||-2|0|3|||17159|12|||1||0|237874676114443178
M1254|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|589|Green|PERL 2014-2016|2015-07-20|2015-07-27|NaT||||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Asian||28|28203|Bachelors Degree|Single|Consultant|28202|1|1|Current/Previous Big|Other Big|Big|General Community|mentor2.0, mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500008321|504312569|504314787|31|0|2|504208036|4|0|2|500833808|10|2|-2||2|1|500014681|-2|500014505, 500015184|-2|0|4|||17159|12|||1|500014681|0|237874676114443178
M1255|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|921|Yellow||2014-08-15|2014-08-29|NaT||||30.3||1|1|1|1|F|Black||12|Yes|Mother|28208|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||28|28205|Masters Degree|Single|Business: Mgt, Admin|28262|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503941222|503931754|31|0|2|503889588|1|0|2|500772492|10|2|-2||2|2||-2||-2|0|4|||17159|12|||1||5424205421938369753|0
M1256|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|700|Red||2014-08-15|2014-08-29|2016-07-29|Volunteer: Time constraint|Volunteer: Time constraint||23||1|1|1|1|F|Black||12|Yes|Mother|28208|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Multi-race (Asian & White)||27|28203|Bachelors Degree|Single|Finance|28211|0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503929747|503931754|31|0|2|503910740|37|0|2|500772491|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1||5424205421938369753|0
M1257|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|230|Green||2014-10-04|2014-10-17|2015-06-04|Volunteer: Moved|Volunteer: Moved||7.6||3|3|2|2|M|Black||12|No|Mother|28211|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||20|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503644180|503646140|31|0|1|503493918|1|0|1|500780600|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1258|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|503|Green||2015-10-09|2015-10-21|NaT||||16.5||3|3|1|1|M|Black||12|No|Mother|28211|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||18|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|503644180|503646140|31|0|1|504327166|31|0|1|500846331|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1259|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1173|Green||2013-12-05|2013-12-20|NaT||||38.5||1|1|1|1|F|Black||12|No|Mother|28215|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||23|28227||Single|Student: College|28202|2|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503638969|503640929|31|0|2|503503174|31|0|2|500736646|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||3723482195151978288|0
M1260|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|319|Green||2014-09-21|2014-09-22|2015-08-07|Volunteer: Moved|Volunteer: Moved||10.5||3|3|2|2|F|Hispanic||12|No|Mother|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503391535|503393392|3|0|2|503497423|1|0|2|500777106|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1261|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|16|Green||2015-11-02|2015-11-03|2015-11-19|Child/Family: Moved|Child/Family: Moved||0.5||3|3|3|3|F|Hispanic||12|No|Mother|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28207|Some College|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503391535|503393392|3|0|2|504306107|1|0|2|500855267|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1262|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1822|Green||2011-08-16|2011-08-31|2016-08-26|Child/Family: Moved|Child/Family: Moved||59.9||1|1|1|1|M|Black||12|No|Mother|28208|K|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||35|28207|Masters Degree|Married|Law: Lawyer|28202|8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|1|0|1|0|277|60|598|500000170|500020910|502431040|502431483|31|0|1|502609637|1|0|1|500550314|10|2|-2||4|1||-2|500004640|-2|0|10|||7496|10|||1||5533634913091743658|0
M1263|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|1312|Green||2012-12-13|2012-12-17|2016-07-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||43.1||2|2|2|2|M|Black||12|Yes|Mother|28205|5|One Parent: Female|Unknown||||Yes||School|General Site|Project Big AND Amachi|Match Support|M|Black||31|28273||Single|Tech: Support, Writing||0|0|Omega Psi Phi|Fraternity/Sorority|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|502766031|502766944|31|0|1|501946079|31|0|1|500669679|10|1|500000295|2128173561|4|1|500004901|-1||-1|0|4|||8694|14|||1||7960300212314874874|0
M1264|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|122|Green|PERL 2014-2016|2015-08-10|2015-08-30|2015-12-30|Child/Family: Moved|Child/Family: Moved||4||1|1|1|1|F|Black||12|No|Mother|28212|4|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||33|28270|Some College|Single|Business|28262|1|3|Other|BBBS Board/Staff|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500017732|504343306|504345530|31|0|2|504109000|31|0|2|500835668|10|2|-2||4|1|500014681|-2||-2|0|10|||7671|13|||1|500014681|7554307376683929204|2876415545463317777
M1265|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1088|Green||2014-03-05|2014-03-15|NaT||||35.7||1|1|1|1|M|Black||12|Yes|Mother|28216|3|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||49|28204|Bachelors Degree|Married|Finance: Accountant|28255|8|0|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020910|503565637|503567522|31|0|1|503604089|1|0|1|500752839|10|2|-2||2|1|500000294|-2|500000294, 500014681|-2|34|2|||7464|9|||1||2979941694006626856|1786514887916898235
M1266|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|609|Green||2014-10-04|2014-10-07|2016-06-07|Volunteer: Moved|Volunteer: Moved||20||1|1|1|1|M|Black||12|No|Mother|28105|3|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|RTBM|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020909|504049262|504051286|31|0|1|503907248|1|0|1|500780579|7|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1267|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|106|Green||2016-11-11|2016-11-21|NaT||||3.5||1|1|2|3|F|Multi-race (Black & White)||11|No|Mother|29715|6|One Parent: Female|$30,000 to $34,999||||No||School|General Site||Match Support|F|Black||53|28226|Bachelors Degree|Single|Business: Mgt, Admin|28217|2|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504890059|504892579|36|0|2|504394474|31|0|2|500927142|10|1|500009132|2128233620|2|1||-1||-1|0|4|||11247|3|||1||1174067921639243853|3166474625198890934
M1268|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-11|2016-11-17|NaT||||3.6||1|1|2|2|F|Black||11|No|GrandMother|28269|6|Grandparents|Less than $10,000||||Yes||School|General Site||Match Support|F|White||35|28226|Bachelors Degree|Married|Finance|28202|0|1|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500021785|504878293|504880813|31|0|2|504632567|1|0|2|500927086|10|1|500009132|2128207318|2|1||-1|500007920, 500011315, 500011316, 500014681|-1|0|4|||12831|3|||1||2611337051335117774|0
M1269|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|302|Green||2014-09-21|2014-09-22|2015-07-21|Volunteer: Moved|Volunteer: Moved||9.9||3|3|2|2|F|Black||11||Father|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503196044|502747550|31|0|2|503509836|31|0|2|500777107|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1270|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|247|Green||2015-10-06|2015-10-06|2016-06-09|Child: Changed school/site|Child: Changed school/site||8.1||3|3|2|2|F|Black||11||Father|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||18|28213|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503196044|502747550|31|0|2|504324154|31|0|2|500844552|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1271|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|301|Green||2014-09-21|2014-09-23|2015-07-21|Volunteer: Moved|Volunteer: Moved||9.9||4|4|2|2|M|Black||11|No|Father|28212||One Parent: Male|Unknown||||No||School|General Site||Match Support|M|Black||20|28277||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502746641|502747550|31|0|1|503540909|31|0|1|500777109|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1272|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|248|Green||2015-10-09|2015-10-09|2016-06-13|Child: Changed school/site|Child: Changed school/site||8.1||4|4|2|2|M|Black||11|No|Father|28212||One Parent: Male|Unknown||||No||School|General Site||Match Support|M|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|502746641|502747550|31|0|1|503907262|1|0|1|500846196|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1273|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|222|Green||2016-06-28|2016-07-28|NaT||||7.3||1|1|1|1|F|Black||11|No|Mother|28215|6|One Parent: Female|$30,000 to $34,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||30|28209|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28204|2|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504671571|504673998|31|0|2|504308223|1|0|2|500898271|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1||7284449467126735125|20998188998147742
M1274|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|106|Green||2016-11-11|2016-11-21|NaT||||3.5||1|1|1|1|F|White||11|No|Mother|29715|6|One Parent: Female|$20,000 to $24,999||||No||School|General Site||Match Support|F|White||50|29710|Bachelors Degree|Married|Business||3|0|Self|Self|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500013781|504890041|504892561|1|0|2|504817368|1|0|2|500927127|10|1|500009132|2128233620|2|1||-1|500007920, 500011315, 500011316|-1|0|4|||7464|9|||1||1174067921639243853|3979721973761636002
M1275|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-04|2016-10-20|NaT||||4.5||1|1|2|2|F|Black||11|No|Mother|28208|6|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||33|28209|Bachelors Degree|Single|Finance|28202|4|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861049|504863568|31|0|2|504354941|1|0|2|500912228|10|1|500009132|2128207318|2|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|7088853613314985400
M1276|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|990|Red||2012-11-20|2012-12-01|2015-08-18|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||32.5||1|1|1|1|M|Black||11|No|Mother|28278|0|One Parent: Female|$35,000 to $39,999||||No||Self|General Community||Match Support|M|White||34|29708|High School Graduate|Single|Business: Mgt, Admin|29730|11|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502527969|502528422|31|0|1|503169378|1|0|1|500662254|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||0|0
M1277|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|196|Green||2014-09-15|2014-12-03|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||6.4||1|1|1|1|M|Black||11|No|Father|28206|5|One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|M|White||28|28211|Bachelors Degree|Single|Finance: Banking|28202|8|0|Ally Financial|Workplace Partner|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503996753|503998768|31|0|1|503911411|1|0|1|500775988|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M1278|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|281|Green||2014-10-04|2014-10-30|2015-08-07|Volunteer: Moved|Volunteer: Moved||9.2||2|2|2|2|F|Black||11|No|Father|28105|4|One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049370|504051394|31|0|2|503517772|1|0|2|500780607|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1279|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|232|Green||2015-10-09|2015-10-21|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.6||2|2|2|2|F|Black||11|No|Father|28105|4|One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||17|28269|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504049370|504051394|31|0|2|504301152|31|0|2|500846352|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1280|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1453|Green||2013-03-12|2013-03-15|NaT||||47.7||1|1|1|1|F|Black||11|No|Mother|28212|4|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Finance|28202|0|4|Relative|Relative|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503259350|503261158|31|0|2|503370160|1|0|2|500687348|10|2|-2||2|1||-2||-2|34|2|||17161|11|||1||7554307376683929204|7044657180546140448
M1281|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|93|Green||2016-11-18|2016-12-04|NaT||||3.1||1|1|1|1|F|Black||11|Yes|Mother|29715|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||36|28277|Juris Doctorate (JD)|Married|Business|29715|1|3|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504908826|504911346|31|0|2|504829966|1|0|2|500929469|10|1|500009132|2128233620|2|1||-1||-1|0|4|||7464|9|||1||1174067921639243853|0
M1282|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|316|Green||2016-04-08|2016-04-25|NaT||||10.4||1|1|1|1|M|White||11|No|Mother|28277|5|One Parent: Female|$60,000 to $74,999||||No||School|General Community||Match Support|M|White||40|28173|Bachelors Degree|Married|Business: Mgt, Admin|33637|9|4|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504240231|504242346|1|0|1|504523981|1|0|1|500888425|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||3090721985630916616|7406803744350640674
M1283|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|676|Green||2013-09-30|2013-09-30|2015-08-07|Volunteer: Moved|Volunteer: Moved||22.2||3|3|1|1|F|Hispanic||11|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503204695|503206461|3|0|2|503506209|1|0|2|500714422|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1284|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|489|Green||2015-10-16|2015-11-04|NaT||||16.1||3|3|1|1|F|Hispanic||11|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|503204695|503206461|3|0|2|504301092|1|0|2|500848809|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1285|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|43|Green||2017-01-06|2017-01-23|NaT||||1.4||2|2|1|1|M|Black||11|No|Mother|28205|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||24|28202|Bachelors Degree|Single|Construction|28217|0|9|BBBS National Site|Web Link|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500015820|503779546|503781523|31|0|1|504625641|1|0|1|500938754|10|1|500000295|2128207319|2|1||-1|500007920, 500011315, 500011316|-1|0|4|||46|2|||1||3935539763241716148|8561594548502006295
M1286|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|204|Green||2015-03-12|2015-03-12|2015-10-02|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.7||2|2|1|1|F|Black||11||Relative: Other|28026||One Parent: Female|Unknown|||Y|Yes||Therapist/Counselor|General Site||Enrollment|F|White||18|28083||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500002335|503669127|503671088|31|0|2|504220439|1|0|2|500818544|5|1|500000296|2128173571|4|1||-1||-1|0|5|||0|4|||1||1550830965009450729|0
M1287|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|116|Green||2016-10-03|2016-11-11|NaT||||3.8||1|1|3|3|M|Black||11|No|Father|28208|6|One Parent: Male|$20,000 to $24,999||||Yes||School|General Site||Match Support|M|White||30|28273|Bachelors Degree|Single|Finance|28202|1|8|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504870344|504872863|31|0|1|503911379|1|0|1|500911991|10|1|500009132|2128207318|2|1||-1||-1|0|4|||12831|3|||1||2611337051335117774|0
M1288|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|137|Green||2016-10-04|2016-10-21|NaT||||4.5||1|1|3|3|M|Black||11|No|Mother|28208|6|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site||Match Support|M|Black||25|28269|Masters Degree|Single|Finance|28202|0|1|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504870349|504872868|31|0|1|504359606|31|0|1|500912557|10|1|500009132|2128207318|2|1||-1|500014681|-1|0|4|||12831|3|||1||2611337051335117774|0
M1289|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|1|1|M|Black||11|No|Mother|28208|6|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site||Match Support|M|Black||29|28027|Bachelors Degree|Married|Business||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504870355|504872868|31|0|1|504798428|31|0|1|500911916|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1290|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|227|Red||2016-02-11|2016-03-14|2016-10-27|Child/Family: Moved|Child/Family: Moved||7.5||2|2|1|1|F|Hispanic||11|No|Mother|28217|3|One Parent: Female|Unknown|||Y|Yes||School|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||32|28277|Bachelors Degree|Single|Business: Sales|28277|1|3|Neighbor/Friend|Neighbor/Friend|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500013781|503779482|503781459|3|0|2|504510616|31|0|2|500879051|10|1|500000295|2128173557|4|3|500007920, 500011315, 500011316|-1|500007920, 500011315, 500011316|-1|0|4|||7496|10|||1||8981704271528751143|0
M1291|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|670|Red|VOL - Mentoring Hispanic Youth|2014-01-17|2014-02-19|2015-12-21|Volunteer: Time constraint|Volunteer: Time constraint||22||2|2|1|1|F|Hispanic||11|No|Mother|28217|3|One Parent: Female|Unknown|||Y|Yes||School|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||27|28262|Bachelors Degree|Single|Student: College||0|9|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020753|503779482|503781459|3|0|2|503108667|31|0|2|500743569|10|1|500000295|2128173557|4|3|500007920, 500011315, 500011316|-1||-1|0|4|||7464|9|||1|500011312|8981704271528751143|0
M1292|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|667|Green||2013-10-08|2013-10-09|2015-08-07|Volunteer: Moved|Volunteer: Moved||21.9||3|3|1|1|F|Hispanic||11|No|Father|28212|1|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502763413|502764325|3|0|2|503577783|1|0|2|500717205|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1293|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|244|Green||2015-10-13|2015-10-13|2016-06-13|Child: Changed school/site|Child: Changed school/site||8||3|3|2|2|F|Hispanic||11|No|Father|28212|1|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|502763413|502764325|3|0|2|503907351|1|0|2|500847613|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1294|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|81|Green||2016-12-16|2016-12-16|NaT||||2.7||1|1|1|1|F|White||11|No|Mother|29715|6|Two Parent|$50,000 to $59,999||||No||School|General Site||Match Support|F|Black||35|28216|Bachelors Degree|Single|Business||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504960112|504962663|1|0|2|504789046|31|0|2|500936175|10|1|500009132|2128233620|2|1||-1||-1|0|4|||7464|9|||1||1174067921639243853|0
M1295|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|376|Green||2014-09-12|2014-09-24|2015-10-05|Child: Changed school/site|Child: Changed school/site||12.4||1|1|1|1|F|Black||11|Yes|Mother|28216|5|One Parent: Female|Unknown||||No||School|General Site||Match Support|F|Black||39|28269||Single|Finance|28202|2|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504013280|504015295|31|0|2|503908838|31|0|2|500775717|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M1296|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|258|Yellow||2016-02-18|2016-02-26|2016-11-10|Child: Graduated|Child: Graduated||8.5||1|1|1|1|F|Black||11|No|Mother|28027|5|Two Parent|Less than $10,000|||Y|Yes||School|General Site|Cabarrus County|Match Support|F|White||18|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504629037|504631448|31|0|2|504619538|1|0|2|500880057|10|1|500000296|2128173571|4|2|500016374|-1|500016374|-1|0|4|||7464|9|||1||3232906304025417619|0
M1297|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|658|Green||2014-06-18|2014-06-30|2016-04-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.6||1|1|1|1|M|Black||11|No|Mother|28216|5|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Enrollment|M|White||31|28210|Masters Degree|Single|Finance|28211|8|1|Recruitment Event|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503686272|503688237|31|0|1|503817633|1|0|1|500766948|5|2|-2||4|1||-2||-2|0|10|||7460|12|||1||5367149751093883357|0
M1298|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1077|Green||2014-03-04|2014-03-26|NaT||||35.4||1|1|1|1|F|Black||11|No|Mother|28216|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|Black||42|28273|Bachelors Degree|Single|Customer Service|28273|4|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503691322|503688237|31|0|2|503763297|31|0|2|500752718|10|2|-2||2|1||-2||-2|0|5|||7464|9|||1||7473714268566895255|0
M1299|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|224|Green||2015-01-22|2015-03-09|2015-10-19|Child/Family: Moved|Child/Family: Moved||7.4||1|1|2|2|M|Black||11|No|Mother|28217|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||28|28207|Bachelors Degree|Single|Finance|28277|1|6|Self|Self|Big|General Site||Enrollment|0|1|1|0|277|60|598|500000170|500020753|504184668|504186777|31|0|1|503338695|1|0|1|500809563|10|1|500000295|2128173557|4|1||-1||-1|0|4|||7464|9|||1||8981704271528751143|0
M1300|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1572|Green||2012-10-23|2012-11-16|NaT||||51.6||1|1|1|1|F|Black||11|No|Mother|28210|2|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||28|28226|Bachelors Degree|Single|Education: Teacher|28173|2|6|TV|Media|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|503143377|503145049|31|0|2|503109316|1|0|2|500649731|10|2|-2||2|1||-2|500000294|-2|0|10|||130|1|||1||4902029756574603597|2940594469294202107
M1301|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|231|Green||2014-10-04|2014-10-17|2015-06-05|Volunteer: Moved|Volunteer: Moved||7.6||3|3|2|2|F|Black||11|No|Mother|28212|2|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503196065|504449560|31|0|2|503497346|1|0|2|500780605|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1302|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|251|Green||2015-10-06|2015-10-06|2016-06-13|Child: Changed school/site|Child: Changed school/site||8.2||3|3|2|2|F|Black||11|No|Mother|28212|2|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503196065|504449560|31|0|2|504308470|1|0|2|500844551|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1303|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|498|Green||2013-12-09|2013-12-17|2015-04-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.4||1|1|1|1|F|Black||11|No|Mother|28217|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||31|28273|Masters Degree|Single|Customer Service|28025|0|6|AA Task Force|Other Big|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016847|503745285|503747257|31|0|2|503655183|31|0|2|500737658|10|1|500000295|2128173557|4|1||-1||-1|0|4|||6247|12|||1||8981704271528751143|0
M1304|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1301|Green||2013-08-02|2013-08-14|NaT||||42.7||1|1|1|1|M|Black||11|No|Mother|28215|1|One Parent: Female|$35,000 to $39,999||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||41|28211|Bachelors Degree|Single|Finance: Banking|28209|5|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|502934728|502936151|31|0|1|503516330|31|0|1|500705674|10|2|-2||2|1||-2|500000294|-2|6854|8|||7464|9|||1||4575902950186762737|0
M1305|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green||2016-11-11|2016-11-28|NaT||||3.3||1|1|1|1|F|White||11|No|GrandMother|29715|6|Grandparents|$20,000 to $24,999||||Yes||Self|General Site||Match Support|F|Black||28|29715|Bachelors Degree|Single|Business|29715|0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504886538|504889058|1|0|2|504829898|31|0|2|500927102|10|1|500009132|2128233620|2|1||-1||-1|0|10|||7464|9|||1||1174067921639243853|0
M1306|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1019|Green||2014-05-07|2014-05-23|NaT||||33.5||2|2|1|1|M|Black||11|No|GrandMother|28210|3|Grandparents|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||34|28210|Masters Degree|Married|Finance: Banking|28202|8|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503609425|503611302|31|0|1|503837417|1|0|1|500762429|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||5711791743715234276|1786514887916898235
M1307|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|389|Green|PERL 2014-2016|2016-01-29|2016-02-12|NaT||||12.8||1|1|1|1|M|Black||11|Yes|Mother|28215|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||29|28262|Some College|Single|Business|28204|0|4|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT, VOL - Thrive - Intro|Match Support|0|1|0|1|277|60|598|500000170|500020753|504230975|504233090|31|0|1|504284612|31|0|1|500876290|10|2|-2||2|1|500000294, 500014681|-2|500008492, 500011315, 500011316, 500014681|-2|0|4|||7462|13|||1|500014681|6077912216232501082|7327400833679234452
M1308|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|415|Red||2014-10-01|2014-10-13|2015-12-02|Volunteer: Time constraint|Volunteer: Time constraint||13.6||1|1|1|1|M|Black||11|Yes|Mother|28215|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Enrollment|M|Black||26|28227|Bachelors Degree|Single|Customer Service||1|3|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503723888|503725860|31|0|1|503858682|31|0|1|500779634|5|2|-2||4|3||-2||-2|0|10|||17101|1|||1||5741767063897867874|8861046674172959830
M1309|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|945|Green||2014-07-14|2014-08-05|NaT||||31||1|1|1|1|F|Black||11|No|Mother|28216|5|One Parent: Female|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Some Other Race||30|28214|Bachelors Degree|Married|Business|28214|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502602926|502603443|31|0|2|503808719|41|0|2|500769460|10|2|-2||2|1||-2||-2|6854|8|||7462|13|||1||2456895876914964961|20998188998147742
M1310|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|116|Green||2016-10-02|2016-11-11|NaT||||3.8||1|1|1|1|F|Black||11|No|Mother|28214|6|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||29|28202|Bachelors Degree|Married|Business: Mgt, Admin|28202|0|3|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861132|504863651|31|0|2|504771994|1|0|2|500911917|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|3200475665780018500
M1311|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|600|Green||2013-11-25|2013-12-19|2015-08-11|Child: Changed school/site|Child: Changed school/site||19.7||1|1|1|1|M|Black||11|No|Mother|28205|2|One Parent: Female|Unknown||||No||School|General Site||Match Support|M|Black||40|28203||Single|Business: Engineer|28244|6|7|Recruitment Event|Self|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503217239|503219020|31|0|1|503666439|31|0|1|500734576|10|1|500000295|2128173561|4|1||-1||-1|0|4|||7458|9|||1||7960300212314874874|0
M1312|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|748|Yellow||2013-07-11|2013-07-30|2015-08-17|Child: Family structure changed|Child: Family structure changed||24.6||1|1|1|1|M|Black||11|Yes|GrandMother|28273|3|Foster Home|$25,000 to $29,999|||Y|Yes||Self|General Community|Amachi|Enrollment|M|White||32|28209|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|5|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500015820|502299232|501806520|31|0|1|503510609|1|0|1|500703319|5|2|-2||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1||0|0
M1313|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2004|Green||2011-08-29|2011-09-11|NaT||||65.8||1|1|2|2|F|Black||11|No|Mother|28205|1|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|White||32|28134|Bachelors Degree|Single|Finance: Banking|28288|0|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502653228|502653964|31|0|2|502192090|1|0|2|500552244|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||6627885846854295604|1018920374251832097
M1314|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|137|Green||2016-10-08|2016-10-21|NaT||||4.5||1|1|1|1|F|Black||11|No|Mother|28208|6|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||25|28202|Bachelors Degree|Single|Business: Mgt, Admin|28202|1|2|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861085|504863604|31|0|2|504391145|1|0|2|500913788|10|1|500009132|2128207318|2|1||-1||-1|0|4|||46|2|||1||2611337051335117774|4554908796282949108
M1315|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-03|2016-10-20|NaT||||4.5||1|1|2|2|F|Black||11|No|Mother|28208|6|One Parent: Female|$10,000 to $14,999||||Yes||Self|General Site||Match Support|F|Black||31|28277|Associate Degree|Single|Finance: Auditor|28202|0|3|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500021785|504870325|504872844|31|0|2|504349862|31|0|2|500912043|10|1|500009132|2128207318|2|1||-1|500014681|-1|0|10|||12831|3|||1||2611337051335117774|0
M1316|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|610|Green||2014-10-04|2014-10-07|2016-06-08|Volunteer: Moved|Volunteer: Moved||20||1|1|1|1|F|Hispanic||11|Yes|Mother|28212|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||19|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504041972|504043990|3|0|2|503897715|1|0|2|500780591|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1317|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|771|Green||2015-01-14|2015-01-26|NaT||||25.3||3|3|2|2|F|Black||11|No|Mother|28216|2|One Parent: Female|Unknown||||Yes|TV|Media|General Community||Match Support|F|Black||48|28203|Bachelors Degree|Married|Business: Mgt, Admin|28202|1|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502324604|502325039|31|0|2|502657850|31|0|2|500808029|10|2|-2||2|1||-2||-2|56|1|||7464|9|||1||7679812394383646966|0
M1318|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1936|Yellow||2010-12-29|2011-01-14|2016-05-03|Volunteer: Time constraint|Volunteer: Time constraint||63.6||1|1|1|1|M|Black||11|No|Mother|28227|4|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|Some Other Race||38|28209|Bachelors Degree|Single|Business: Mgt, Admin|28205|5|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502211032|502211462|31|0|1|502276859|41|0|1|500508474|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1||6505995099520362521|1937926248155442003
M1319|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|237|Red||2014-05-28|2014-06-13|2015-02-05|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.8||1|1|1|1|M|Black||11|No|Mother|28216|3|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||62|28210|Bachelors Degree|Divorced|Business: Engineer|28202|35|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503492511|503494379|31|0|1|503852376|1|0|1|500764721|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1||2456895876914964961|0
M1320|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|266|Green|Cabarrus County|2016-06-14|2016-06-14|NaT||||8.7||1|1|1|1|F|White||11|No|GrandMother|28124|5|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community|Cabarrus County|Match Support|F|White||45|28025|Some College||Business|28262|1|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504635786|504638197|1|0|2|504662207|1|0|2|500896660|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|1345826867198613426|0
M1321|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|214|Green|Cabarrus County|2016-08-01|2016-08-05|NaT||||7||1|1|1|1|F|Black||11|No|Mother|28027|4|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||35|28027|Masters Degree|Married|Medical: Nurse||0|6|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504026659|504028677|31|0|2|504744796|31|0|2|500901331|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|3|||7464|9|||1|500016374|6810228174639243761|0
M1322|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2199|Green||2011-02-18|2011-02-28|NaT||||72.2||1|1|1|1|F|Black||11|No|Mother|28216||One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||29|28207|Bachelors Degree|Single|Human Services: Non-Profit|28212|1|4|Newspaper|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|502274606|502275038|31|0|2|502441954|1|0|2|500518627|10|2|-2||2|1||-2||-2|6854|8|||129|1|||1||0|0
M1323|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|527|Green|PERL 2014-2016|2015-01-13|2015-02-10|2016-07-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||17.3||1|1|2|2|F|Black||11|No|Mother|28206|4|One Parent: Female|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|Hispanic||36|28210|Bachelors Degree|Married|Finance: Accountant|28203|4|0|BBBS National Site|Web Link|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|504100771|504102805|31|0|2|504000676|3|0|2|500807798|10|1|500000295|2128173561|4|1|500014681|-1|500014681|-1|0|4|||46|2|||1|500014681|7960300212314874874|0
M1324|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|149|Green|PERL 2014-2016|2014-12-09|2014-12-16|2015-05-14|Child/Family: Time constraints|Child/Family: Time constraints||4.9||2|2|2|2|M|Black||11|No|GrandMother|28270|3|Grandparents|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|M|White||57|28105|Bachelors Degree|Married|Business: Sales|28203|11|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500018987|503650948|503652908|31|0|1|504063702|1|0|1|500802395|5|2|-2||4|1|500014681|-2|500000294|-2|0|10|||17159|12|||1|500014681|4726905079488957916|0
M1325|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|165|Green||2016-09-23|2016-09-23|NaT||||5.4||1|1|1|1|F|Black||11|No|Mother|28212|5|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||37|28227|Bachelors Degree|Married|Business: Mgt, Admin|28173|10|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504357732|504359958|31|0|2|504576046|1|0|2|500909829|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1||4487969519148815281|6692528426538080183
M1326|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|642|Green||2013-10-15|2013-10-17|2015-07-21|Volunteer: Moved|Volunteer: Moved||21.1||2|2|1|1|F|Black||11|No|Relative: Other|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28207||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503644199|503646159|31|0|2|503540939|1|0|2|500719603|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1327|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|235|Green||2015-10-09|2015-10-22|2016-06-13|Child: Changed school/site|Child: Changed school/site||7.7||2|2|2|2|F|Black||11|No|Relative: Other|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||17|28269|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503644199|503646159|31|0|2|504296433|31|0|2|500846365|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1328|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|525|Green|PERL 2014-2016|2015-09-23|2015-09-29|NaT||||17.2||1|1|1|1|M|Black||11|No|Mother|28214|4|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28273|Bachelors Degree|Single|Insurance|28226|7|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|504153965|504156015|31|0|1|504372591|1|0|1|500841770|10|2|-2||2|1|500014681|-2||-2|0|4|||7464|9|||1|500014681|7089569121628268952|0
M1329|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1362|Green||2013-06-11|2013-06-14|NaT||||44.7||1|1|3|3|F|Hispanic||11|No|Mother|28269|2|Two Parent|Unknown|||Y|Yes||Relative|General Community||Match Support|F|Hispanic||37|28203|Some College|Single|Education: Teacher|28217|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020753|503470937|502831178|3|0|2|500188541|3|0|2|500700189|10|2|-2||2|1||-2|500000294|-2|0|3|||2238|7|||1||6713311931049891381|0
M1330|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|103|Green||2016-11-11|2016-11-24|NaT||||3.4||1|1|1|1|F|White||11|No|Father|29715|6|One Parent: Male|$50,000 to $59,999||||Yes||Self|General Site||Match Support|F|White||38|28277|Juris Doctorate (JD)|Married|Law: Lawyer||6|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504886558|504889078|1|0|2|504822645|1|0|2|500927134|10|1|500009132|2128233620|2|1||-1||-1|0|10|||7464|9|||1||1174067921639243853|0
M1331|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-21|2016-11-30|NaT||||3.2||1|1|2|2|F|Black||11|Yes|Mother|28211|5|Two Parent|Less than $10,000|||Y|Yes||Relative|General Site||Match Support|F|Black||18|28213|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504944637|504947188|31|0|2|504324154|31|0|2|500929894|10|1|500000296|2128173564|2|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1332|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|104|Green||2016-11-23|2016-11-23|NaT||||3.4||1|1|1|1|M|Multi-race (Black & White)||11|No|Mother|29715|6|One Parent: Female|$50,000 to $59,999||||Yes||School|General Site||Match Support|M|White||68|28208|Masters Degree|Married|Finance|29715|2|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504908775|504911295|36|0|1|504806684|1|0|1|500930711|10|1|500009132|2128233620|2|1||-1||-1|0|4|||7464|9|||1||1174067921639243853|6156547733130613405
M1333|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|589|Green||2014-10-04|2014-10-22|2016-06-02|Child: Graduated|Child: Graduated||19.4||1|1|1|1|M|Hispanic||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28210||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020908|504041849|504043867|3|0|1|503995703|1|0|1|500780598|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1334|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|515|Green||2015-01-26|2015-01-29|2016-06-27|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||16.9||1|1|1|1|M|Black||11|No|GrandMother|28025|4|Grandparents|Unknown||||Yes||School|General Site|Cabarrus County|Enrollment|F|White||18|28036||Single|Student: High School||0|0||High School Partner|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504110036|504112070|31|0|1|504043678|1|0|2|500810175|5|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||0|4|||1||3575183301237417432|0
M1335|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|659|Green||2013-09-30|2013-09-30|2015-07-21|Volunteer: Moved|Volunteer: Moved||21.7||2|2|1|1|F|Black||11|Yes|Father|28212|3|One Parent: Male|Unknown||||Yes||School|General Site|Amachi|Match Support|F|Black||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503629844|503631783|31|0|2|503608281|31|0|2|500714467|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1336|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|231|Green||2015-10-09|2015-10-22|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.6||2|2|2|2|F|Black||11|Yes|Father|28212|3|One Parent: Male|Unknown||||Yes||School|General Site|Amachi|Match Support|F|White||18|28207|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503629844|503631783|31|0|2|504307866|1|0|2|500846367|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1337|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|265|Green||2014-09-22|2014-09-25|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.7||1|1|3|3|M|Black||11|No|Father|28208|4|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|M|White||30|28202|Bachelors Degree|Single|Finance: Accountant|28202|2|0|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|504030027|504015306|31|0|1|503908898|1|0|1|500777117|10|1|500009132|2128173561|4|1||-1||-1|0|4|||12831|3|||1||7960300212314874874|0
M1338|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|600|Green|PERL 2014-2016|2015-01-06|2015-02-05|2016-09-27|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19.7||3|3|2|2|M|Hispanic||11|No|Mother|28206|5|One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|M|Hispanic||28|28217|Bachelors Degree|Single|Finance|28202|2|5|Self|Self|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500016270|503408595|503410452|3|0|1|503490264|3|0|1|500806665|10|1|500000295|2128173561|4|1|500011312, 500014681|-1|500014681|-1|0|4|||7464|9|||1|500014681|7960300212314874874|0
M1339|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-11|2016-12-02|NaT||||3.1||1|1|2|2|M|Hispanic||11|No|Father|29715|6|One Parent: Male|$30,000 to $34,999||||No||School|General Site||Match Support|M|White||40|28273||Married|Finance|28217|10|0|LPL Financial|Workplace Partner|Big|General Site|VOL - PreMatch|Match Support|0|1|0|1|277|60|598|500000170|500013781|504870394|504872913|3|0|1|504557665|1|0|1|500927099|10|1|500009132|2128233620|2|1||-1|500007920|-1|0|4|||11247|3|||1||1174067921639243853|0
M1340|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|267|Green|PERL 2014-2016|2014-09-12|2014-09-23|2015-06-17|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.8||1|1|1|1|M|Black||11|No|Mother|28206|4|One Parent: Female|Unknown|||Y|Yes||School|General Site|PERL 2014-2016|Match Support|M|White||33|28269|Bachelors Degree|Married|Tech: Management|28202|3|6|Ally Financial|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500016270|503996736|503998751|31|0|1|503880784|1|0|1|500775712|10|1|500009132|2128173561|4|1|500014681|-1|500014681|-1|0|4|||12831|3|||1|500014681|7960300212314874874|0
M1341|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|806|Green|PERL 2014-2016|2014-12-19|2014-12-22|NaT||||26.5||1|1|1|1|M|Black||11|No|Mother|28226|3|One Parent: Female|$30,000 to $34,999||||No||School|General Community|PERL 2014-2016|Match Support|M|White||34|28214|Bachelors Degree||Transport: Flight Attendant|21804|7|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500018851|504083467|504085496|31|0|1|504003996|1|0|1|500805363|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681|4726905079488957916|1427172337358308252
M1342|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|55|Green||2017-01-08|2017-01-11|NaT||||1.8||2|2|1|1|F|Black||11|No|Mother|28217|6|Two Parent|$20,000 to $24,999||||Yes||Relative|General Site||Match Support|F|Some Other Race||33|28210|Bachelors Degree|Married|Finance|28205|1|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504861175|504863694|31|0|2|504952358|41|0|2|500938917|10|1|500009132|2128207318|2|1||-1||-1|0|3|||7464|9|||1||2611337051335117774|0
M1343|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|75|Green||2016-10-04|2016-10-20|2017-01-03|Volunteer: Time constraint|Volunteer: Time constraint||2.5||2|2|3|3|F|Black||11|No|Mother|28217|6|Two Parent|$20,000 to $24,999||||Yes||Relative|General Site||Match Support|F|White||28|28203|Bachelors Degree|Single|Finance|28202|0|6|Ally Financial|Workplace Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504861175|504863694|31|0|2|504349844|1|0|2|500912231|10|1|500009132|2128207318|4|1||-1||-1|0|3|||12831|3|||1||2611337051335117774|0
M1344|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1042|Green||2014-04-16|2014-04-30|NaT||||34.2||1|1|1|1|M|Black||11|No|Mother|28216|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||29|28202|Bachelors Degree|Single|Finance|28202|1|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020910|503503497|503505371|31|0|1|503775803|1|0|1|500759857|10|2|-2||2|1|500000294|-2|500000294|-2|0|10|||7464|9|||1||6077912216232501082|0
M1345|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|651|Green||2013-10-07|2013-10-07|2015-07-20|Volunteer: Moved|Volunteer: Moved||21.4||2|2|1|1|M|Hispanic||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503637763|503639718|3|0|1|503507441|1|0|1|500716283|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1346|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|240|Green||2015-10-09|2015-10-13|2016-06-09|Child: Changed school/site|Child: Changed school/site||7.9||2|2|2|2|M|Hispanic||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28211|Some College|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503637763|503639718|3|0|1|504307795|1|0|1|500846370|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1347|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|138|Green||2016-10-04|2016-10-20|NaT||||4.5||1|1|1|1|F|Black||11|No|Mother|28208|6|Two Parent|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|Black||35|28213|Masters Degree|Married|Business|28202|2|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504878263|504880783|31|0|2|504797062|31|0|2|500912540|10|1|500009132|2128207318|2|1||-1||-1|0|4|||7464|9|||1||2611337051335117774|0
M1348|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|651|Green||2013-10-07|2013-10-07|2015-07-20|Volunteer: Moved|Volunteer: Moved||21.4||3|3|1|1|M|Multi-race (Black & White)||11|No|Father|28211|1|One Parent: Male|Unknown||||No||School|General Site||Match Support|M|White||20|28277|Some High School||Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|502749239|502750151|36|0|1|503507342|1|0|1|500716287|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1349|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|244|Green||2015-10-09|2015-10-13|2016-06-13|Child: Changed school/site|Child: Changed school/site||8||3|3|2|2|M|Multi-race (Black & White)||11|No|Father|28211|1|One Parent: Male|Unknown||||No||School|General Site||Match Support|M|White||18|28036|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|502749239|502750151|36|0|1|503905466|1|0|1|500846261|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1350|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|428|Green||2015-12-14|2016-01-04|NaT||||14.1||1|1|1|1|M|Black||11|Yes|Mother|28208|5|One Parent: Female|Less than $10,000||||Yes||Relative|General Site||Match Support|M|Black||37|28277|Bachelors Degree|Married|Arts, Entertainment, Sports|28277|1|0|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504526251|504528583|31|0|1|504475303|31|0|1|500867619|10|1|500000295|2128207319|2|1||-1||-1|0|3|||18809|8|||1||3935539763241716148|0
M1351|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|426|Yellow||2014-12-02|2014-12-02|2016-02-01|Volunteer: Time constraint|Volunteer: Time constraint||14||1|1|1|1|F|Black||11||Mother|28031|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||30|28031|Bachelors Degree|Married|Medical: Nurse|28203|0|6|BBBS National Site|Web Link|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|504134537|504136574|31|0|2|503852298|1|0|2|500800216|10|1|500000295|2128173570|4|2||-1||-1|0|4|||46|2|||1||8034889377453131101|0
M1352|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|362|Green||2014-09-29|2014-10-09|2015-10-06|Child: Changed school/site|Child: Changed school/site||11.9||1|1|1|1|M|White||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504005669|504007684|1|0|1|503908386|1|0|1|500778963|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1353|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green||2016-11-28|2016-11-28|NaT||||3.3||1|1|1|1|F|White||11|No|Mother|29715|6|Two Parent|$30,000 to $34,999|Yes: Active|No||Yes||School|General Site||Match Support|F|White||26|28203|Bachelors Degree|Single|Finance|29175|0|6|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504942804|504945355|1|0|2|504807056|1|0|2|500931105|10|1|500009132|2128233620|2|1||-1||-1|0|4|||7464|9|||1||1174067921639243853|5471818036158225409
M1354|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|973|Red|Amachi|2012-04-13|2012-05-23|2015-01-21|Volunteer: Moved|Volunteer: Moved||32|Y|1|1|1|1|M|Black||11|Yes|Mother|28278||One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community|Amachi|Match Support|F|White||34|29710|Bachelors Degree|Married|Education: Teacher||0|6|Relative|Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502464508|502211737|31|0|1|502901720|1|0|2|500609874|10|2|500003586||4|3|500000294|-2||-2|0|10|||17161|11|||1|500000294|0|0
M1355|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|113|Green||2016-11-02|2016-11-14|NaT||||3.7||1|1|1|1|F|Black||11|No|Mother|28269|6|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||39|28269|Bachelors Degree|Single|Govt|28202|1|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504628103|504630514|31|0|2|504469742|31|0|2|500922796|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1||1320477920662455183|4825213036474521167
M1356|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|649|Green|PERL 2014-2016, Cabarrus County|2015-05-11|2015-05-28|NaT||||21.3||1|1|1|1|M|Black||11|No|Mother|28027|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||31|28027|Juris Doctorate (JD)|Married|Law: Lawyer|28036|2|10|Igniting Breakfast|Special Event|Big|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|502426625|502502446|31|0|1|504274174|1|0|1|500826502|10|2|500016307||2|1|500014681, 500016374|-2|500000294, 500014681, 500016374|-2|0|10|||17266|8|||1|500014681, 500016374|7075115687862385692|2581014289501540602
M1357|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|455|Green||2013-11-27|2013-12-19|2015-03-19|Child/Family: Moved|Child/Family: Moved||14.9||1|1|1|1|F|Black||11|No|Mother|2649|4|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Education: Teacher|28012|3|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500015820|503569115|503570990|31|0|2|503619714|1|0|2|500735248|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||4903779310522421428|7674215580094440446
M1358|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|134|Green||2016-10-12|2016-10-24|NaT||||4.4||1|1|1|1|M|Multi-race (Black & White)||11|No|Mother|28212|6|One Parent: Female|$50,000 to $59,999||||Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||22|28202|Bachelors Degree|Single|Tech: Sales, Mktg|28202|0|2|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|503623886|503625775|36|0|1|504803107|1|0|1|500915035|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||2811191761055817959|5499465424599250965
M1359|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|1147|Green|VOL - Mentoring Hispanic Youth|2013-12-09|2013-12-17|2017-02-06|Child: Graduated|Child: Graduated||37.7||1|1|1|1|M|Hispanic||11|No|Mother|28217|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||26|28210|Bachelors Degree|Married|Business: Sales|28234|0|5|Recruitment Event|BBBS Board/Staff|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|503745242|503747214|3|0|1|503480703|1|0|1|500737636|10|1|500000295|2128173557|4|1||-1|500000294|-1|0|4|||7462|13|||1|500011312|8981704271528751143|0
M1360|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1819|Yellow||2012-02-08|2012-03-14|NaT||||59.8||1|1|1|1|F|Black||11|No|GrandMother|28205||Grandparents|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||40|28227|Masters Degree|Married|Tech: Support, Writing|28262|11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502859181|500187987|31|0|2|502638002|1|0|2|500597079|10|2|-2||2|2||-2||-2|0|10|||7462|13|||1||7960300212314874874|0
M1361|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|386|Green||2014-07-09|2014-07-23|2015-08-13|Volunteer: Time constraint|Volunteer: Time constraint||12.7||1|1|1|1|F|Black||11|No|Mother|28208|5|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||RTBM|F|White||28|28211|Bachelors Degree|Single|Child/Day Care Worker||0|8|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503795417|503797394|31|0|2|503762193|1|0|2|500769015|7|2|-2||4|1||-2||-2|0|5|||17159|12|||1||5386346637278076349|2141487034287122220
M1362|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|572|Green||2014-03-12|2014-03-26|2015-10-19|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||18.8||2|2|1|1|M|Black||11|No|Mother|28025|4|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||73|28226|PHD|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503741920|503743892|31|0|1|503696505|1|0|1|500754344|10|2|-2||4|1|500016374|-2||-2|0|10|||7464|9|||1||0|5503100293073900724
M1363|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|19|Green||2017-01-23|2017-02-16|NaT||||0.6||2|2|1|1|M|Black||11|No|Mother|28025|4|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||30|28075|Bachelors Degree|Married|Business: Sales|28213|6|3|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|503741920|503743892|31|0|1|504976126|1|0|1|500941524|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||17159|12|||1||0|5503100293073900724
M1364|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green||2016-11-11|2016-11-28|NaT||||3.3||1|1|1|1|M|White||11|No|Mother|29715|6|One Parent: Female|$50,000 to $59,999||||No||School|General Site||Match Support|M|White||36|28202||Single|Business: Mgt, Admin||6|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504870414|504872933|1|0|1|504787136|1|0|1|500927126|10|1|500009132|2128233620|2|1||-1||-1|0|4|||7464|9|||1||1174067921639243853|0
M1365|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|98|Green||2016-10-24|2016-11-29|NaT||||3.2||1|1|1|1|F|Black||11|No|Mother|28209|5|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||23|28203|Bachelors Degree||Finance: Accountant|28031|0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504662612|504665039|31|0|2|504595097|1|0|2|500918825|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||6627885846854295604|2719955880210213907
M1366|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|464|Green||2013-11-18|2013-11-20|2015-02-27|Child: Graduated|Child: Graduated||15.2||1|1|1|1|M|Black||11|No|Mother|28216|3|One Parent: Female|Unknown|||Y|Yes||Self|General Site||Match Support|M|White||29|28209|Bachelors Degree|Single|Business: Engineer|28208|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500008321|503718051|503720018|31|0|1|503489016|1|0|1|500732255|10|1|-1||4|1||-1||-1|0|10|||7496|10|||1||8568001799025358453|0
M1367|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1786|Green||2012-03-20|2012-04-16|NaT||||58.7||2|2|2|2|F|Black||11|No|Mother|28208|3|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|Black||41|28209|Bachelors Degree|Single|Finance: Banking|28255|0|6|TV|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502298007|502234907|31|0|2|501202092|31|0|2|500605225|10|2|-2||2|1|500004640|-2||-2|0|10|||130|1|||1||2611337051335117774|5656517387001249169
M1368|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|368|Green||2014-12-04|2015-01-30|2016-02-02|Volunteer: Moved|Volunteer: Moved||12.1||2|2|1|1|M|Black||11|No|Mother|28205|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||33|28206|Masters Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504059510|503637389|31|0|1|504000163|31|0|1|500801345|10|1|500000295|2128173561|4|1||-1||-1|0|4|||46|2|||1||7960300212314874874|0
M1369|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|79|Green||2016-02-22|2016-05-03|2016-07-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||2.6||2|2|1|1|M|Black||11|No|Mother|28205|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||27|28203|Bachelors Degree|Single|Finance: Banking|28244|1|2|Self|Self|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500016270|504059510|503637389|31|0|1|504359587|31|0|1|500880682|10|1|500000295|2128173561|4|1||-1|500007920, 500011315, 500011316|-1|0|4|||7464|9|||1||7960300212314874874|0
M1370|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|519|Green||2015-03-18|2015-04-16|2016-09-16|Child: Lost interest|Child: Lost interest||17.1||1|1|1|1|F|Black||11|No|Father|28205|4|One Parent: Male|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Black||56|28216|High School Graduate|Married|Unemployed||0|0|United Way|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|504221885|504223999|31|0|2|504188499|31|0|2|500819243|10|2|-2||4|1||-2||-2|0|4|||16263|6|||1||5822146217251000296|0
M1371|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1442|Green||2013-03-13|2013-03-26|NaT||||47.4||1|1|1|1|M|White||11|No|Mother|28269|3|Other/Unknown|$15,000 to $19,999||||Yes||School|General Community||Match Support|M|White||47|28278|Bachelors Degree|Married|Finance: Banking|28210|0|8|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502842247|502843540|1|0|1|503305101|1|0|1|500687640|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||967246839551912690|2094153948849884702
M1372|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|608|Green||2014-10-04|2014-10-07|2016-06-06|Volunteer: Moved|Volunteer: Moved||20||2|2|1|1|F|Hispanic||11|No|Father|28212|3|One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049252|504051276|3|0|2|503901627|1|0|2|500780589|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1373|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-16|2016-11-30|NaT||||3.2||2|2|2|2|F|Hispanic||11|No|Father|28212|3|One Parent: Male|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||18|28173|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504049252|504051276|3|0|2|504297141|31|0|2|500928423|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1374|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|374|Green||2014-09-29|2014-09-30|2015-10-09|Child: Changed school/site|Child: Changed school/site||12.3||2|2|2|2|M|Black||11||Mother|28217|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503198334|503200089|31|0|1|503907463|1|0|1|500778747|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1375|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|967|Green|VOL - Mentoring Hispanic Youth|2014-07-08|2014-07-14|NaT||||31.8||1|1|1|1|F|Hispanic||11|Yes|GrandMother|28216|2|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||30|28203|Masters Degree|Single|Medical: Pharmacist|28213|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503904008|503906008|3|0|2|503820652|1|0|2|500768869|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1|500011312|3664007741235143067|0
M1376|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|148|Green|PERL 2014-2016|2016-09-06|2016-10-10|NaT||||4.9||1|1|1|1|M|Black||11|No|Mother|28210|5|One Parent: Female|$50,000 to $59,999||||No||Self|General Community|PERL 2014-2016|Match Support|M|Native Hawaiian or Other Pacific Islander||26|28209|Bachelors Degree|Single|Business: Engineer|28202|1|8|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504714089|504716526|31|0|1|504679648|5|0|1|500906166|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|500014681|4902029756574603597|3402014428779854546
M1377|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|368|Green||2015-10-05|2015-10-19|2016-10-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12.1||2|2|1|1|F|Black||11|No|Mother|28203|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||33|28210|PHD|Single|Medical|28105|1|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|504388136|504390375|31|0|2|504360253|1|0|2|500844373|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1||8568001799025358453|2876415545463317777
M1378|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|76|Green||2016-12-08|2016-12-21|NaT||||2.5||2|2|2|2|F|Black||11|No|Mother|28203|6|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||26|28210|Bachelors Degree|Single|Medical: Admin|28209|1|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500013781|504388136|504390375|31|0|2|503869569|1|0|2|500934047|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||8568001799025358453|2876415545463317777
M1379|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|400|Green||2016-01-06|2016-02-01|NaT||||13.1||1|1|5|5|M|Hispanic||11|No|Mother|28217|5|Two Parent|$20,000 to $24,999||||Yes||School|General Site||Match Support|M|White||48|28209|Bachelors Degree|Married|Business: Mgt, Admin|28217|21|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504526331|504528663|3|0|1|500994796|1|0|1|500870411|10|1|500000295|2128207319|2|1||-1||-1|0|4|||7464|9|||1||3935539763241716148|0
M1380|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|791|Red||2014-04-10|2014-04-29|2016-06-28|Volunteer: Moved|Volunteer: Moved||26||2|2|1|1|F|Hispanic||11|No|Mother|28212|2|Two Parent|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||29|28206|Masters Degree|Single|Finance: Accountant|28210|3|0|United Way|Service Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017777|502619308|502619917|3|0|2|503710698|1|0|2|500759246|10|2|-2||4|3||-2|500000294|-2|0|10|||16263|6|||1||2417657944362725638|0
M1381|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1042|Green||2014-04-21|2014-04-30|NaT||||34.2||1|1|1|1|M|Black||11|No|Mother|28215|2|One Parent: Female|$45,000 to $49,999||||No||Self|General Community||Match Support|M|White||37|28205|Bachelors Degree|Married|Finance|28205|0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503545940|503547815|31|0|1|503804018|1|0|1|500760430|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1||0|3402014428779854546
M1382|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|159|Green|PERL 2014-2016|2016-09-14|2016-09-29|NaT||||5.2||1|1|1|1|F|Black||11|No|Mother|28031|4|Two Parent|$15,000 to $19,999|||Y|No||School|General Community|PERL 2014-2016|Match Support|F|White||44|28031|Masters Degree|Married|Education||0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500017732|504577421|504579758|31|0|2|504771021|1|0|2|500907629|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681|0|7137064858903755892
M1383|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|587|Green||2014-10-04|2014-10-28|2016-06-06|Volunteer: Moved|Volunteer: Moved||19.3||2|2|1|1|M|Hispanic||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049238|504051262|3|0|1|503907477|1|0|1|500780597|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1384|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|M|Hispanic||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504049238|504051262|3|0|1|504297082|1|0|1|500929312|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1385|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|241|Red|PERL 2014-2016|2015-06-28|2015-06-28|2016-02-24|Child/Family: Time constraints|Child/Family: Time constraints||7.9||1|1|2|2|M|Black||11|No|Mother|28226|3|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500013781|504198439|504200550|31|0|1|504230177|1|0|1|500831539|10|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||7462|13|||1|500014681|6368218764956286027|0
M1386|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|617|Green||2013-11-10|2013-11-11|2015-07-21|Volunteer: Moved|Volunteer: Moved||20.3||2|2|1|1|F|Multi-race (Black & White)||11|No|Mother|28211|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503704249|503706214|36|0|2|503497234|1|0|2|500729568|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1387|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|181|Green||2015-10-09|2015-10-21|2016-04-19|Child/Family: Moved|Child/Family: Moved||5.9||2|2|2|2|F|Multi-race (Black & White)||11|No|Mother|28211|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|503704249|503706214|36|0|2|504303308|1|0|2|500846337|10|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1388|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|216|Green||2016-02-18|2016-02-26|2016-09-29|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||7.1||2|2|1|1|M|Black||11|No|Mother|28025|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|Cabarrus County|Match Support|M|White||19|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504619450|504621861|31|0|1|504619589|1|0|1|500880034|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||643003066716863548|0
M1389|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|112|Green|Cabarrus County|2016-10-17|2016-11-15|NaT||||3.7||2|2|1|1|M|Black||11|No|Mother|28025|5|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|Cabarrus County|Match Support|M|Black||17|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504619450|504621861|31|0|1|504884038|31|0|1|500916292|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|643003066716863548|0
M1390|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|726|Green||2015-03-03|2015-03-12|NaT||||23.9||1|1|1|1|M|Black||11|No|Mother|28215|3|One Parent: Female|$30,000 to $34,999||||Yes||School|General Community||Match Support|M|Black||44|28173|Masters Degree|Married|Tech: Computer/Programmer|28202|7|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503794892|503796869|31|0|1|504175530|31|0|1|500816649|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||5741767063897867874|3643651798871536206
M1391|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|613|Green||2014-10-07|2014-10-09|2016-06-13|Volunteer: Moved|Volunteer: Moved||20.1||2|2|1|1|F|Black||11|No|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504041768|504043786|31|0|2|503907444|1|0|2|500781516|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1392|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|90|Green||2016-11-18|2016-12-07|NaT||||3||2|2|2|2|F|Black||11|No|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||17|28269|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504041768|504043786|31|0|2|504296433|31|0|2|500929353|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1393|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|48|Green||2016-12-05|2017-01-18|NaT||||1.6||1|1|2|2|F|Hispanic||11|No|Father|28211|5|One Parent: Male|$20,000 to $24,999|||Y|Yes||Self|General Site||Match Support|F|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504937026|504939577|3|0|2|504303240|1|0|2|500933236|10|1|500000296|2128173564|2|1||-1||-1|0|10|||0|4|||1||2762897743412756173|0
M1394|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|499|Green||2015-10-16|2015-10-20|2017-03-02|Volunteer: Time constraint|Volunteer: Time constraint||16.4||1|1|1|1|M|Black||11|No|Mother|28212|4|One Parent: Female|$15,000 to $19,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|White||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504468539|504470812|31|0|1|504306056|1|0|1|500848710|10|1|500000296|2128173564|4|1|500014068|-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1395|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|350|Red||2016-03-02|2016-03-22|NaT||||11.5||1|1|1|1|F|Black||11|No|Mother|28208|5|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site||Match Support|F|White||28|28205|Bachelors Degree|Single|Journalist/Media|28217|3|8|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504526307|504528639|31|0|2|504441484|1|0|2|500882703|10|1|500000295|2128207319|2|3||-1||-1|0|4|||46|2|||1||3935539763241716148|0
M1396|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|498|Green||2014-03-12|2014-04-08|2015-08-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||16.4||1|1|2|2|F|Black||11|No|Mother|28209|K|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||28|28212|Masters Degree|Single|Customer Service|28202|3|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503418236|503420100|31|0|2|503671882|31|0|2|500754333|10|1|-1||4|1||-1||-2|0|4|||7464|9|||1||8568001799025358453|0
M1397|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|403|Green||2015-12-18|2016-01-29|NaT||||13.2||1|1|1|1|M|Hispanic||11|No|Mother|28208|4|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||45|28227|Some College|Divorced|Self-Employed, Entrepreneur|28277|15|0|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504531588|504533921|3|0|1|504127246|1|0|1|500868809|10|1|500000295|2128207319|2|1||-1||-1|0|4|||17159|12|||1||3935539763241716148|0
M1398|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|313|Green||2014-11-09|2014-12-04|2015-10-13|Child: Changed school/site|Child: Changed school/site||10.3||1|1|2|2|F|Black||11|No|Mother|28213|3|Two Parent|Unknown||||No||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504093590|504095620|31|0|2|503907351|1|0|2|500793663|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1399|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|593|Green||2014-10-04|2014-10-22|2016-06-06|Volunteer: Moved|Volunteer: Moved||19.5||1|1|1|1|M|Black||11|No|Father|28212|3|One Parent: Male|Unknown|||Y|Yes||School|General Site||RTBM|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504042013|504044031|31|0|1|503999137|1|0|1|500780599|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1400|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|11|Green||2017-02-20|2017-02-24|NaT||||0.4||1|1|1|1|F|Black||11|No|Mother|28208|4|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Black||23|28208|Associate Degree|Single|Medical||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504970052|504972603|31|0|2|504743981|31|0|2|500947288|10|1|500000295|2128207319|2|1||-1||-1|0|4|||7464|9|||1||3935539763241716148|0
M1401|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-22|2016-11-30|NaT||||3.2||1|1|3|3|F|White||11|No|Father|28211|5|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Site||Match Support|F|White||18|28207|Some College|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504952387|504954938|1|0|2|504306107|1|0|2|500930367|10|1|500000296|2128173564|2|1||-1||-1|0|10|||0|4|||1||2762897743412756173|0
M1402|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|289|Green||2014-10-04|2014-10-22|2015-08-07|Volunteer: Moved|Volunteer: Moved||9.5||3|3|2|2|M|Hispanic||11|No|Mother|28203||One Parent: Female|Unknown||||No||School|General Site||Match Support|M|White||20|28226||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503214533|503646168|3|0|1|503540968|1|0|1|500780612|10|1|||4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1403|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|343|Green||2015-10-09|2015-10-26|2016-10-03|Child: Changed school/site|Child: Changed school/site||11.3||3|3|2|2|M|Hispanic||11|No|Mother|28203||One Parent: Female|Unknown||||No||School|General Site||Match Support|M|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503214533|503646168|3|0|1|504307950|1|0|1|500846334|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1404|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|758|Green||2013-09-25|2013-09-30|2015-10-28|Volunteer: Time constraint|Volunteer: Time constraint||24.9||2|2|1|1|M|Black||11||Mother|28208|4|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|Black||30|28027|Bachelors Degree|Married|Business: Clerical|28282|3|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020990|502982459|502983913|31|0|1|503565143|31|0|1|500713173|10|2|-2||4|1|500014681|-2||-2|0|10|||7464|9|||1||5548059939346196746|7044657180546140448
M1405|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|228|Green|PERL 2014-2016|2016-07-13|2016-07-22|NaT||||7.5||2|2|1|1|M|Black||11||Mother|28208|4|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||24|28204|Bachelors Degree||Arts, Entertainment, Sports|28201|0|8|Local TV|Media|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|502982459|502983913|31|0|1|504669593|1|0|1|500899540|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7438|1|||1|500014681|5548059939346196746|7044657180546140448
M1406|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|165|Green||2015-04-20|2015-05-04|2015-10-16|Child/Family: Moved|Child/Family: Moved||5.4||1|1|1|1|M|Black||11|Yes|Mother|28217|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||67|28277||Married|Retired||0|0|Other|Service Organization|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500020753|504184746|504186855|31|0|1|504183176|31|0|1|500824006|10|1|500000295|2128173557|4|1||-1||-1|0|4|||7452|6|||1||8981704271528751143|0
M1407|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|549|Red|PERL 2014-2016|2015-01-23|2015-02-06|2016-08-08|Child: Severity of challenges|Child: Severity of challenges||18||1|1|1|1|M|White||11|No|Mother|28081|3|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Hispanic||31|28083|Some College|Married|Business: Mgt, Admin||14|3|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500020753|504059549|504061573|1|0|1|504109643|3|0|2|500809931|10|2|-2||4|3|500014681, 500016374|-2|500014681, 500016374|-2|0|5|||46|2|||1|500014681|8568001799025358453|2141487034287122220
M1408|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|655|Green||2013-09-09|2013-09-20|2015-07-07|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||21.5||2|2|1|1|F|Black||11|Yes|Mother|28206|4|One Parent: Female|Unknown|||Y|Yes||Self|General Site||Match Support|F|Black||65|28110|Masters Degree|Single|Human Services||7|0|Self|Self|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500016270|503515718|503517589|31|0|2|503443502|31|0|2|500709607|10|1|500000295|2128173561|4|1||-1||-1|0|10|||7464|9|||1||7960300212314874874|0
M1409|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|248|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2015-10-27|2015-11-16|2016-07-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||8.1||2|2|1|1|F|Black||11|Yes|Mother|28206|4|One Parent: Female|Unknown|||Y|Yes||Self|General Site||Match Support|F|White||32|28207|Bachelors Degree|Single|Finance: Auditor|28202|8|10|Current/Previous Big|Other Big|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500016270|503515718|503517589|31|0|2|504368058|1|0|2|500852488|10|1|500000295|2128173561|4|1||-1|500007920, 500011315, 500011316|-1|0|10|||17159|12|||1|500007920, 500011315, 500011316|7960300212314874874|0
M1410|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|264|Green||2016-05-24|2016-06-16|NaT||||8.7||1|1|1|1|F|Black||11|No|Mother|28216|4|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||27|28209|Bachelors Degree|Single|Medical|28054|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504628520|504630931|31|0|2|504409458|1|0|2|500894207|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||2456895876914964961|7044657180546140448
M1411|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|231|Green||2014-10-04|2014-10-17|2015-06-05|Volunteer: Moved|Volunteer: Moved||7.6||3|3|2|2|M|Hispanic||11|Yes|Mother|28212||One Parent: Female|Unknown||||Yes||School|General Site|Amachi|Match Support|M|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503418298|503420158|3|0|1|503497508|1|0|1|500780602|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1412|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|518|Green||2015-10-06|2015-10-06|NaT||||17||3|3|1|1|M|Hispanic||11|Yes|Mother|28212||One Parent: Female|Unknown||||Yes||School|General Site|Amachi|Match Support|M|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|503418298|503420158|3|0|1|504303764|1|0|1|500844550|10|1|500000296|2128173564|2|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1413|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|766|Green|PERL 2014-2016, Cabarrus County|2015-01-22|2015-01-31|NaT||||25.2||2|2|1|1|F|White||11|No|Father|28081|4|One Parent: Male|Unknown||||Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||32|28226|Bachelors Degree|Married|Business: Mgt, Admin|10006|1|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|503634724|503636659|1|0|2|504107959|1|0|2|500809650|10|2|-2||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||17159|12|||1|500014681, 500016374|6810228174639243761|1786514887916898235
M1414|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|985|Green||2014-06-09|2014-06-26|NaT||||32.4||1|1|2|2|M|Black||11|No|Mother|28269|5|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||49|28031|Associate Degree||Customer Service||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503543014|503544889|31|0|1|503546166|1|0|1|500765902|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||220177803211026571|8243619853090168866
M1415|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|277|Green||2014-10-04|2014-10-17|2015-07-21|Volunteer: Moved|Volunteer: Moved||9.1||3|3|2|2|F|Hispanic||11|No|Mother|28227|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503254195|503256000|3|0|2|503608280|1|0|2|500780606|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1416|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|509|Green||2015-10-09|2015-10-15|NaT||||16.7||3|3|1|1|F|Hispanic||11|No|Mother|28227|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|503254195|503256000|3|0|2|504386413|1|0|2|500846388|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1417|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|378|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-10|2016-02-23|NaT||||12.4||1|1|1|1|M|Black||11|No|Mother|28262|3|One Parent: Female|$30,000 to $34,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504295805|504298006|31|0|1|504337975|1|0|1|500878715|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1|500007920, 500011315, 500011316|7102230088759381237|5923747279518652886
M1418|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|55|Green||2016-12-13|2017-01-11|NaT||||1.8||1|1|1|1|F|Black||11|No|Mother|28208|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||24|28203|Bachelors Degree|Single|Finance|28255|0|6|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504617847|504620258|31|0|2|504580008|1|0|2|500935128|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7462|13|||1||5711791743715234276|8408514790530965815
M1419|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1964|Green||2011-04-08|2011-04-14|2016-08-29|Child/Family: Moved|Child/Family: Moved||64.5||1|1|1|1|F|Black||11|No|Mother|28273||One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||61|28211|Bachelors Degree|Widowed|Real Estate: Realtor|28207|16|0|Other|BBBS Board/Staff|Big|General Community|Amachi, Project Big|Match Support|1|0|1|0|277|60|598|500000170|500017777|502425281|502425720|31|0|2|502529075|1|0|2|500530096|10|2|-2||4|1||-2|500000294, 500004640|-2|0|10|||7671|13|||1||0|0
M1420|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2191|Green||2011-02-24|2011-03-08|NaT||||72||1|1|1|1|F|Multi-race (Hispanic & White)||11|No|GrandMother|28210|K|Grandparents|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||31|28211|Bachelors Degree|Single|Finance: Banking|28255|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|1|0|0|1|277|60|598|500000170|500020753|502458411|502458858|35|0|2|502479222|1|0|2|500520070|10|2|-2||2|1||-2|500000294, 500004640|-2|6854|8|||7496|10|||1||0|0
M1421|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|25|Green|Cabarrus County|2017-02-03|2017-02-10|NaT||||0.8||2|2|1|1|M|Black||11|No|Mother|28025|4|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Cabarrus County|Match Support|M|White||56|28075|PHD|Married|Education: College Professor|28223|5|6|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504637328|504639739|31|0|1|504995988|1|0|1|500944447|10|2|500016307||2|1|500016374|-2|500016374|-2|0|4|||17159|12|||1|500016374|3575183301237417432|7044657180546140448
M1422|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|191|Yellow||2016-03-11|2016-03-22|2016-09-29|Child/Family: Moved|Child/Family: Moved||6.3||2|2|1|1|M|Black||11|No|Mother|28025|4|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Cabarrus County|Match Support|F|White||17|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504637328|504639739|31|0|1|504583576|1|0|2|500884254|10|1|500000296|2128173571|4|2|500016374|-2|500016374|-1|0|4|||7464|9|||1||3575183301237417432|7044657180546140448
M1423|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|62|Red|PERL 2014-2016|2015-02-12|2015-02-27|2015-04-30|Child: Severity of challenges|Child: Severity of challenges||2||1|1|1|1|M|Black||11|No|Mother|28202|2|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||26|28205|Bachelors Degree|Single|Business: Sales|28205|1|1|BBBS National Site|Web Link|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500008321|504003061|504005076|31|0|1|504169596|1|0|1|500813623|10|2|-2||4|3|500014681|-2||-2|34|2|||46|2|||1|500014681|6368218764956286027|8861782924354204409
M1424|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1439|Green|Amachi|2012-05-25|2012-06-11|2016-05-20|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||47.3||1|1|1|1|F|Black||11|Yes|Mother|28216|2|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||Enrollment|F|White||28|28202|Bachelors Degree|Single|Finance: Banking||0|9|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|502948870|503287812|31|0|2|502984009|1|0|2|500616576|5|2|-2||4|1||-2||-2|0|10|||7496|10|||1|500000294|6065435025527210335|0
M1425|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|601|Green||2013-10-08|2013-10-11|2015-06-04|Volunteer: Moved|Volunteer: Moved||19.7||1|1|1|1|M|Black||11|Yes|Mother|28204|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|M|White||20|28278|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503644166|503646126|31|0|1|503497274|1|0|1|500717211|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1426|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|208|Green|PERL 2014-2016, Cabarrus County|2016-08-09|2016-08-11|NaT||||6.8||1|1|1|1|F|Black||11|No|Mother|28025|4|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||25|28027|Some College|Single|Business: Sales||0|6|Community Engagement|Special Event|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504711954|504714390|31|0|2|504718024|1|0|2|500902765|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|34|2|||18809|8|||1|500014681, 500016374|0|7044657180546140448
M1427|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|576|Green||2013-10-15|2013-10-22|2015-05-21|Child/Family: Moved|Child/Family: Moved||18.9||1|1|1|1|F|Black||11|Yes|Mother|28227|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503637696|503639656|31|0|2|503540493|1|0|2|500719607|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1428|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1035|Green||2014-04-07|2014-05-07|NaT||||34||1|1|1|1|M|Black||11|No|Mother|28206|1|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||31|28204|Bachelors Degree|Single|Business|28262|1|9|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503381519|503383388|31|0|1|503803833|1|0|1|500758686|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||392688197545050058|5081726734274569781
M1429|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|90|Green||2016-11-30|2016-12-07|NaT||||3||1|1|2|2|F|Hispanic||11|No|Mother|28212|5|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504944612|504504693|3|0|2|504297059|1|0|2|500931725|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1430|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|154|Green||2014-10-07|2014-10-28|2015-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.1||1|1|1|1|F|Black||11|No|Mother|28206|2|One Parent: Female|Unknown||||No||School|General Site||Match Support|F|Black||24|28215||Single|Student: High School|28223|0|0|Recruitment Event|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503217195|503218976|31|0|2|503695805|31|0|2|500781086|10|1|500000295|2128173561|4|1||-1||-1|0|4|||7458|9|||1||7960300212314874874|0
M1431|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|495|Green||2015-01-30|2015-01-30|2016-06-08|Volunteer: Moved|Volunteer: Moved||16.3||2|2|2|2|F|Black||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28222|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504184145|504186254|31|0|2|503907282|1|0|2|500811308|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1432|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|F|Black||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504184145|504186254|31|0|2|504308470|1|0|2|500929304|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1433|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|113|Green||2016-10-24|2016-11-14|NaT||||3.7||1|1|1|1|M|Black||11|Yes|Mother|28217|4|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|M|White||27|28278||Single|Business|28208|0|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504456498|504458770|31|0|1|504766383|1|0|1|500918854|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||0|5597049740348738
M1434|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|511|Green||2015-10-05|2015-10-13|NaT||||16.8||2|2|1|1|F|Black||11|No|Mother|28269|5|One Parent: Female|$50,000 to $59,999|||Y|No||School|General Community||Match Support|F|Black||41|28216|Bachelors Degree|Single|Business|28282|2|11|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504243465|504245581|31|0|2|504365625|31|0|2|500844251|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||0|2806833304218536184
M1435|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|56|Green||2015-04-23|2015-04-30|2015-06-25|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||1.8||2|2|1|1|F|Black||11|No|Mother|28269|5|One Parent: Female|$50,000 to $59,999|||Y|No||School|General Community||Match Support|F|White||27|28202|Some College|Single|Transport: Flight Attendant||2|1|Local TV|Media|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500017732|504243465|504245581|31|0|2|504173742|1|0|2|500824646|10|2|-2||4|1||-2||-2|0|4|||7438|1|||1||0|2806833304218536184
M1436|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|153|Green||2014-10-07|2014-10-21|2015-03-23|Child/Family: Moved|Child/Family: Moved||5||1|1|1|1|M|Hispanic||11|Yes|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||RTBM|1|0|1|0|277|60|598|500000170|500019116|504049414|504031221|3|0|1|503898561|1|0|1|500781528|10|1|||4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1437|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|994|Green||2013-11-13|2013-12-09|2016-08-29|Child: Lost interest|Child: Lost interest||32.7||1|1|1|1|M|Black||11|No|Mother|28227|3|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|M|White||38|28203||Single|Finance|28202|16|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503067218|503068877|31|0|1|503526377|1|0|1|500730492|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1||8979408036987322141|7701000190042603388
M1438|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|1547|Green||2012-12-11|2012-12-11|NaT||||50.8||1|1|1|1|M|Black||11|Yes|Mother|28217|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||55|28078|Some College|Married|Business: Sales|28217|24|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|1|0|0|1|277|60|598|500000170|500021785|503329148|503330982|31|0|1|503225539|1|0|1|500668735|10|1|500000295|2128173557|2|1||-1||-1|0|4|||7496|10|||1||8981704271528751143|0
M1439|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1006|Green||2014-05-19|2014-06-05|NaT||||33.1||1|1|1|1|M|Black||11|No|Mother|28205|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||49|28205|Masters Degree|Domestic Partner|Business: Mgt, Admin|28277|3|9|Agency Sponsored|Special Event|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503737886|503739858|31|0|1|503844296|1|0|1|500763770|10|2|-2||2|1||-2||-2|0|10|||16426|8|||1||421482027904269589|0
M1440|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|920|Green||2014-08-30|2014-08-30|NaT||||30.2||1|1|1|1|F|Black||11|No|Mother|28205|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||37|28105|Masters Degree|Single|Education: Teacher||2|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020910|503764144|503739858|31|0|2|503784339|31|0|2|500773966|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||421482027904269589|0
M1441|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1007|Green|Cabarrus County|2014-05-05|2014-06-04|NaT||||33.1||1|1|1|1|M|Black||11|No|Mother|28083|2|One Parent: Female|$45,000 to $49,999|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|Black||50|28075|Masters Degree|Married|Law|28212|25|1|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|503694415|503696380|31|0|1|503723380|31|0|1|500762190|10|2|500016307||2|1|500016374|-2|500016374|-2|34|2|||7464|9|||1|500016374|6720734052660262632|8084353152153143886
M1442|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2016-12-06|2017-01-30|NaT||||1.2||1|1|1|1|M|Black||11|No|Mother|28202|4|One Parent: Female|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||50|28210|Bachelors Degree|Married|Finance|28202|15|0|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504700175|504702604|31|0|1|504649796|1|0|1|500933583|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||18809|8|||1||6368218764956286027|6761707515712559257
M1443|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|837|Green||2014-11-12|2014-11-21|NaT||||27.5||1|1|1|1|M|Black||11|Yes|Mother|28227|3|One Parent: Female|$30,000 to $34,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||29|28210|Bachelors Degree|Single|Tech: Sales, Mktg|28262|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503956230|503958239|31|0|1|504026743|31|0|1|500795032|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1||0|8913351025023100786
M1444|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|601|Green||2014-10-07|2014-10-14|2016-06-06|Volunteer: Moved|Volunteer: Moved||19.7||2|2|1|1|F|Black||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049221|504051245|31|0|2|503897618|1|0|2|500781526|10|1|500000296|2128173564|4|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1445|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-18|2016-11-30|NaT||||3.2||2|2|2|2|F|Black||11|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504049221|504051245|31|0|2|504306171|1|0|2|500929334|10|1|500000296|2128173564|2|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1446|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|762|Red||2015-01-24|2015-01-28|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25||1|1|1|1|M|Black||11|No|GrandMother|28215|1|One Parent: Female|$35,000 to $39,999|||Y|Yes||School|General Community||Enrollment|M|White||26|28205|Bachelors Degree|Single|Business: Mgt, Admin|28205|1|7|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500020753|503853254|503855248|31|0|1|504163053|1|0|1|500809956|5|2|-2||4|3||-2|500000294|-2|0|4|||17159|12|||1||3723482195151978288|0
M1447|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|398|Green||2016-01-05|2016-02-03|NaT||||13.1||1|1|1|1|F|Black||11|No|Mother|28208|5|One Parent: Female|$15,000 to $19,999||||Yes||Relative|General Site||Match Support|F|Black||35|28278|Masters Degree|Married|Homemaker|10801|0|0|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504526285|504528617|31|0|2|504530191|31|0|2|500870373|10|1|500000295|2128207319|2|1||-1||-1|0|3|||17159|12|||1||3935539763241716148|0
M1448|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|712|Yellow||2015-03-10|2015-03-26|NaT||||23.4||1|1|1|1|F|Black||11|No|Mother|28227|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||29|28226|Bachelors Degree|Single|Finance: Accountant|28202|0|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504194601|504184323|31|0|2|504032490|1|0|2|500817776|10|2|-2||2|2||-2||-2|0|4|||7464|9|||1||8452412398369747552|5822555200185981373
M1449|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|1027|Green||2014-05-13|2014-05-15|NaT||||33.7||1|1|2|2|M|Black||11|No|Mother|28031|5|One Parent: Female|Unknown||||Yes||Relative|General Site||Match Support|M|Black||58|28216|Bachelors Degree|Married|Business: Mgt, Admin|27701|30|0|AA Task Force|Special Event|Big|General Site|mentor2.0 2015|Match Support|1|0|0|1|277|60|598|500000170|500015820|503505378|503507249|31|0|1|503796728|31|0|1|500763163|10|1|500000295|2128173570|2|1||-1|500015184|-1|0|3|||11098|8|||1||8034889377453131101|0
M1450|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1044|Green||2014-04-16|2014-04-28|NaT||||34.3||1|1|1|1|M|Black||11|No|Mother|28273|5|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|White||30|28101|Bachelors Degree|Single|Landscaper/Groundskeeper|28269|3|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503446279|503448145|31|0|1|503842555|1|0|1|500759862|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||4208486535559819469|2042734412389339558
M1451|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|92|Green||2016-11-11|2016-12-05|NaT||||3||3|3|1|1|M|Black||11|No|Mother|28262|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||53|28269|Bachelors Degree|Married|Tech: Computer/Programmer|28202|23|0|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|503585510|503587387|31|0|1|504817967|1|0|1|500926954|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1||836952159905822963|5766455966581408090
M1452|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|246|Green||2015-08-11|2015-08-12|2016-04-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.1||3|3|1|1|M|Black||11|No|Mother|28262|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||27|28262|Bachelors Degree|Single|Arts, Entertainment, Sports|28202|0|1|Local TV|Media|Big|General Community|VOL - PreMatch|Match Support|0|1|1|0|277|60|598|500000170|500017732|503585510|503587387|31|0|1|504179374|31|0|1|500835906|10|2|-2||4|1||-2|500007920|-2|0|10|||7438|1|||1||836952159905822963|5766455966581408090
M1453|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|272|Green||2014-10-22|2014-10-22|2015-07-21|Volunteer: Moved|Volunteer: Moved||8.9||2|2|2|2|M|Hispanic||11|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||Relative|General Site||Match Support|M|White||20|28226|Some High School||Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504078916|504080945|3|0|1|503497302|1|0|1|500786376|10|1|500000296|2128173564|4|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1454|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|497|Green||2015-10-09|2015-10-27|NaT||||16.3||2|2|1|1|M|Hispanic||11|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||Relative|General Site||Match Support|M|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504078916|504080945|3|0|1|504311135|1|0|1|500846348|10|1|500000296|2128173564|2|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1455|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1487|Green|Cabarrus County|2013-01-30|2013-02-09|NaT||||48.9||1|1|1|1|M|White||11|No|Mother|28083|3|One Parent: Female|Unknown||||Yes||Self|General Community|Cabarrus County|Match Support|M|White||59|28025|Some College|Married|Business: Sales|28025|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502656083|502656820|1|0|1|503108132|1|0|1|500678455|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|0|0
M1456|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1285|Green||2013-08-27|2013-08-30|NaT||||42.2||1|1|1|1|M|Black||11|Yes|Mother|28217|1|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||28|28209|Bachelors Degree||Finance|28202|2|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500017732|502920379|502921794|31|0|1|503497697|1|0|1|500708164|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||0|0
M1457|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|RTBM|119|Green|Cabarrus County|2016-11-01|2016-11-08|NaT||||3.9||1|1|1|1|F|Black||11|No|Mother|28025|5|One Parent: Female|$35,000 to $39,999||||Yes|BBBS National Site|Web Link|General Community|Cabarrus County|RTBM|F|White||15|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504875300|504877820|31|0|2|504877937|1|0|2|500922404|7|1|500000296|2128173571|2|1|500016374|-2|500016374|-1|34|2|||7464|9|||1|500016374|3575183301237417432|6156547733130613405
M1458|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|403|Green||2016-01-04|2016-01-29|NaT||||13.2||1|1|1|1|F|Hispanic||11|No|Mother|28208|4|Two Parent|Unknown||||Yes||Relative|General Site||Match Support|F|Black||25|28269|Bachelors Degree|Single|Customer Service||0|2|Current/Previous Big|Other Big|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500015820|504531004|504533336|3|0|2|504455232|31|0|2|500870062|10|1|500000295|2128207319|2|1||-1|500007920, 500011315, 500011316|-1|0|3|||17159|12|||1||3935539763241716148|0
M1459|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|544|Green|PERL 2014-2016|2015-08-26|2015-09-10|NaT||||17.9||1|1|1|1|M|Black||11|No|Mother|28203|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28202|Bachelors Degree|Single|Retail: Sales|28209|4|5|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504039192|504041210|31|0|1|504344501|1|0|1|500837420|10|2|-2||2|1|500014681|-2||-2|0|4|||17159|12|||1|500014681|8568001799025358453|7044657180546140448
M1460|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|327|Green||2015-04-29|2015-04-29|2016-03-21|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||10.7||1|1|1|1|F|Black||11|No|Mother|28212|3|One Parent: Female|$25,000 to $29,999||||Yes||School|General Community||Match Support|F|White||26|28205||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500017732|504231007|504233122|31|0|2|504163497|1|0|2|500825416|10|2|-2||4|1||-2||-2|0|4|||17159|12|||1||7554307376683929204|8136849793711030748
M1461|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|322|Green||2016-04-08|2016-04-19|NaT||||10.6||1|1|1|1|M|White||11|No|Mother|28277|4|One Parent: Female|$75,000 to $99,999||||No||School|General Community||Match Support|M|White||53|28270|Masters Degree|Married|Self-Employed, Entrepreneur||15|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504581060|504583394|1|0|1|504503934|1|0|1|500888341|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||0|5081726734274569781
M1462|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|952|Green||2014-06-10|2014-07-29|NaT||||31.3||1|1|1|1|F|Black||11|No|Mother|28226|2|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||46|28207|Bachelors Degree|Married|Arts, Entertainment, Sports|28209|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503867922|503126373|31|0|2|503834583|1|0|2|500766160|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||4903779310522421428|6991424324982091759
M1463|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|647|Green||2014-12-02|2014-12-22|2016-09-29|Volunteer: Time constraint|Volunteer: Time constraint||21.3||1|1|1|1|F|Some Other Race||11|No|Mother|28208|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Enrollment|F|White||24|28209|Bachelors Degree|Single|Business|28207|0|2|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500021785|504004518|504006533|41|0|2|504055712|1|0|2|500800042|5|2|-2||4|1||-2||-2|0|4|||46|2|||1||7581500809034284566|0
M1464|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1206|Red||2012-02-01|2012-03-06|2015-06-25|Volunteer: Moved|Volunteer: Moved||39.6||1|1|1|1|F|Black||11|No|Mother|28205|K|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||26|28269|Some College||Medical|28216|0|3|Recruitment Event|BBBS Board/Staff|Big|General Community|Project Big|Match Support|1|0|1|0|277|60|598|500000170|500008321|502782687|502783868|31|0|2|502760157|31|0|2|500595472|10|2|-2||4|3||-2|500004640|-2|0|10|||7462|13|1207|5|1||5822146217251000296|0
M1465|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|269|Yellow|PERL 2014-2016|2014-09-19|2014-09-29|2015-06-25|Child/Family: Moved|Child/Family: Moved||8.8||1|1|1|1|F|Black||11|No|Mother|28234|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Multi-race (Black & White)||41|28270|Associate Degree|Divorced|Law: Security Officer|28262|1|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500008321|503296668|503298492|31|0|2|503922155|36|0|2|500777025|10|2|-2||4|2|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681|7554307376683929204|34077960614894405
M1466|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|463|Green||2015-11-19|2015-11-30|NaT||||15.2||1|1|1|1|F|Hispanic||11|No|Father|28212|4|Two Parent|$20,000 to $24,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504524360|504526691|3|0|2|504302471|1|0|2|500861415|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1467|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|35|Green||2017-01-10|2017-01-31|NaT||||1.1||2|2|1|1|F|Black||11|No|Mother|28217|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||27|28273|Bachelors Degree|Single|Finance|28202|3|3|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504126227|504128262|31|0|2|504846755|31|0|2|500939318|10|2|-2||2|1|500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||8981704271528751143|2141487034287122220
M1468|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|464|Green||2015-01-09|2015-01-26|2016-05-04|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||15.2||2|2|1|1|F|Black||11|No|Mother|28217|5|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||24|28213||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500021785|504126227|504128262|31|0|2|504042887|31|0|2|500807321|10|2|-2||4|1|500007920, 500011315, 500011316|-2||-2|0|4|||46|2|||1||8981704271528751143|2141487034287122220
M1469|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|561|Red||2014-07-11|2014-07-29|2016-02-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.4||2|2|1|1|F|Black||11|No|Mother|28277|3|One Parent: Female|$30,000 to $34,999|||Y|No||School|General Community||Enrollment|F|Black||31|28270|Bachelors Degree|Single|Business: Sales||0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503388408|503390265|31|0|2|503761210|31|0|2|500769224|5|2|-2||4|3||-2||-2|0|4|||7464|9|||1||5893332617597240023|3318470209175146344
M1470|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|670|Green||2013-05-01|2013-05-16|2015-03-17|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||22||1|1|1|1|M|Black||11|No|Mother|28215||One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|White||29|28208|Bachelors Degree|Single|Law: Police Officer|28216|3|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|502882555|501090456|31|0|1|503438025|1|0|1|500695316|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1||5741767063897867874|4753237757252407321
M1471|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|504|Green||2015-10-09|2015-10-20|NaT||||16.6||1|1|1|1|M|Black||11|No|Mother|28212|4|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|M|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504441613|504443869|31|0|1|504310955|1|0|1|500846394|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1472|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|281|Green||2014-10-10|2014-10-30|2015-08-07|Volunteer: Moved|Volunteer: Moved||9.2||2|2|2|2|F|White||10|No|Mother|28211|1|Two Parent|Unknown||||Yes||School|General Site||RTBM|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503229456|503231244|1|0|2|503603496|1|0|2|500782500|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1473|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1078|Green||2014-03-12|2014-03-25|NaT||||35.4||1|1|1|1|M|Black||10|No|Mother|28227|1|One Parent: Female|$45,000 to $49,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||26|28202|Bachelors Degree|Single|Consultant|28244|2|5|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503411965|503413822|31|0|1|503792970|1|0|1|500754286|10|2|-2||2|1||-2||-2|34|2|||46|2|||1||5388127382485844452|4204211518705620145
M1474|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1249|Green||2013-09-26|2013-10-05|NaT||||41||1|1|1|1|M|Black||10|Yes|Mother|28216|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||27|28203|Bachelors Degree|Single|Real Estate: Realtor|28202|4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|503383959|503554371|31|0|1|503572248|1|0|1|500713580|10|2|-2||2|1|500000294|-2|500000294|-2|0|10|||46|2|||1||3664007741235143067|1698789781793629886
M1475|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|595|Green||2014-10-07|2014-10-21|2016-06-07|Volunteer: Moved|Volunteer: Moved||19.5||2|2|1|1|F|White||10|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049169|504051193|1|0|2|504002563|1|0|2|500781522|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1476|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|F|White||10|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28207|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504049169|504051193|1|0|2|504307866|1|0|2|500929305|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1477|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|541|Red||2015-07-14|2015-07-27|2017-01-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||17.8||1|1|1|1|F|Black||10|No|Mother|28208|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Enrollment|F|Black||24|28262||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|504274120|504276320|31|0|2|504255905|31|0|2|500832878|5|2|-2||4|3||-2||-2|0|4|||17159|12|||1||7284449467126735125|2053394993324953440
M1478|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|155|Green||2016-09-22|2016-10-03|NaT||||5.1||2|2|1|1|M|Multi-race (Black & Hispanic)||10|No|Mother|28036|4|One Parent: Female|$10,000 to $14,999||||Yes||School|General Community||Match Support|M|White||45|28031|Some College|Separated|Business: Sales|27405|10|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment|Match Support|0|1|0|1|277|60|598|500000170|500017732|504658548|504451923|38|0|1|504789938|1|0|1|500909808|10|2|-2||2|1||-2|500007920, 500011316|-2|0|4|||17159|12|||1||0|5081726734274569781
M1479|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|140|Green||2016-04-01|2016-04-11|2016-08-29|Child: Changed school/site|Child: Changed school/site||4.6||2|2|2|2|M|Multi-race (Black & Hispanic)||10|No|Mother|28036|4|One Parent: Female|$10,000 to $14,999||||Yes||School|General Community||Match Support|M|Black||21|28035|Some College|Single|Student: College||0|0|Self|Self|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504658548|504451923|38|0|1|504629735|31|0|1|500887477|10|1|500000295|2128173570|4|1||-2||-1|0|4|||7464|9|||1||0|5081726734274569781
M1480|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|274|Green||2014-10-04|2014-11-06|2015-08-07|Volunteer: Moved|Volunteer: Moved||9||3|3|2|2|F|Hispanic||10|No|Mother|28105|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503206081|503663066|3|0|2|503497526|1|0|2|500780604|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1481|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|348|Green||2015-10-09|2015-10-21|2016-10-03|Child: Changed school/site|Child: Changed school/site||11.4||3|3|2|2|F|Hispanic||10|No|Mother|28105|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||18|28227|Some High School|Single|Student: College||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500022905|503206081|503663066|3|0|2|504296357|1|0|2|500846341|10|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1482|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|489|Green|PERL 2014-2016, Cabarrus County|2015-10-27|2015-11-04|NaT||||16.1||1|1|1|1|F|Multi-race (Hispanic & Asian)||10|No|Mother|28081|5|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||40|28025||Married|Self-Employed, Entrepreneur||11|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504432726|504434981|40|0|2|504430061|1|0|2|500852606|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7464|9|||1|500014681, 500016374|2437132833506538679|3993797463174785246
M1483|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1785|Green|Amachi|2012-04-05|2012-04-17|NaT||||58.6||1|1|1|1|F|Black||10|No|Mother|28206|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|F|White||28|28208|Bachelors Degree|Single|Business: Marketing|28269|0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502869627|502871029|31|0|2|502932955|1|0|2|500608271|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|500000294|392688197545050058|2053394993324953440
M1484|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|381|Green||2015-05-03|2015-05-04|2016-05-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.5||2|2|1|1|M|Black||10|Yes|Mother|28213|3|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||31|28105|Bachelors Degree|Married|Consultant|43215|1|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504240016|504242131|31|0|1|504155486|1|0|1|500825676|10|2|-2||4|1|500000294|-2||-2|0|10|||17159|12|||1||6065435025527210335|3326174373441625173
M1485|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|42|Green||2017-01-10|2017-01-24|NaT||||1.4||2|2|1|1|M|Black||10|Yes|Mother|28213|3|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|Black||29|28211|Bachelors Degree|Single|Business: Engineer|28212|3|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504240016|504242131|31|0|1|504911868|31|0|1|500939329|10|2|-2||2|1|500000294|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||6065435025527210335|3326174373441625173
M1486|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1079|Yellow||2013-02-13|2013-02-26|2016-02-10|Child: Lost interest|Child: Lost interest||35.4||1|1|1|1|F|White||10|No|Mother|28226|1|One Parent: Female|$25,000 to $29,999||||No||School|General Community||Match Support|F|White||27|28207|Bachelors Degree|Single|Arts, Entertainment, Sports|28207|0|0|Billboard|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503297711|503299535|1|0|2|503353908|1|0|2|500681652|10|2|-2||4|2||-2||-2|0|4|||125|1|||1||4902029756574603597|866643722990487659
M1487|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|519|Green||2015-09-28|2015-10-05|NaT||||17.1||1|1|1|1|M|Black||10|No|Mother|28213|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Consultant|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504179804|504181918|31|0|1|504337207|1|0|1|500842586|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||9080589164524051479|7044657180546140448
M1488|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|811|Green||2014-12-02|2014-12-17|NaT||||26.6||1|1|1|1|M|Black||10|No|Mother|28208|3|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||29|28203|Masters Degree|Married|Business|28202|0|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|504058316|504060340|31|0|1|503984749|1|0|1|500800274|10|2|-2||2|1||-2||-2|34|2|||7462|13|||1||6065435025527210335|8456769937733544110
M1489|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|418|Green|PERL 2014-2016|2016-01-04|2016-01-14|NaT||||13.7||1|1|1|1|F|Black||10|No|Mother|28203|3|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||25|28209|Bachelors Degree|Single|Business|28277|1|0|Bowl For Kids Sake|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504388295|504390534|31|0|2|504404378|1|0|2|500870013|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||132|8|||1|500014681|7284449467126735125|2141487034287122220
M1490|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|567|Red||2015-03-08|2015-04-13|2016-10-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.6||1|1|1|1|M|Black||10|No|Mother|28212|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Business|33701|2|11|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|504122670|504124721|31|0|1|504179830|1|0|1|500817495|10|2|-2||4|3||-2||-2|0|4|||46|2|||1||5386346637278076349|0
M1491|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|841|Green||2014-11-10|2014-11-17|NaT||||27.6||1|1|1|1|M|Black||10|No|Mother|28105|2|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|White||44|28211|Bachelors Degree|Married|Business: Human Resources|28255|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|504030099|504032117|31|0|1|503994598|1|0|1|500793822|10|2|-2||2|1||-2||-2|0|4|||7671|13|||1||7134583514356134698|0
M1492|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|292|Green||2014-12-01|2015-01-15|2015-11-03|Volunteer: Time constraint|Volunteer: Time constraint||9.6||1|1|2|2|M|Black||10|No|Mother|28206|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||27|28262|Associate Degree|Divorced|Medical: Nurse|28203|1|0|Self|Self|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500016270|504005675|504007690|31|0|1|502635965|31|0|1|500799927|10|1|500000295|2128173561|4|1||-1||-1|0|4|||7464|9|||1||7960300212314874874|0
M1493|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|138|Green|PERL 2014-2016|2016-09-13|2016-10-20|NaT||||4.5||1|1|1|1|M|Black||10|No|Mother|28216|4|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28203|Bachelors Degree|Single|Finance: Banking|28281|3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504647175|504649586|31|0|1|504759286|1|0|1|500907299|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||17159|12|||1|500014681|2324686837245224089|7044657180546140448
M1494|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1245|Green|Cabarrus County|2013-09-19|2013-10-09|NaT||||40.9||1|1|1|1|M|Black||10|Yes|Mother|28083|K|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||33|28269|Bachelors Degree|Single|Retail: Sales|28027|0|6|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502776079|502777258|31|0|1|503573272|1|0|1|500711993|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|370020301266015142|0
M1495|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|569|Green||2014-12-03|2014-12-03|2016-06-24|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||18.7||1|1|1|1|F|White||10|No|Father|28083||Other Relative|Unknown||||Yes||School|General Site|Cabarrus County|Enrollment|F|White||66|28025||Married|Retired||0|0|Bowl For Kids Sake|Special Event|Big|General Site|Cabarrus County|Enrollment|1|0|1|0|277|60|598|500000170|500012459|504073587|504075616|1|0|2|503904297|1|0|2|500800825|5|1|500000295|2128212919|4|1|500016374|-1|500016374|-1|0|4|||132|8|||1||2437132833506538679|0
M1496|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|167|Green|Cabarrus County|2016-03-29|2016-04-15|2016-09-29|Child/Family: Moved|Child/Family: Moved||5.5||1|1|1|1|F|Black||10|No|Mother|28025|4|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Site|Cabarrus County|Match Support|F|White||18|28081|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504666129|504668556|31|0|2|504583619|1|0|2|500886774|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|3|||7464|9|||1|500016374|3324851395989241799|0
M1497|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|118|Green|Cabarrus County|2016-11-01|2016-11-09|NaT||||3.9||1|1|1|1|F|White||10|No|Mother|28027|4|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|Cabarrus County|Match Support|F|White||17|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504907815|504910335|1|0|2|504878315|1|0|2|500922402|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|3232906304025417619|7335049822486282493
M1498|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|738|Green||2015-02-09|2015-02-28|NaT||||24.2||3|3|1|1|F|Black||10|Yes|Aunt|28227|3|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||69|28104||Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502643841|502255582|31|0|2|504076732|1|0|2|500812797|10|2|-2||2|1|500000294|-2||-2|0|10|||46|2|||1||2056258660718146620|0
M1499|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|102|Green||2014-10-15|2014-10-20|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||3.4||3|3|1|1|F|Black||10|Yes|Aunt|28227|3|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||53|28215||Married|Unemployed||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|502643841|502255582|31|0|2|503991357|31|0|2|500783837|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1||2056258660718146620|0
M1500|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|353|Green||2014-10-21|2014-10-21|2015-10-09|Child: Changed school/site|Child: Changed school/site||11.6||1|1|2|2|F|Black||10|No|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||Relative|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504078931|504080960|31|0|2|503905510|1|0|2|500785765|10|1|500000296|2128173564|4|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1501|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|111|Green||2016-10-24|2016-11-16|NaT||||3.6||1|1|1|1|F|Black||10|No|Mother|28211|5|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||39|28277|Masters Degree|Married|Education||3|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504835647|504838149|31|0|2|504545759|31|0|2|500918758|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1||6627885846854295604|8726431331992650796
M1502|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|16|Green|Cabarrus County|2017-02-09|2017-02-19|NaT||||0.5||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28027|5|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|Black||54|28075|Masters Degree|Married|Business||0|9|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504819474|504821973|36|0|1|505001672|31|0|1|500945474|10|2|500016307||2|1||-2|500016374|-2|0|10|||7464|9|||1|500016374|1550830965009450729|0
M1503|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|417|Green||2013-11-18|2014-01-06|2015-02-27|Child: Graduated|Child: Graduated||13.7||1|1|2|2|F|Hispanic||10|No|Mother|28209|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Asian||49|28210|Masters Degree|Married|Education: Teacher||0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|1|0|1|0|277|60|598|500000170|500008321|503718011|503719978|3|0|2|503281135|4|0|2|500732119|10|1|-1||4|1||-1|500015184|-1|0|4|||7462|13|||1||8568001799025358453|0
M1504|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|943|Green||2013-06-25|2013-07-03|2016-02-01|Volunteer: Moved|Volunteer: Moved||31||1|1|1|1|F|Black||10|No|Mother|28211||One Parent: Female|Unknown|||Y|Yes||Self|General Community||Enrollment|F|Black||46|28256|Associate Degree|Single|Finance: Banking||7|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|502610111|501288299|31|0|2|501041084|31|0|2|500701839|5|2|-2||4|1||-2||-2|0|10|||46|2|||1||1158671944891395407|0
M1505|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|645|Green||2014-04-07|2014-05-20|2016-02-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.2||2|2|1|1|F|Multi-race (Black & White)||10|No|Mother|28115|3|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|White||46|28211|Bachelors Degree|Married|Finance|28105|11|4|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500018851|503076808|503078467|36|0|2|503688665|1|0|2|500758530|10|2|-2||4|1||-2|500000294|-2|0|10|||46|2|||1||7857548027029642592|8690133977366715726
M1506|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1407|Green||2013-04-30|2013-04-30|NaT||||46.2||1|1|1|1|F|Black||10|No|Mother|28278|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||29|28205|Masters Degree|Single|Finance|28203|0|6|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020752|503389942|503239061|31|0|2|503191064|1|0|2|500695067|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||8050480174690503915|7044657180546140448
M1507|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|504|Green||2015-10-09|2015-10-20|NaT||||16.6||1|1|1|1|F|Hispanic||10|No|Mother|28212|4|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504442301|504444557|3|0|2|504296402|1|0|2|500846393|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1508|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|265|Yellow||2016-01-07|2016-01-08|2016-09-29|Child/Family: Moved|Child/Family: Moved||8.7||1|1|2|3|F|Black||10|No|Mother|28083||One Parent: Female|$30,000 to $34,999||||Yes||School|General Site|Cabarrus County|Match Support|F|Black||28|28083|Bachelors Degree|Single|Law|28147|0|2|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504530688|504533020|31|0|2|504528677|31|0|2|500870768|10|1|500000295|2128232374|4|2|500016374|-1|500016374|-2|0|4|||7496|10|||1||2043334928777030191|0
M1509|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|482|Green||2015-10-21|2015-11-11|NaT||||15.8||1|1|1|1|M|Black||10|Yes|Mother|28216|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community|Amachi|Match Support|M|Black||41|28214|Some College|Married|Business|28287|0|3|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504207638|504209750|31|0|1|504357457|31|0|1|500850393|10|2|-2||2|1|500000294|-2||-2|0|4|||17159|12|||1||2979941694006626856|7674215580094440446
M1510|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|119|Green||2014-09-30|2014-10-06|2015-02-02|Child/Family: Moved|Child/Family: Moved||3.9||1|1|2|2|M|Black||10|Yes|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500019116|504041737|504043755|31|0|1|503901650|1|0|1|500779466|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1511|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2017-01-10|2017-01-30|NaT||||1.2||1|1|1|1|F|Multi-race (Black & White)||10|No|Mother|28213|5|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||38|28202|Bachelors Degree|Single|Business|28202|0|2|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504888357|504890877|36|0|2|504850919|1|0|2|500939317|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1||836952159905822963|4855845956679832355
M1512|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|494|Green||2015-10-08|2015-10-30|NaT||||16.2||1|1|1|1|F|Black||10|No|Mother|28216|4|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|F|Black||31|28216|Bachelors Degree|Single|Arts, Entertainment, Sports|28202|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504345626|504347850|31|0|2|504373316|31|0|2|500845709|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||7679812394383646966|1712849328738258411
M1513|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|42|Green||2017-01-18|2017-01-24|NaT||||1.4||1|1|1|1|M|Hispanic||10|No|Mother|28027|4|Two Parent|Unknown||||Yes||School|General Site|Cabarrus County|Match Support|M|White||76|28075||Married|Business||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504975900|504978451|3|0|1|504998038|1|0|1|500940723|10|1|500000295|2128212924|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||3232906304025417619|0
M1514|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|98|Green||2016-11-18|2016-11-29|NaT||||3.2||1|1|2|2|M|Hispanic||10|No|Mother|28211|5|Two Parent|$15,000 to $19,999||||Yes||School|General Site||Match Support|M|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504932738|504935289|3|0|1|504307950|1|0|1|500929299|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1515|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|779|Green|PERL 2014-2016|2015-01-08|2015-01-18|NaT||||25.6||1|1|1|1|F|Black||10|Yes|Mother|28208|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||27|29730|Bachelors Degree|Married|Finance|28277|3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504115691|504117725|31|0|2|504068384|1|0|2|500807126|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681|7857548027029642592|0
M1516|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1327|Green||2013-07-09|2013-07-19|NaT||||43.6||1|1|1|1|F|Hispanic||10|No|Mother|28217|1|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||35|28273|Masters Degree|Single|Finance: Accountant|28201|9|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020753|503355399|503348836|3|0|2|503428702|1|0|1|500703056|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||0|0
M1517|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|372|Green||2014-06-23|2014-07-16|2015-07-23|Volunteer: Health|Volunteer: Health||12.2||3|3|1|1|F|Black||10|No|GrandMother|28083|1|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||37|28027|Some College|Married|Business: Mgt, Admin|28255|2|6|Local Print|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503585540|503587420|31|0|2|503798839|1|0|2|500767384|10|2|-2||4|1|500014681|-2||-2|34|2|||7439|1|||1||6810228174639243761|0
M1518|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|140|Red|PERL 2014-2016|2015-10-07|2015-10-26|2016-03-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.6||3|3|1|1|F|Black||10|No|GrandMother|28083|1|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||22|28081||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500020753|503585540|503587420|31|0|2|504301494|1|0|2|500845172|10|2|-2||4|3|500014681|-2||-2|34|2|||17159|12|||1|500014681|6810228174639243761|0
M1519|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|601|Green||2014-10-07|2014-10-21|2016-06-13|Volunteer: Moved|Volunteer: Moved||19.7||1|1|1|1|F|Black||10|Yes|Mother|28105|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504050657|504052681|31|0|2|503929917|1|0|2|500781524|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||0|0
M1520|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|858|Green||2014-10-29|2014-10-31|NaT||||28.2||1|1|1|1|M|Black||10|No|Mother|28208|5|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|M|White||40|28204|Bachelors Degree|Single|Business|28027|8|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503931637|503933644|31|0|1|504068281|1|0|1|500789322|10|2|-2||2|1||-2||-2|0|4|||46|2|||1||7089569121628268952|8626610080771140821
M1521|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|88|Green||2016-12-06|2016-12-09|NaT||||2.9||1|1|1|1|M|Black||10|No|Mother|28031|5|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|M|White||20|28035||Single|Education|20901|12|6|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504848419|504850921|31|0|1|504941003|1|0|1|500933672|10|1|500000295|2128173570|2|1||-1||-1|0|4|||7464|9|||1||8034889377453131101|0
M1522|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|448|Green||2015-11-23|2015-12-15|NaT||||14.7||1|1|1|1|M|Black||10|Yes|Mother|28217|5|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|M|White||69|28277|Masters Degree|Widowed|Retired||0|0|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504517631|504519932|31|0|1|504284567|1|0|1|500862686|10|1|500000295|2128173557|2|1|500007920, 500011315, 500011316|-1||-1|0|4|||17159|12|||1||8981704271528751143|0
M1523|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1421|Green||2013-04-02|2013-04-16|NaT||||46.7||1|1|1|1|F|Black||10|Yes|Mother|28212|1|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||29|28202|Bachelors Degree|Single|Business|28226|1|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503246892|503248691|31|0|2|503350295|1|0|2|500691065|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1||2762897743412756173|0
M1524|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1301|Yellow||2012-06-15|2012-06-21|2016-01-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||42.7||2|2|1|1|F|Black||10|No|Mother|28215|1|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||37|28270|Bachelors Degree|Single|Finance: Banking||0|0|Recruitment Event|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500013781|502688939|501750989|31|0|2|503023856|1|0|2|500619498|10|2|-2||4|2||-2||-2|0|10|||7458|9|||1||8568001799025358453|0
M1525|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|658|Green|PERL 2014-2016|2015-04-29|2015-05-19|NaT||||21.6||1|1|1|1|F|White||10|No|GrandMother|28210|3|Other Relative|Unknown||||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||28|28205|Some College|Single|Transport: Driver|28277|8|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|504234369|503470938|1|0|2|504116244|35|0|2|500825294|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||46|2|||1|500014681|6898335769881586649|7044657180546140448
M1526|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|196|Green||2016-08-16|2016-08-23|NaT||||6.4||1|1|1|1|M|Black||10|No|Mother|28277|3|One Parent: Female|$40,000 to $44,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||45|28210|Masters Degree|Divorced|Finance: Banking|28202|10|11|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504022991|504025006|31|0|1|504545438|31|0|1|500903682|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1||5893332617597240023|5969614404793803539
M1527|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|770|Green||2015-01-14|2015-01-27|NaT||||25.3||1|1|1|1|M|Black||10|No|Mother|28262|4|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Tech: Engineer|28027|3|11|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020752|503801691|503803668|31|0|1|504142324|1|0|1|500808169|10|2|-2||2|1||-2|500000294|-2|0|10|||17159|12|||1||7127394271070859649|386356889061704511
M1528|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1226|Green||2013-06-27|2013-07-10|2016-11-17|Volunteer: Time constraint|Volunteer: Time constraint||40.3|Y|2|2|1|1|M|Black||10|No|Mother|28269|5|One Parent: Female|$40,000 to $44,999||||No||School|General Community||Match Support|M|White||34|28078|Bachelors Degree|Married|Business: Mgt, Admin|28262|2|10|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017732|502543702|502544155|31|0|1|503346987|1|0|1|500702244|10|2|-2||4|1||-2|500000294|-2|0|4|||7464|9|||1||0|6418092831698127977
M1529|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|15|Green||2017-01-23|2017-02-20|NaT||||0.5||2|2|1|1|M|Black||10|No|Mother|28269|5|One Parent: Female|$40,000 to $44,999||||No||School|General Community||Match Support|M|White||23|28269|Bachelors Degree|Single|Business: Engineer|28104|1|5|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|502543702|502544155|31|0|1|504874916|1|0|1|500941320|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||0|6418092831698127977
M1530|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2015|Green||2011-08-12|2011-08-31|NaT||||66.2||1|1|1|1|F|Black||10|No|Mother|28269|2|One Parent: Female|$40,000 to $44,999||||No||School|General Community||Match Support|F|White||29|28202|Bachelors Degree|Single|Service: Hotel||0|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|502544010|502544463|31|0|2|502641777|1|0|2|500549950|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||0|5468286809853673926
M1531|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|250|Green|Cabarrus County|2016-06-20|2016-06-30|NaT||||8.2||1|1|1|1|M|Multi-race (Hispanic & White)||10|No|Mother|28025|3|One Parent: Female|Unknown|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28027|Bachelors Degree|Single|Business|28027|2|4|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504553935|504556269|35|0|1|504682974|1|0|1|500897234|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|34|2|||7464|9|||1|500016374|3380316005507597709|8216069172157856234
M1532|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|609|Green||2014-10-04|2014-10-06|2016-06-06|Volunteer: Moved|Volunteer: Moved||20||2|2|1|1|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504041835|504043867|3|0|1|503895081|1|0|1|500780581|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1533|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28277|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504041835|504043867|3|0|1|504303741|1|0|1|500929317|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1534|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|287|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-04-19|2016-05-24|NaT||||9.4||1|1|1|1|F|Black||10|No|Mother|28208|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||29|28210|Bachelors Degree|Single|Business: Sales|28269|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504556546|504558880|31|0|2|504283498|1|0|2|500889681|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1|500007920, 500011315, 500011316|5473689050106799364|6084148439133243542
M1535|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|419|Green||2015-06-24|2015-06-30|2016-08-22|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||13.8||1|1|2|2|M|White||10|No|Mother|28277|3|One Parent: Female|$40,000 to $44,999|||Y|Yes||Self|General Community||Match Support|M|White||57|28105|Bachelors Degree|Married|Business: Sales|28203|11|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|503921502|503891297|1|0|1|504063702|1|0|1|500831159|10|2|-2||4|1||-2|500000294|-2|0|10|||17159|12|||1||7444351539618566014|6156547733130613405
M1536|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|665|Green||2015-04-15|2015-05-12|NaT||||21.8||1|1|1|1|F|White||10|No|Mother|28277|4|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|F|White||29|29708|Bachelors Degree|Married|Medical|28105|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503889301|503891297|1|0|2|504021478|1|0|2|500823483|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||7444351539618566014|6156547733130613405
M1537|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green||2016-11-18|2016-12-05|NaT||||3||2|2|2|2|M|Hispanic||10|No|Father|28211|3|Two Parent|Unknown||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|Asian||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504495775|504498060|3|0|1|504376009|4|0|1|500929354|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M1538|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|328|Green||2015-11-01|2015-11-11|2016-10-04|Child: Changed school/site|Child: Changed school/site||10.8||2|2|2|2|M|Hispanic||10|No|Father|28211|3|Two Parent|Unknown||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|Asian||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504495775|504498060|3|0|1|504376009|4|0|1|500854809|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M1539|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|313|Green|PERL 2014-2016, Cabarrus County|2016-04-07|2016-04-28|NaT||||10.3||1|1|1|1|M|White||10|No|GrandMother|28124|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||35|28027|Bachelors Degree|Single|Tech: Computer/Programmer|28202|2|6|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, mentor2.0, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504640447|504638197|1|0|1|504266263|1|0|1|500888255|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014505, 500016374|-2|0|4|||17159|12|||1|500014681, 500016374|1345826867198613426|0
M1540|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|741|Green||2015-02-25|2015-02-25|NaT||||24.3||2|2|1|1|M|Hispanic||10|Yes|Mother|28031|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||21|28035||Single|Student: College||0|0|Kappa Alpha Psi|Fraternity/Sorority|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|503720519|503722491|3|0|1|504207546|1|0|1|500815623|10|1|500000295|2128173570|2|1||-1||-1|0|4|||8693|14|||1||8034889377453131101|0
M1541|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|357|Green||2014-10-04|2014-10-14|2015-10-06|Child: Changed school/site|Child: Changed school/site||11.7||2|2|1|1|M|Black||10|Yes|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site|Amachi|Match Support|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503281864|503263744|31|0|1|503897642|1|0|1|500780592|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1542|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1286|Green||2013-08-13|2013-08-29|NaT||||42.3||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28212|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||28|28207|PHD|Married|Medical: Healthcare Worker|28025|2|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503569406|503567063|38|0|2|503534366|1|0|2|500706542|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||7127394271070859649|0
M1543|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|117|Green|Cabarrus County|2016-11-07|2016-11-10|NaT||||3.8||1|1|1|1|F|Black||10|No|Mother|28081|5|One Parent: Female|Unknown||||No||School|General Site|Cabarrus County|Match Support|F|White||17|28269||Single|Student: High School||0|0|Other|BBBS Board/Staff|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504918317|504920837|31|0|2|504932049|1|0|2|500925583|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7671|13|||1|500016374|0|0
M1544|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1042|Green||2014-04-14|2014-04-30|NaT||||34.2||1|1|1|1|M|Black||10|No|Mother|28214|5|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||45|28214|Masters Degree|Married|Business|28207|3|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502931159|502932575|31|0|1|503802032|1|0|1|500759587|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||8452412398369747552|0
M1545|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1329|Green||2013-06-10|2013-07-17|NaT||||43.7||1|1|1|1|M|Black||10|No|Mother|28215|1|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|M|White||30|28203|Bachelors Degree|Single|Finance|28202|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503402178|503404035|31|0|1|503468005|1|0|1|500700142|10|2|-2||2|1||-2||-2|0|3|||7496|10|||1||314687390558932914|7044657180546140448
M1546|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|720|Red||2013-09-18|2013-09-26|2015-09-16|Child: Lost interest|Child: Lost interest||23.7||1|1|1|1|F|Black||10|No|Mother|28212|2|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||Match Support|F|Black||38|28262|Masters Degree|Divorced|Finance|28202|3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503586001|503587878|31|0|2|503568168|31|0|2|500711704|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||5822146217251000296|5304581627889532800
M1547|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|720|Red||2013-09-18|2013-09-26|2015-09-16|Child: Lost interest|Child: Lost interest||23.7||1|1|1|1|F|Black||10|No|Mother|28212|2|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|F|Black||47|28269|Bachelors Degree|Married|Medical: Nurse|28078|8|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503586069|503587878|31|0|2|503541572|31|0|2|500711744|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1||5822146217251000296|5304581627889532800
M1548|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|426|Red|PERL 2014-2016|2015-02-10|2015-02-17|2016-04-18|Volunteer: Moved|Volunteer: Moved||14||1|1|1|1|F|White||10|No|Mother|28078|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community|PERL 2014-2016|Enrollment|F|White||38|28031|Some College|Single|Real Estate: Realtor|28031|8|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500008321|504134912|504136949|1|0|2|503909509|1|0|2|500813035|5|2|-2||4|3|500014681|-2|500014681|-2|0|4|||46|2|||1|500014681|7777315526213898088|0
M1549|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|81|Green||2016-12-16|2016-12-16|NaT||||2.7||1|1|2|2|F|Black||10|No|Mother|29715|6|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|Black||31|28216|Masters Degree|Single|Customer Service|28217|1|6|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500013781|504970032|504972583|31|0|2|504037091|31|0|2|500936280|10|1|500009132|2128233620|2|1||-1||-1|0|4|||11247|3|||1||1174067921639243853|0
M1550|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|574|Green||2014-11-11|2014-11-11|2016-06-07|Volunteer: Moved|Volunteer: Moved||18.9||2|2|2|2|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504095778|504178353|3|0|1|503916388|1|0|1|500794487|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||0|0
M1551|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28211|Some College|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504095778|504178353|3|0|1|504307795|1|0|1|500929326|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||0|0
M1552|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|503|Green||2015-01-21|2015-01-21|2016-06-07|Volunteer: Moved|Volunteer: Moved||16.5||2|2|2|2|M|Hispanic||10|No|Mother|28212||One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504176244|504178353|3|0|1|503901671|1|0|1|500809239|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1553|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|M|Hispanic||10|No|Mother|28212||One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28203|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504176244|504178353|3|0|1|504324165|1|0|1|500929314|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1554|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|31|Green|Cabarrus County|2017-01-27|2017-02-04|NaT||||1||1|1|1|1|M|Black||10|No|Mother|28027|5|One Parent: Female|$15,000 to $19,999||||Yes||School|General Community|Cabarrus County|Match Support|M|Black||34|28227|Juris Doctorate (JD)|Separated|Law: Lawyer|28227|9|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504937135|504939686|31|0|1|504694440|31|0|1|500942634|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|500016374|1550830965009450729|0
M1555|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|531|Green|PERL 2014-2016|2015-09-10|2015-09-23|NaT||||17.4||2|2|1|1|M|Black||10|No|Mother|28214|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||25|28227|Bachelors Degree|Single|Insurance|28277|1|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503779386|503781363|31|0|1|504333970|31|0|1|500839160|10|2|-2||2|1|500014681|-2||-2|0|4|||7464|9|||1|500014681|7554307376683929204|1546374315672654438
M1556|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|494|Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2015-10-08|2015-10-30|NaT||||16.2|Y|1|1|1|1|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28204|Masters Degree|Married|Consultant||0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|504254978|504257111|3|0|1|504379733|1|0|1|500845639|10|2|-2||2|1|500014681|-2|500014681|-2|0|5|||46|2|||1|500011312, 500014681|9080589164524051479|0
M1557|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|139|Green||2016-10-02|2016-10-19|NaT||||4.6||1|1|3|3|F|Black||10|No|Mother|28208|6|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|Black||30|28270|Masters Degree|Single|Finance|28202|0|1|Duke Energy|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504875019|504877539|31|0|2|504396349|31|0|2|500911911|10|1|500009132|2128207318|2|1||-1||-1|0|4|||16705|3|||1||2611337051335117774|0
M1558|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|350|Green|Cabarrus County|2016-02-29|2016-03-22|NaT||||11.5||1|1|1|1|F|Black||10|No|Mother|28025|4|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|Cabarrus County|Match Support|F|Black||18|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504605286|504607697|31|0|2|504579876|31|0|2|500882081|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|3324851395989241799|0
M1559|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|98|Green||2014-10-04|2014-10-17|2015-01-23|Volunteer: Time constraint|Volunteer: Time constraint||3.2||3|3|2|2|M|Hispanic||10|No|Mother|28212|1|One Parent: Female|Unknown||||No||School|General Site||Match Support|M|White||19|28205|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503214548|503216323|3|0|1|503500393|1|0|1|500780601|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1560|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|232|Green||2015-02-02|2015-02-09|2015-09-29|Child: Changed school/site|Child: Changed school/site||7.6||3|3|2|2|M|Hispanic||10|No|Mother|28212|1|One Parent: Female|Unknown||||No||School|General Site||Match Support|M|White||19|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503214548|503216323|3|0|1|503901650|1|0|1|500811548|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1561|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|105|Green||2016-11-22|2016-11-22|NaT||||3.4||1|1|2|2|F|White||10|No|Mother|28212|5|Two Parent|$30,000 to $34,999||||No||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504896389|504898909|1|0|2|504301129|1|0|2|500930399|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1562|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|869|Green||2014-10-09|2014-10-20|NaT||||28.6||1|1|1|1|M|Black||10|No|Mother|28031|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||21|28031|Some College|Single|Student: College||0|0|Kappa Alpha Psi|Fraternity/Sorority|Big|General Site||Match Support|1|0|0|1|277|60|598|500000170|500015820|503630433|503632372|31|0|1|504025162|31|0|1|500782178|10|1|500000295|2128173570|2|1||-1||-1|0|4|||8693|14|||1||8034889377453131101|0
M1563|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|366|Green||2015-05-19|2015-05-19|2016-05-19|Volunteer: Time constraint|Volunteer: Time constraint||12||1|1|1|1|F|Black||10|No|Mother|28212|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community|Amachi|Enrollment|F|White||31|28031|Associate Degree|Married|Business: Marketing||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500018851|504205503|504207614|31|0|2|504191463|1|0|2|500827528|5|2|-2||4|1|500000294|-2|500000294|-2|0|4|||7438|1|||1||392688197545050058|7500593753197857009
M1564|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|470|Green|PERL 2014-2016|2015-11-06|2015-11-23|NaT||||15.4||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28208|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||30|28204|Some College|Single|Medical|28208|3|3|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504278828|504281028|38|0|2|504354967|35|0|2|500857068|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500014681|967246839551912690|2378213070582218846
M1565|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|62|Green||2017-01-02|2017-01-04|NaT||||2||1|1|1|1|F|Hispanic||10|No|Mother|28212|5|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||19|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504976138|504978689|3|0|2|504709284|1|0|2|500937876|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1566|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|7|Green||2017-02-10|2017-02-28|NaT||||0.2||1|1|1|1|M|Black||10|No|Mother|28277|5|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|M|White||31|28277|Masters Degree|Married|Finance: Accountant|28273|0|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504838542|504838321|31|0|1|504930064|1|0|1|500945724|10|2|-2||2|1|500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||1078778250813636816|2742327884002010428
M1567|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|88|Green||2016-12-05|2016-12-09|NaT||||2.9||1|1|1|1|M|White||10|No|Mother|28031|5|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Site||Match Support|M|White||36|28036|Masters Degree|Married|Finance: Banking|28210|6|0|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504951152|504953703|1|0|1|504775091|1|0|1|500933275|10|1|500000295|2128173570|2|1||-1||-1|0|3|||17159|12|||1||8034889377453131101|0
M1568|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|111|Green|PERL 2014-2016, Cabarrus County|2016-11-15|2016-11-16|NaT||||3.6||1|1|1|1|M|White||10|No|Mother|28081|5|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||25|28027||Married|Medical: Healthcare Worker||0|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|504862022|504864541|1|0|1|504930361|1|0|1|500927996|10|2|-2||2|1|500014681, 500016374|-2|500014681, 500016374|-2|34|2|||7671|13|||1|500014681, 500016374|6810228174639243761|2036270106764562772
M1569|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|155|Green||2016-09-07|2016-10-03|NaT||||5.1||1|1|1|1|M|Black||10|No|GrandMother|28212|4|One Parent: Female|$10,000 to $14,999|||Y|No||School|General Community|PERL 2014-2016|Match Support|M|White||48|28211|Masters Degree|Married|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504592676|504595050|31|0|1|504742988|1|0|1|500906468|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1||0|0
M1570|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|321|Green|PERL 2014-2016|2015-10-27|2015-11-13|2016-09-29|Volunteer: Time constraint|Volunteer: Time constraint||10.5||2|2|2|2|F|Black||10|Yes|Mother|28027|4|Other/Unknown|Unknown||||Yes||School|General Site|Amachi, Cabarrus County, PERL 2014-2016|Enrollment|F|White||31|28025||Married|Retail: Mgt|28025|5|0|Recruitment Event|Workplace Partner|Big|General Site|Cabarrus County, PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500012459|504137677|504139717|31|0|2|504026893|1|0|2|500852587|5|1|500000295|2128212924|4|1|500000294, 500014681, 500016374|-1|500014681, 500016374|-1|0|4|||7446|3|||1|500014681|3232906304025417619|0
M1571|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Enrollment|294|Yellow||2014-12-03|2014-12-11|2015-10-01|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||9.7||2|2|1|1|F|Black||10|Yes|Mother|28027|4|Other/Unknown|Unknown||||Yes||School|General Site|Amachi, Cabarrus County, PERL 2014-2016|Enrollment|F|Black||29|28025||Living w/ Significant Other|Retail: Sales|28027|0|0|Recruitment Event|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500012459|504137677|504139717|31|0|2|504032683|31|0|2|500801052|5|1|500000295|2128212924|4|2|500000294, 500014681, 500016374|-1||-1|0|4|||7446|3|||1||3232906304025417619|0
M1572|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|318|Green||2014-09-21|2014-09-23|2015-08-07|Volunteer: Moved|Volunteer: Moved||10.4||3|3|2|2|F|Black||10|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503315297|503317130|31|0|2|503507566|1|0|2|500777108|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1573|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|83|Green||2015-10-09|2015-10-15|2016-01-06|Child/Family: Moved|Child/Family: Moved||2.7||3|3|2|2|F|Black||10|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503315297|503317130|31|0|2|504308458|1|0|2|500846385|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1574|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|607|Green||2014-10-04|2014-10-08|2016-06-06|Volunteer: Moved|Volunteer: Moved||19.9||2|2|1|1|F|Black||10|No|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049186|504065687|31|0|2|503898609|1|0|2|500780590|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1575|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-18|2016-11-30|NaT||||3.2||2|2|2|2|F|Black||10|No|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||18|28227|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504049186|504065687|31|0|2|504302535|31|0|2|500929350|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1576|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|279|Green||2014-10-10|2014-10-14|2015-07-20|Volunteer: Moved|Volunteer: Moved||9.2||3|3|2|2|F|Black||10|Yes|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504063660|504065687|31|0|2|503507139|1|0|2|500782501|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1577|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||3|3|2|2|F|Black||10|Yes|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504063660|504065687|31|0|2|504307828|1|0|2|500929288|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1578|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|395|Green||2015-10-09|2015-10-16|2016-11-14|Volunteer: Time constraint|Volunteer: Time constraint||13||3|3|1|1|F|Black||10|Yes|Mother|28211|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28203|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504063660|504065687|31|0|2|504306023|1|0|2|500846383|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1579|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|616|Green||2014-09-29|2014-09-30|2016-06-07|Volunteer: Moved|Volunteer: Moved||20.2||3|3|1|1|M|Hispanic||10|No|Mother|28211|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020909|503229418|503231198|3|0|1|503907312|1|0|1|500778740|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1580|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||3|3|2|2|M|Hispanic||10|No|Mother|28211|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|503229418|503231198|3|0|1|504310910|1|0|1|500928398|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1581|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1225|Green||2013-10-24|2013-10-29|NaT||||40.2||1|1|1|1|M|Black||10|No|Mother|28215|2|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|White||29|28211|Bachelors Degree|Single|Business: Marketing|28262|3|0|Recruitment Event|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|502934732|502936151|31|0|1|503537424|1|0|1|500722866|10|2|-2||2|1||-2|500000294|-2|0|10|||7458|9|||1||4575902950186762737|0
M1582|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|295|Green|PERL 2014-2016|2014-12-11|2014-12-11|2015-10-02|Volunteer: Time constraint|Volunteer: Time constraint||9.7||3|3|1|1|F|Multi-race (Black & Hispanic)||10||Mother|28025||One Parent: Female|Unknown||||Yes||School|General Site|Cabarrus County, PERL 2014-2016|Match Support|F|White||19|28031|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500002335|504106223|504108257|38|0|2|504043405|1|0|2|500803670|10|1|500000296|2128173571|4|1|500014681, 500016374|-1|500014681|-1|0|4|||0|4|||1|500014681|5208542183136337346|0
M1583|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|244|Yellow||2016-02-09|2016-02-26|2016-10-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8||3|3|1|1|F|Multi-race (Black & Hispanic)||10||Mother|28025||One Parent: Female|Unknown||||Yes||School|General Site|Cabarrus County, PERL 2014-2016|Match Support|F|White||18|28025|Some High School|Single|Student: College||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504106223|504108257|38|0|2|504579772|1|0|2|500878416|10|1|500000296|2128173571|4|2|500014681, 500016374|-1|500016374|-1|0|4|||7464|9|||1||5208542183136337346|0
M1584|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|119|Green|Cabarrus County|2016-10-31|2016-11-08|NaT||||3.9||3|3|2|2|F|Multi-race (Black & Hispanic)||10||Mother|28025||One Parent: Female|Unknown||||Yes||School|General Site|Cabarrus County, PERL 2014-2016|Match Support|F|Hispanic||17|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504106223|504108257|38|0|2|504579805|3|0|2|500921828|10|1|500000296|2128173571|2|1|500014681, 500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|5208542183136337346|0
M1585|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|97|Green|Amachi|2015-09-11|2015-09-23|2015-12-29|Child: Lost interest|Child: Lost interest||3.2||1|1|1|1|F|Black||10|Yes|GrandMother|28217|4|Grandparents|Less than $10,000|||Y|Yes||School|General Community|Amachi|Match Support|F|White||32|28277|Masters Degree|Divorced|Tech: Computer/Programmer|28277|0|3|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017732|504195472|504197572|31|0|2|504222207|1|0|2|500839514|10|2|-2||4|1|500000294|-2|500000294|-2|0|4|||7464|9|||1|500000294|7857548027029642592|0
M1586|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|198|Green||2016-03-11|2016-03-15|2016-09-29|Child/Family: Moved|Child/Family: Moved||6.5||1|1|2|2|M|Black||10|No|Mother|28025|3|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|Cabarrus County|Match Support|F|White||17|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504652703|504655124|31|0|1|504629049|1|0|2|500884395|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||643003066716863548|0
M1587|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|627|Green||2013-10-08|2013-11-01|2015-07-21|Volunteer: Moved|Volunteer: Moved||20.6||3|3|1|1|F|Hispanic||10|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503204707|503206461|3|0|2|503497191|1|0|2|500717215|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1588|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|509|Green||2015-10-09|2015-10-15|NaT||||16.7||3|3|1|1|F|Hispanic||10|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|503204707|503206461|3|0|2|504302580|1|0|2|500846390|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1589|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|62|Green||2016-11-22|2017-01-04|NaT||||2||1|1|2|2|F|Black||10|Yes|Mother|28229|5|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|Black||17|28269|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504951143|504953694|31|0|2|504301152|31|0|2|500930449|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1590|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|221|Yellow|PERL 2014-2016|2015-01-23|2015-01-30|2015-09-08|Child/Family: Moved|Child/Family: Moved||7.3||1|1|1|1|M|Hispanic||10|No|Mother|28025|2|Two Parent|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|White||31|29732||Single|Retail: Mgt||0|0|Recruitment Event|Workplace Partner|Big|General Site|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500012459|504167666|504169774|3|0|1|504035902|1|0|2|500809874|10|1|500000295|2128212924|4|2|500014681|-1|500014681|-1|0|4|||7446|3|||1|500014681|3232906304025417619|0
M1591|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1115|Green||2013-07-11|2013-07-30|2016-08-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||36.6||1|1|1|1|M|White||10|No|Mother|28210|2|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|Asian||29|28134|Masters Degree|Single|Finance: Accountant|28202|1|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500021785|503471046|503472912|1|0|1|503489178|4|0|1|500703315|10|2|-2||4|1||-2|500000294|-2|0|10|||7496|10|||1||2272605169937511837|8528216325355383116
M1592|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1475|Green||2013-02-14|2013-02-21|NaT||||48.5||1|1|1|1|M|Black||10|No|Mother|28217|4|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|M|White||28|28209|Masters Degree|Single|Finance: Accountant||0|6|Relative|Relative|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502778215|502610737|31|0|1|503291713|1|0|1|500682140|10|2|-2||2|1||-2||-2|0|3|||17161|11|||1||5386346637278076349|0
M1593|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|489|Green||2015-10-16|2015-11-04|NaT||||16.1||1|1|1|1|F|Asian||10|No|Father|28212|3|Two Parent|$30,000 to $34,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504478043|504480317|4|0|2|504306207|1|0|2|500848721|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1594|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|605|Green||2014-10-07|2014-10-17|2016-06-13|Volunteer: Moved|Volunteer: Moved||19.9||1|1|1|1|M|Hispanic||10|No|Mother|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|M|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504050669|504052693|3|0|1|503925833|1|0|1|500781520|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1595|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|603|Red||2013-06-13|2013-06-26|2015-02-19|Volunteer: Time constraint|Volunteer: Time constraint||19.8||2|2|1|1|F|Black||10||Mother|28216|4|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||55|28209|Some College|Divorced|Business: Clerical|28273|20|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503259551|503261359|31|0|2|503371077|1|0|2|500700569|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1||8568001799025358453|7044657180546140448
M1596|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|593|Green||2015-06-26|2015-07-23|NaT||||19.5||2|2|1|1|F|Black||10||Mother|28216|4|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Business: Human Resources|28202|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503259551|503261359|31|0|2|504219483|1|0|2|500831431|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1||8568001799025358453|7044657180546140448
M1597|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|402|Green|Cabarrus County|2016-01-22|2016-01-30|NaT||||13.2||1|1|1|1|F|Multi-race (Hispanic & White)||10|No|Mother|28025|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||25|28269||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504532725|504535058|35|0|2|503951023|1|0|2|500874940|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||7496|10|||1|500016374|643003066716863548|2141487034287122220
M1598|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|167|Green||2016-09-01|2016-09-21|NaT||||5.5||1|1|1|1|M|White||10|No|Mother|28226|3|One Parent: Female|$35,000 to $39,999|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||30|28226|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|1|Other|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504379951|504382189|1|0|1|504736110|1|0|1|500905929|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316|-2|0|10|||7671|13|||1||5893332617597240023|1706608681384859512
M1599|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|335|Green||2015-10-16|2015-11-04|2016-10-04|Child: Changed school/site|Child: Changed school/site||11||1|1|2|2|M|Black||10|No|Mother|28215|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|M|White||18|28211||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504443661|504445917|31|0|1|504311367|1|0|1|500848820|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1600|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|572|Green||2015-07-23|2015-08-13|NaT||||18.8||1|1|1|1|F|Black||10|No|Mother|28216|2|One Parent: Female|$30,000 to $34,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||34|28031||Single|Self-Employed, Entrepreneur||9|8|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504186133|504188242|31|0|2|504122609|1|0|2|500834256|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1||2056258660718146620|8136849793711030748
M1601|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|49|Green||2016-11-29|2017-01-17|NaT||||1.6||2|2|1|1|F|Black||10|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504449710|504451966|31|0|2|504708194|1|0|2|500931395|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1602|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|420|Green||2015-10-05|2015-10-06|2016-11-29|Volunteer: Time constraint|Volunteer: Time constraint||13.8||2|2|1|1|F|Black||10|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504449710|504451966|31|0|2|504311336|1|0|2|500844172|10|1|500000296|2128173564|4|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1603|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|303|Green||2015-03-28|2015-03-29|2016-01-26|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||10||1|1|2|2|M|Black||10|No|Mother|28213|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||Therapist/Counselor|General Community||Enrollment|M|Black||35|28273|Some College|Married|Business: Marketing|28203|1|1|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500018987|504005000|504007015|31|0|1|504241664|31|0|1|500820944|5|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|5|||46|2|||1||4013586283864837776|1044653023923149817
M1604|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|228|Green|PERL 2014-2016|2015-11-09|2016-01-14|2016-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.5||1|1|1|1|F|Black||10|No|Mother|28056|4|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||RTBM|F|White||30|28209|Bachelors Degree|Single|Finance: Banking|28211|3|2|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500017777|504407275|504409521|31|0|2|504393547|1|0|2|500857377|7|2|-2||4|1||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|500014681|7679812394383646966|0
M1605|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|346|Yellow||2015-04-07|2015-04-20|2016-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.4||2|2|1|1|F|Black||10|No|Mother|28206|2|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Enrollment|F|White||29|28205|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|3|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503834826|503836805|31|0|2|504139505|1|0|2|500822171|5|2|-2||4|2||-2||-2|0|10|||17159|12|||1||421482027904269589|0
M1606|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|148|Green||2016-09-20|2016-10-10|NaT||||4.9||1|1|2|2|M|Black||10|Yes|Mother|28214|4|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||30|28209|Bachelors Degree|Married|Real Estate: Realtor|28217|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504759201|504761658|31|0|1|504322037|1|0|1|500908756|10|2|-2||2|1|500014681|-2||-2|0|10|||46|2|||1||6095563712459522926|7105699653014118193
M1607|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|968|Green||2013-11-26|2013-11-26|2016-07-21|Volunteer: Moved|Volunteer: Moved||31.8||2|2|1|1|M|Black||10|No|Mother|28031|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||22|28035|Some College|Single|Student: College||0|0|Self|Self|Big|General Site|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500015820|503720474|503252163|31|0|1|503638772|31|0|1|500735056|10|1|500000295|2128173570|4|1||-1|500000294|-1|0|4|||7464|9|||1||8034889377453131101|0
M1608|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|155|Green||2016-09-26|2016-10-03|NaT||||5.1||2|2|1|1|M|Black||10|No|Mother|28031|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||20|28035||Single|Student: College||0|0|Self|Self|Big|General Site|VOL - PreMatch|Match Support|0|1|0|1|277|60|598|500000170|500015820|503720474|503252163|31|0|1|504685604|31|0|1|500910306|10|1|500000295|2128173570|2|1||-1|500007920|-1|0|4|||7464|9|||1||8034889377453131101|0
M1609|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|494|Green||2015-10-23|2015-10-30|NaT||||16.2||1|1|1|1|F|Hispanic||10|No|Mother|28212|3|Two Parent|$30,000 to $34,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504478270|504480544|3|0|2|504307889|1|0|2|500851485|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1610|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|374|Red||2014-10-29|2014-11-21|2015-11-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.3||1|1|1|1|M|White||10|No|Mother|28270|1|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Enrollment|M|White||28|28270|Bachelors Degree|Living w/ Significant Other|Law: Police Officer|28211|0|9|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|503873009|503875005|1|0|1|503953864|1|0|1|500789610|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1||5790136262762328632|3810421262203348915
M1611|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1778|Green||2012-03-21|2012-04-24|NaT||||58.4||1|1|1|1|F|Black||10|No|GrandMother|28208||Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||31|28209|Masters Degree|Single|Medical: Healthcare Worker|28079|0|4|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|502946633|502948059|31|0|2|502893902|1|0|2|500605537|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1||0|3402014428779854546
M1612|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|988|Green||2014-06-12|2014-06-23|NaT||||32.5||1|1|1|1|F|Black||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|Black||35|28104|Some College|Single|Medical: Healthcare Worker|28105|2|7|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500020910|503582752|502908938|31|0|2|503771996|31|0|2|500766377|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||5741767063897867874|4374719395834495975
M1613|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1141|Green|Cabarrus County|2014-01-17|2014-01-21|NaT||||37.5||1|1|1|1|F|White||10|No|Father|28081|4|One Parent: Male|Unknown|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|White||50|28226|Bachelors Degree||Human Services: Non-Profit|28208|0|6|Self|Self|Big|General Community|Cabarrus County|Enrollment|1|0|0|1|277|60|598|500000170|500013781|503634722|503636659|1|0|2|503597445|1|0|2|500743535|10|2|-2||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|4619448746907815971|1786514887916898235
M1614|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|813|Green||2014-12-01|2014-12-15|NaT||||26.7||1|1|1|1|M|Black||10|No|Mother|28206|1|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||28|28203|Masters Degree|Single|Business|28277|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503671417|503673378|31|0|1|504022116|1|0|1|500799802|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1||7987165241089060600|1558599596122179496
M1615|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|661|Yellow||2013-04-19|2013-04-22|2015-02-12|Child/Family: Moved|Child/Family: Moved||21.7||1|1|1|1|F|Black||10|No|Mother|28216|2|One Parent: Female|$10,000 to $14,999|||Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||28|28205|Bachelors Degree|Single|Business|28255|0|3|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500015820|503230851|503232639|31|0|2|503317475|1|0|2|500693795|5|2|-2||4|2||-2|500000294|-2|6854|8|||7464|9|||1||7960300212314874874|3866301893856809726
M1616|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|498|Green||2015-10-16|2015-10-26|NaT||||16.4||1|1|1|1|F|Hispanic||10|No|Father|28212|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504468544|503779890|3|0|2|504297069|1|0|2|500848783|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1617|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|379|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-09|2016-02-22|NaT||||12.5||1|1|1|1|F|Multi-race (Black & White)||10|Yes|Foster Parent|28216|4|One Parent: Female|$40,000 to $44,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||45|28208|Bachelors Degree|Single|Education: Teacher|28208|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504498650|504500981|36|0|2|504131389|31|0|2|500878445|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1|500007920, 500011315, 500011316|2456895876914964961|0
M1618|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|700|Green||2015-03-30|2015-03-30|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||23||1|1|1|1|F|Black||10|Yes|Mother|28273|2|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Black||29|28269||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|504165894|504167953|31|0|2|504138163|31|0|2|500821104|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1||5711791743715234276|5161383151676749743
M1619|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|120|Green||2016-10-17|2016-10-26|2017-02-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||3.9||1|1|1|1|M|Black||10|No|Mother|28208|3|One Parent: Female|$35,000 to $39,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business|28203|2|9|BBBS National Site|Web Link|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020910|503401421|503403278|31|0|1|504818783|1|0|1|500916185|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-1|34|2|||46|2|||1||7508998544817094399|5096023753338979088
M1620|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|496|Green||2015-10-16|2015-10-28|NaT||||16.3||1|1|1|1|M|Black||10|No|Mother|28212|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site|VOL - HSBigs|Match Support|M|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504442284|504444540|31|0|1|504302566|1|0|1|500848813|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1621|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|349|Yellow|Cabarrus County|2016-03-09|2016-03-23|NaT||||11.5||1|1|1|1|M|Black||10|No|Mother|28027|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||35|28083|High School Graduate|Married|Medical||8|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504563369|504565703|31|0|1|504600175|1|0|1|500883737|10|2|500016307||2|2|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|500016374|3325175628848876741|6200244613298520712
M1622|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|664|Green||2015-05-08|2015-05-13|NaT||||21.8||1|1|1|1|F|White||10|No|Mother|28214|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|F|White||28|28206|Bachelors Degree|Single|Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504231269|504233379|1|0|2|503927707|1|0|2|500826291|10|2|-2||2|1||-2||-2|0|3|||46|2|||1||7089569121628268952|0
M1623|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|105|Green||2016-11-18|2016-11-22|NaT||||3.4||1|1|1|1|M|Black||10|No|Mother|28211|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Site||Match Support|F|White||16|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504412845|504415101|31|0|1|504727827|1|0|2|500929294|10|1|500000296|2128173564|2|1||-1||-1|0|10|||0|4|||1||2762897743412756173|0
M1624|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|517|Red|VOL - Mentoring Hispanic Youth|2015-03-19|2015-03-31|2016-08-29|Child: Family structure changed|Child: Family structure changed||17||1|1|1|1|M|Hispanic||10|No|Mother|28214|2|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|VOL - Mentoring Hispanic Youth|Match Support|M|Hispanic||40|28277|Bachelors Degree|Married|Insurance|28277|8|0|Current/Previous Big|Other Big|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|0|1|1|0|277|60|598|500000170|500017777|504059287|504061304|3|0|1|504210666|3|0|1|500819684|10|2|-2||4|3|500011312|-2|500011312|-2|0|5|||17159|12|||1|500011312|5604470640552265812|0
M1625|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|300|Green|PERL 2014-2016|2015-11-30|2015-12-04|2016-09-29|Child/Family: Moved|Child/Family: Moved||9.9||1|1|6|6|F|Black||10|No|Mother|28083|3|One Parent: Female|Unknown||||Yes||Relative|General Site|Cabarrus County, PERL 2014-2016|Match Support|F|Black||38|28269|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500012459|504530709|504533041|31|0|2|500189256|31|0|2|500863845|10|1|500000295|2128232374|4|1|500014681, 500016374|-1|500007920, 500011315, 500011316, 500016374|-1|0|3|||7464|9|1360|3|1|500014681|2043334928777030191|0
M1626|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1197|Red||2013-06-10|2013-06-18|2016-09-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||39.3||1|1|1|1|M|Black||10|Yes|GrandMother|28208|0|One Parent: Female|$10,000 to $14,999|||Y|Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Enrollment|M|White||29|28269|Masters Degree|Living w/ Significant Other|Business: Mgt, Admin|28203|0|7|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|503144476|503146148|31|0|1|503453981|1|0|1|500700084|5|2|-2||4|3|500000294|-2|500000294|-2|7294|13|||7464|9|||1||7679812394383646966|1786514887916898235
M1627|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|27|Green||2017-01-11|2017-02-08|NaT||||0.9||1|1|1|1|M|Black||10|No|Mother|28211|2|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|M|Black||38|28227|Bachelors Degree|Single|Business: Marketing|28202|4|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504417080|504419332|31|0|1|504872445|31|0|1|500939553|10|2|-2||2|1|500007920, 500011315, 500011316, 500014681|-2|500007920, 500011315, 500011316|-2|0|5|||46|2|||1||5367149751093883357|2763237020791144915
M1628|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|677|Green|PERL 2014-2016|2015-04-11|2015-04-30|NaT||||22.2||1|1|2|2|M|Multi-race (Black & Hispanic)||10|Yes|GrandMother|28208|1|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community|Amachi, PERL 2014-2016|Match Support|M|Asian||33|28204|Bachelors Degree|Married|Business: Engineer|28007|3|9|Man Up Campaign|Media|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|503433219|503227914|38|0|1|503890372|4|0|1|500822826|10|2|-2||2|1|500000294, 500014681|-2|500000294, 500014681|-2|0|10|||17101|1|||1|500014681|8998367770661215127|7044657180546140448
M1629|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|902|Green||2014-09-12|2014-09-17|NaT||||29.6||1|1|1|1|M|Multi-race (Black & Hispanic)||10|No|Mother|28212|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||27|28211|Bachelors Degree|Single|Finance|29715|1|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503836529|503838508|38|0|1|503876514|1|0|1|500775633|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1||2762897743412756173|7044657180546140448
M1630|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|482|Green|PERL 2014-2016|2015-10-29|2015-11-11|NaT||||15.8||1|1|1|1|F|Black||10|No|Mother|28216|3|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Hispanic||26|28031|Bachelors Degree|Single|Tech: Research/Design|28117|0|8|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504390954|504393193|31|0|2|504231700|3|0|2|500853984|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1|500014681|2979941694006626856|3650724132819756420
M1631|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|573|Green||2014-04-03|2014-04-25|2015-11-19|Volunteer: Time constraint|Volunteer: Time constraint||18.8||1|1|1|1|M|Black||10|Yes|Mother|28216|1|One Parent: Female|$45,000 to $49,999|||Y|Yes||Self|General Community||Match Support|M|White||33|28031|Bachelors Degree|Single|Tech: Engineer|28081|6|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503662361|503664337|31|0|1|503740772|1|0|1|500758213|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||3664007741235143067|7044657180546140448
M1632|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|908|Green||2014-08-20|2014-09-11|NaT||||29.8||1|1|1|1|M|Black||10|No|Mother|28217|1|One Parent: Female|$25,000 to $29,999|||Y|Yes||Relative|General Community||Match Support|M|White||47|28278|Bachelors Degree|Married|Business: Mgt, Admin|29732|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503835875|503837854|31|0|1|503926804|1|0|1|500772936|10|2|-2||2|1||-2||-2|0|3|||17159|12|||1||0|7560981454869879219
M1633|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|105|Green||2016-11-17|2016-11-22|NaT||||3.4||1|1|1|1|F|Some Other Race||10|No|Mother|28212|3|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504933441|504935992|41|0|2|504712714|1|0|2|500929159|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1634|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|927|Green||2014-01-02|2014-01-17|2016-08-01|Volunteer: Moved|Volunteer: Moved||30.5||2|2|1|1|M|Black||10|No|Mother|28078|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||22|28031|Some College|Single|Student: College||0|0|Kappa Alpha Psi|Fraternity/Sorority|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500015820|503471483|503473349|31|0|1|503641249|31|0|1|500740954|10|1|500000295|2128173570|4|1||-1||-1|0|4|||8693|14|||1||8034889377453131101|0
M1635|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|155|Green||2016-09-21|2016-10-03|NaT||||5.1||2|2|1|1|M|Black||10|No|Mother|28078|5|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||21|28035||Single|Student: College||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|503471483|503473349|31|0|1|504631163|31|0|1|500909237|10|1|500000295|2128173570|2|1||-1||-1|0|4|||7464|9|||1||8034889377453131101|0
M1636|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|153|Green||2016-03-29|2016-04-29|2016-09-29|Volunteer: Time constraint|Volunteer: Time constraint||5||2|2|2|2|M|Black||10|No|Mother|28202|3|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||RTBM|M|White||31|28203|Bachelors Degree|Single|Construction|28208|1|1|Igniting Breakfast|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500021785|503804106|503712061|31|0|1|502255664|1|0|1|500886730|7|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|10|||17266|8|||1||6368218764956286027|5056473444237941296
M1637|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|380|Green||2014-09-24|2014-09-29|2015-10-14|Volunteer: Moved|Volunteer: Moved||12.5||2|2|1|1|M|Black||10|No|Mother|28202|3|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||RTBM|M|White||25|28209|Bachelors Degree|Single|Tech: Computer/Programmer|28202|0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503804106|503712061|31|0|1|503988181|1|0|1|500777910|7|2|-2||4|1||-2||-2|0|10|||7464|9|||1||6368218764956286027|5056473444237941296
M1638|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|12|Green||2017-02-03|2017-02-23|NaT||||0.4||1|1|2|2|M|Black||10|No|Mother|28214|2|One Parent: Female|$25,000 to $29,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|504486089|504488364|31|0|1|502643791|3|0|1|500944356|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1||0|6570326659017849719
M1639|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|288|Yellow||2014-10-22|2014-11-10|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||9.5||1|1|1|1|F|Black||10|No|Mother|28203|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||RTBM|F|White||34|28203|Masters Degree|Single|Business||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|504051221|504053245|31|0|2|503972520|1|0|2|500786442|7|2|-2||4|2||-2||-2|0|4|||17159|12|||1||8568001799025358453|7044657180546140448
M1640|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1421|Green||2013-04-15|2013-04-16|NaT||||46.7||1|1|1|1|F|Black||10|No|Mother|28215|2|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community||Match Support|F|White||33|28210|Bachelors Degree|Single|Tech: Support, Writing|28217|0|6|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503224812|503226552|31|0|2|503385277|1|0|2|500692915|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1||2417657944362725638|0
M1641|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|495|Green||2015-10-29|2015-10-29|NaT||||16.3||1|1|1|1|F|Black||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|White||18|28173|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504495854|504498139|31|0|2|504303214|1|0|2|500853665|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1642|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-31|2016-10-31|NaT||||4.2||1|1|1|1|M|Black||10|Yes|Mother|28208|3|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|M|Black||46|28277|Some College|Married|Business|28277|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504401349|504403590|31|0|1|504856770|31|0|1|500921965|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||0|4309014537710246316
M1643|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|503|Green||2015-10-16|2015-10-21|NaT||||16.5||1|1|1|1|F|Black||10|No|Mother|28211|3|One Parent: Female|Less than $10,000||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504476395|504478669|31|0|2|504302545|1|0|2|500848846|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1644|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|182|Green||2016-08-18|2016-09-06|NaT||||6||1|1|1|1|M|Black||10|Yes|Mother|28212|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|White||24|28202|Bachelors Degree|Single|Finance: Banking|28202|0|2|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504260162|504262304|31|0|1|504639207|1|0|1|500903992|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||0|4802885652788112046
M1645|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|236|Green||2016-06-29|2016-07-14|NaT||||7.8||2|2|1|1|F|Black||10|No|Mother|28208|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||39|28278|Masters Degree|Married|Business: Human Resources|28217|1|7|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|503589761|503591638|31|0|2|504552375|1|0|2|500898409|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1||976372749760822282|7044657180546140448
M1646|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|718|Yellow||2013-10-11|2013-10-28|2015-10-16|Volunteer: Health|Volunteer: Health||23.6||2|2|1|1|F|Black||10|No|Mother|28208|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Child/Day Care Worker|28214|10|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|503589761|503591638|31|0|2|503582412|1|0|2|500718535|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1||976372749760822282|7044657180546140448
M1647|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|554|Green||2014-03-27|2014-03-27|2015-10-02|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.2||3|3|1|1|M|Black||10|No|Mother|28025||Other/Unknown|Unknown||||No||Therapist/Counselor|General Site|Cabarrus County|Match Support|M|White||20|28215|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500002335|503669403|503671364|31|0|1|503553049|1|0|1|500757038|10|1|500000296|2128173571|4|1|500016374|-1||-1|0|5|||0|4|||1||4085045877112350207|0
M1648|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|412|Green|Cabarrus County|2016-01-14|2016-01-20|NaT||||13.5||3|3|1|1|M|Black||10|No|Mother|28025||Other/Unknown|Unknown||||No||Therapist/Counselor|General Site|Cabarrus County|Match Support|M|White||17|28036|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|503669403|503671364|31|0|1|504549032|1|0|1|500872045|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|5|||0|4|||1|500016374|4085045877112350207|0
M1649|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|105|Green||2016-11-22|2016-11-22|NaT||||3.4||1|1|2|2|M|Black||10|No|Mother|28212|4|Two Parent|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28209|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504896413|504898933|31|0|1|504296421|1|0|1|500930418|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|5708657394834009072
M1650|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|171|Yellow||2015-02-04|2015-02-27|2015-08-17|Child/Family: Moved|Child/Family: Moved||5.6||1|1|1|1|F|Black||10|No|Mother|28206|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Business: Sales||0|10|Recruitment Event|BBBS Board/Staff|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500015820|504168597|504170705|31|0|2|504161094|1|0|2|500812001|10|2|-2||4|2||-2||-2|0|4|||7462|13|||1||4863631750424600365|7044657180546140448
M1651|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|876|Green||2013-03-11|2013-03-27|2015-08-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.8||1|1|1|1|M|Black||10|No|Mother|28205|1|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||34|28203|Masters Degree|Single|Real Estate: Realtor||5|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503001538|503003032|31|0|1|503380945|1|0|1|500686972|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1||7987165241089060600|7044657180546140448
M1652|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|388|Green|Cabarrus County|2016-02-01|2016-02-13|NaT||||12.7||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28025|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||28|28027|Masters Degree|Single|Govt|28273|3|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504468562|504470835|36|0|1|504556956|31|0|1|500876668|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|500016374|5173041326630627506|7044657180546140448
M1653|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1392|Green||2013-04-04|2013-05-15|NaT||||45.7||1|1|1|1|M|Multi-race (Black & White)||10||Mother|28226|1|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Multi-race (Asian & White)||35|28209|Bachelors Degree|Single|Business: Mgt, Admin||1|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503321228|503323062|36|0|1|503412979|37|0|1|500691563|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||5893332617597240023|7044657180546140448
M1654|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|189|Green||2016-08-10|2016-08-30|NaT||||6.2||1|1|2|2|M|Black||10|No|Mother|28277|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||51|28277|Bachelors Degree|Married|Finance|28277|0|0|Igniting Breakfast|Special Event|Big|General Community|mentor2.0, mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500017732|504660516|504662943|31|0|1|503922166|1|0|1|500902981|10|2|-2||2|1||-2|500014505, 500014506|-2|0|10|||17266|8|||1||7617270550840231462|7044657180546140448
M1655|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|366|Green||2015-03-24|2015-04-13|2016-04-13|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12||1|1|1|1|F|Black||10|No|Mother|28206|2|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||23|28262||Single|Student: College||0|0|Current/Previous Big|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500018851|504211769|504213882|31|0|2|504100154|1|0|2|500820237|10|2|-2||4|1||-2||-2|0|5|||17159|12|||1||7960300212314874874|0
M1656|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|91|Green||2016-11-18|2016-12-06|NaT||||3||2|2|2|2|F|Multi-race (Black & Hispanic)||10|No|Father|28212|3|Two Parent|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504495820|504498105|38|0|2|504297164|1|0|2|500929291|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1657|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|341|Green||2015-10-29|2015-10-29|2016-10-04|Child: Changed school/site|Child: Changed school/site||11.2||2|2|2|2|F|Multi-race (Black & Hispanic)||10|No|Father|28212|3|Two Parent|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504495820|504498105|38|0|2|504297164|1|0|2|500853876|10|1|500000296|2128173564|4|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1658|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1099|Green||2014-02-03|2014-03-04|NaT||||36.1||1|1|1|1|M|Black||10|No|Mother|28226|1|One Parent: Female|$20,000 to $24,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Some Other Race||38|28277|Masters Degree|Married|Finance: Banking|28228|7|0|Big For A Day|Special Event|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503650774|503652734|31|0|1|503526078|41|0|1|500746685|10|2|-2||2|1||-2||-2|34|2|||16422|8|||1||4726905079488957916|894086896518290414
M1659|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|572|Green|PERL 2014-2016|2014-10-15|2014-10-22|2016-05-16|Volunteer: Time constraint|Volunteer: Time constraint||18.8||1|1|1|1|F|Black||10|No|Mother|28213|2|One Parent: Female|$30,000 to $34,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||32|28270|Associate Degree|Married|Arts, Entertainment, Sports|28203|3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500018851|503995241|503997256|31|0|2|503924249|1|0|2|500783860|10|2|-2||4|1|500014681|-2|500014681|-2|34|2|||17159|12|||1|500014681|0|7045146654760389673
M1660|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|334|Green||2015-10-28|2015-11-04|2016-10-03|Child: Changed school/site|Child: Changed school/site||11||1|1|2|2|F|Black||10|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500022905|504449730|504451986|31|0|2|504307828|1|0|2|500853505|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1661|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|722|Green||2015-03-08|2015-03-16|NaT||||23.7||1|1|1|1|M|Black||10|No|Mother|28211|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||31|28209|Bachelors Degree|Married|Medical|70112|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503314773|503314167|31|0|1|504176084|1|0|1|500817494|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||2762897743412756173|4253272603994307857
M1662|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|588|Green||2015-07-23|2015-07-28|NaT||||19.3||1|1|1|1|M|Black||10||GrandMother|28213|2|Grandparents|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||28|28204||Single|Finance: Accountant|28277|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503022461|501332937|31|0|1|504323998|1|0|1|500834322|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||6065435025527210335|0
M1663|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|118|Green|Cabarrus County|2016-10-31|2016-11-09|NaT||||3.9||1|1|1|1|F|Black||10|No|Mother|28025|4|Two Parent|Unknown|Yes: Active|No||Yes||School|General Site|Cabarrus County|Match Support|F|Asian||17|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504918193|504920713|31|0|2|504884057|4|0|2|500921836|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|5208542183136337346|0
M1664|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|155|Green||2016-09-16|2016-10-03|NaT||||5.1||1|1|1|1|M|Black||10|No|Mother|28273|3|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||33|28273|Bachelors Degree|Married|Tech: Computer/Programmer|28262|9|4|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504391010|504393249|31|0|1|504614273|1|0|1|500908114|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||1834158761762606452|703802826159951755
M1665|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|811|Green||2014-12-08|2014-12-17|NaT||||26.6||2|2|1|1|F|Black||10|Yes|GrandMother|28031|4|Grandparents|Unknown|||Y|Yes||School|General Site||Match Support|F|White||46|28078|Some College|Married|Govt|28031|7|3|Current/Previous Big|Other Big|Big|General Site||Match Support|1|0|0|1|277|60|598|500000170|500015820|503873448|503875444|31|0|2|503889163|1|0|2|500802076|10|1|500000295|2128173570|2|1||-1||-1|0|4|||17159|12|||1||8034889377453131101|0
M1666|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|227|Green||2015-10-29|2015-10-29|2016-06-12|Volunteer: Moved|Volunteer: Moved||7.5||1|1|2|2|M|Asian||10|No|Mother|28262|3|Two Parent|$10,000 to $14,999|||Y|Yes||School|General Site|VOL - HSBigs|RTBM|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504495871|504498156|4|0|1|503901733|1|0|2|500853684|7|1|500000296|2128173564|4|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1667|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1006|Green||2014-06-02|2014-06-05|NaT||||33.1||1|1|1|1|M|Black||10|No|Mother|28262|4|One Parent: Female|$50,000 to $59,999|Yes: Active|No||No||Self|General Community||Match Support|M|Black||46|28078||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503468785|503470651|31|0|1|503856524|31|0|1|500765157|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1||4356567821563751981|786532283575222488
M1668|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|644|Green||2013-10-08|2013-11-01|2015-08-07|Volunteer: Moved|Volunteer: Moved||21.2||2|2|1|1|F|Hispanic||10|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503391580|503393421|3|0|2|503509851|1|0|2|500717213|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1669|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|503|Green||2015-10-09|2015-10-21|NaT||||16.5||2|2|1|1|F|Hispanic||10|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|503391580|503393421|3|0|2|504303256|1|0|2|500846326|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1670|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|329|Yellow||2014-04-04|2014-04-10|2015-03-05|Volunteer: Time constraint|Volunteer: Time constraint||10.8||2|2|1|1|M|Black||10|Yes|Mother|28216|1|One Parent: Female|Less than $10,000||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||43|28269|Bachelors Degree|Married|Business: Marketing|28262|2|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|503565647|503567522|31|0|1|503577080|1|0|1|500758415|10|2|-2||4|2|500000294|-2||-2|34|2|||7464|9|1360|3|1||2979941694006626856|1786514887916898235
M1671|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|708|Green||2015-03-19|2015-03-30|NaT||||23.3||2|2|2|2|M|Black||10|Yes|Mother|28216|1|One Parent: Female|Less than $10,000||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||42|28205|Bachelors Degree|Married|Arts, Entertainment, Sports|28205|14|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020910|503565647|503567522|31|0|1|503865770|1|0|1|500819520|10|2|-2||2|1|500000294|-2|500000294|-2|34|2|||17159|12|||1||2979941694006626856|1786514887916898235
M1672|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|509|Green||2015-10-14|2015-10-15|NaT||||16.7||1|1|1|1|M|Black||10|No|Mother|28211|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|VOL - HSBigs|Match Support|M|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504297445|504299659|31|0|1|504306075|1|0|1|500847670|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|3260639349613832803
M1673|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green||2015-10-29|2015-11-11|NaT||||15.8||1|1|1|1|F|Hispanic||10|No|Father|28212|3|Two Parent|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504495828|504498113|3|0|2|504296415|1|0|2|500854002|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1674|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|659|Green||2013-09-30|2013-09-30|2015-07-21|Volunteer: Moved|Volunteer: Moved||21.7||2|2|1|1|F|Hispanic||10|No|Mother|28212|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28207||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503637758|503639718|3|0|2|503498727|1|0|2|500714444|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1675|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|503|Green||2015-10-09|2015-10-21|NaT||||16.5||2|2|1|1|F|Hispanic||10|No|Mother|28212|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|503637758|503639718|3|0|2|504297025|1|0|2|500846328|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1676|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|537|Green||2014-11-05|2014-11-05|2016-04-25|Child/Family: Moved|Child/Family: Moved||17.6||1|1|1|1|F|Black||10|No|Mother|28212|4|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||19|28205|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020909|504101686|504103720|31|0|2|503907516|31|0|2|500792058|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1677|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|519|Yellow||2014-03-10|2014-03-24|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||17.1||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28081|K|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||51|28027|Some College|Married|Business: Marketing|28027|1|5|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503461190|503463056|36|0|1|503672434|1|0|1|500753717|10|2|||4|2||-2||-2|0|10|||7464|9|||1||0|4022520458090739403
M1678|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|736|Yellow||2015-01-29|2015-02-23|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.2||1|1|1|1|M|Multi-race (Black & White)||10|Yes|Mother|28204|1|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||26|28216|Bachelors Degree|Single|Tech: Engineer|28078|0|4|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503812210|503814187|36|0|1|504084695|1|0|1|500810906|10|2|-2||4|2||-2||-2|0|10|||46|2|||1||7960300212314874874|7044657180546140448
M1679|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|659|Green||2013-09-30|2013-09-30|2015-07-21|Volunteer: Moved|Volunteer: Moved||21.7||2|2|1|1|M|Hispanic||10|No|Mother|28212|K|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||20|29715|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503418294|503420158|3|0|1|503507180|1|0|1|500714485|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1680|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|473|Green||2015-10-16|2015-11-20|NaT||||15.5||2|2|1|1|M|Hispanic||10|No|Mother|28212|K|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||18|28078|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|503418294|503420158|3|0|1|504311115|1|0|1|500848822|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1681|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green|VOL - HSBigs|2016-11-16|2016-11-28|NaT||||3.3||1|1|1|1|F|Hispanic||10|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504932802|504935353|3|0|2|504718131|1|0|2|500928280|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1|500014068|2762897743412756173|0
M1682|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|455|Green||2015-11-30|2015-12-08|NaT||||14.9||1|1|1|1|M|Black||10|No|Mother|28208|2|One Parent: Female|Less than $10,000|||Y|Yes|TV|Media|General Community||Match Support|M|White||27|28203|Bachelors Degree|Single|Insurance|21202|2|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504046908|504048929|31|0|1|504349113|1|0|1|500863535|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|56|1|||17159|12|||1||976372749760822282|7044657180546140448
M1683|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|747|Red|PERL 2014-2016|2014-08-26|2014-09-18|2016-10-04|Child: Family structure changed|Child: Family structure changed||24.5||1|1|2|2|M|Multi-race (Black & White)||10|Yes|Mother|28025|1|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016, VOL - Incarcerated Parents|Match Support|M|Asian||27|28075|Bachelors Degree|Single|Finance: Banking|28202|3|0|Local Print|Media|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500020753|503681425|503683390|36|0|1|503786945|4|0|1|500773494|10|2|-2||4|3|500007918, 500014681, 500016374|-2|500014681, 500016374|-2|34|2|||7439|1|||1|500014681|5173041326630627506|2141487034287122220
M1684|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|18|Green||2017-02-06|2017-02-17|NaT||||0.6||1|1|1|1|M|Black||10|No|Mother|28269|3|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|M|White||24|28208|Bachelors Degree|Single|Tech: Management|28203|0|5|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504811851|504814332|31|0|1|504883582|1|0|1|500944658|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|3|||7464|9|||1||6077912216232501082|7044657180546140448
M1685|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|96|Green||2014-10-04|2014-10-17|2015-01-21|Child/Family: Moved|Child/Family: Moved||3.2||2|2|2|2|M|Hispanic||10|No|Mother|28212||One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||19|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503241971|503243768|3|0|1|503901671|1|0|1|500780608|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1686|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|105|Green||2016-10-21|2016-11-22|NaT||||3.4||2|2|1|1|F|Black||10|No|Mother|28215|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||27|28204|Masters Degree||Business: Human Resources|28202|0|3|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|503602769|503604646|31|0|2|504787610|31|0|2|500918350|10|2|-2||2|1|500007920, 500011315, 500011316, 500014681|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||1158671944891395407|1786514887916898235
M1687|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|413|Green||2014-10-23|2014-11-10|2015-12-28|Volunteer: Moved|Volunteer: Moved||13.6||2|2|1|1|F|Black||10|No|Mother|28215|4|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||25|28213|Bachelors Degree|Single|Finance: Banking|28216|0|10|Billboard|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020990|503602769|503604646|31|0|2|503919845|31|0|2|500787263|10|2|-2||4|1|500007920, 500011315, 500011316, 500014681|-2||-2|0|10|||125|1|||1||1158671944891395407|1786514887916898235
M1688|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|244|Green|Cabarrus County|2016-07-05|2016-07-06|NaT||||8||1|1|1|1|F|Hispanic||10|No|Mother|28027|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|White||47|28081||Married|Finance: Banking||18|5|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504724296|504726733|3|0|2|504746325|1|0|2|500898734|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|500016374|3232906304025417619|0
M1689|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|200|Red|PERL 2014-2016|2015-04-30|2015-05-14|2015-11-30|Volunteer: Time constraint|Volunteer: Time constraint||6.6||1|1|1|1|M|Black||10|No|Mother|28212|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|PERL 2014-2016|Enrollment|M|White||28|28105|Bachelors Degree|Married|Tech: Computer/Programmer|28272|2|7|Local TV|Media|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500008321|504122686|504124721|31|0|1|504171365|1|0|1|500825432|5|2|-2||4|3|500014681|-2|500014681|-2|0|4|||7438|1|||1|500014681|5386346637278076349|0
M1690|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|182|Green||2015-11-11|2015-11-16|2016-05-16|Child/Family: Moved|Child/Family: Moved||6||1|1|1|1|M|Black||10|No|Mother|28031|2|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||23|28036|Some College|Single|Student: College||0|0|Self|Self|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504462301|504464559|31|0|1|503680396|31|0|1|500858694|10|1|500000295|2128173570|4|1||-1||-1|0|4|||7464|9|||1||8034889377453131101|0
M1691|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|496|Green||2015-10-16|2015-10-28|NaT||||16.3||1|1|1|1|F|Hispanic||10|No|Mother|28212|3|Two Parent|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504478000|504480274|3|0|2|504306150|1|0|2|500848855|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1692|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|496|Yellow|Cabarrus County|2015-10-19|2015-10-28|NaT||||16.3||1|1|2|2|M|Black||9|No|Mother|28027|4|One Parent: Female|$75,000 to $99,999||||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|Black||34|28269|Some College|Married|Business|28025|5|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County, mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500022817|503911799|503913806|31|0|1|503956879|31|0|1|500849358|10|2|500016307||2|2|500016374|-2|500014506, 500016374|-2|34|2|||7671|13|||1|500016374|0|0
M1693|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|372|Yellow||2016-02-23|2016-02-29|NaT||||12.2||2|2|1|1|M|White||9|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||22|28215|Some College|Single|Finance|28215|0|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|503661137|503646117|1|0|1|504531427|1|0|1|500881061|10|2|-2||2|2||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||2762897743412756173|0
M1694|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|580|Green||2013-10-15|2013-11-01|2015-06-04|Volunteer: Moved|Volunteer: Moved||19.1||2|2|1|1|M|White||9|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||20|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503661137|503646117|1|0|1|503507155|1|0|1|500719614|10|1|500000296|2128173564|4|1||-2||-1|0|4|||0|4|||1||2762897743412756173|0
M1695|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|82|Green||2016-12-05|2016-12-15|NaT||||2.7||2|2|1|1|M|White||9|No|Mother|28212|4|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||42|28205|Bachelors Degree||Business|28202|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|503644157|503646117|1|0|1|504605644|1|0|1|500932984|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||2762897743412756173|0
M1696|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|604|Green||2013-10-07|2013-10-08|2015-06-04|Volunteer: Moved|Volunteer: Moved||19.8||2|2|1|1|M|White||9|No|Mother|28212|4|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503644157|503646117|1|0|1|503500364|1|0|1|500716294|10|1|500000296|2128173564|4|1||-2||-1|0|4|||0|4|||1||2762897743412756173|0
M1697|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|496|Green||2015-10-16|2015-10-28|NaT||||16.3||1|1|1|1|M|Black||9|Yes|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|M|White||18|28207|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504441601|504443857|31|0|1|504306403|1|0|1|500848814|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1698|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|508|Green||2015-10-15|2015-10-16|NaT||||16.7||1|1|1|1|M|Black||9|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|M|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504449694|504451950|31|0|1|504311015|1|0|1|500848540|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1699|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1477|Green||2013-02-18|2013-02-19|NaT||||48.5||1|1|1|1|F|Black||9|No|Father|28213|K|One Parent: Male|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Black||56|28269|Bachelors Degree|Single|Business: Mgt, Admin|28262|25|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503226693|503228481|31|0|2|503035671|31|0|2|500682567|10|2|500014421||2|1||-2||-2|0|4|||7671|13|||1||7679812394383646966|5605796235524810842
M1700|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|927|Green||2014-07-17|2014-08-23|NaT||||30.5||1|1|3|3|F|Black||9|No|Mother|28213|1|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|Black||29|28262|Bachelors Degree|Single|Student: College||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503883171|503885167|31|0|2|502138981|31|0|2|500769877|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1||6713311931049891381|7044657180546140448
M1701|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|222|Green|PERL 2014-2016|2016-07-21|2016-07-28|NaT||||7.3||1|1|1|1|F|Black||9|No|Mother|28217||One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Some Other Race||25|28208|Bachelors Degree|Single|Business: Sales|28278|0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504601619|504604030|31|0|2|504611053|41|0|2|500900279|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||46|2|||1|500014681|0|727731964632783453
M1702|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|609|Green||2014-10-04|2014-10-07|2016-06-07|Volunteer: Moved|Volunteer: Moved||20||2|2|1|1|F|Black||9|No|Mother|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Some Other Race||18|28173|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504042033|504044051|31|0|2|503916425|41|0|2|500780588|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1703|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|2|2|F|Black||9|No|Mother|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504042033|504044051|31|0|2|504303791|1|0|2|500929329|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1704|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|957|Green||2014-07-09|2014-07-24|NaT||||31.4||1|1|1|1|M|Black||9|Yes|Mother|28262|1|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|M|White||31|28117|Bachelors Degree|Single|Finance: Accountant|28677|0|5|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503587467|503587387|31|0|1|503886373|1|0|1|500768974|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1||836952159905822963|5766455966581408090
M1705|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|119|Green|Cabarrus County|2016-10-31|2016-11-08|NaT||||3.9||1|1|2|2|F|Black||9|Yes|Mother|28083|4|Two Parent|$30,000 to $34,999|Yes: Active|No||No||School|General Site|Cabarrus County|Match Support|F|White||17|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504918404|504920924|31|0|2|504629049|1|0|2|500921816|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|0|0
M1706|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|198|Green||2016-02-09|2016-02-26|2016-09-11|Volunteer: Time constraint|Volunteer: Time constraint||6.5||2|2|1|1|F|White||9|No|Father|28027|3|One Parent: Male|Less than $10,000||||Yes||School|General Site|Cabarrus County|Match Support|F|White||17|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504600029|504602440|1|0|2|504579912|1|0|2|500878405|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||6810228174639243761|0
M1707|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|119|Green|Cabarrus County|2016-11-01|2016-11-08|NaT||||3.9||2|2|1|1|F|White||9|No|Father|28027|3|One Parent: Male|Less than $10,000||||Yes||School|General Site|Cabarrus County|Match Support|F|White||17|28083|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504600029|504602440|1|0|2|504884009|1|0|2|500922401|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|6810228174639243761|0
M1708|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|797|Green||2014-05-21|2014-05-31|2016-08-05|Volunteer: Moved|Volunteer: Moved||26.2||1|1|1|1|M|Black||9|No|Mother|28208|1|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||31|28277|Bachelors Degree|Single|Finance: Economist|28277|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503778456|503780433|31|0|1|503787440|1|0|1|500763996|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1||4356567821563751981|4365185292611375158
M1709|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|372|Green|Cabarrus County|2016-02-09|2016-02-29|NaT||||12.2||1|1|1|1|F|White||9|No|Mother|28027|3|Two Parent|$30,000 to $34,999||||Yes||School|General Site|Cabarrus County|Match Support|F|Hispanic||18|28025|Some High School|Single|Student: College||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504619564|504621975|1|0|2|504579789|3|0|2|500878410|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|6810228174639243761|0
M1710|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|332|Green||2015-10-09|2015-10-26|2016-09-22|Volunteer: Moved|Volunteer: Moved||10.9||1|1|1|1|M|Black||9|No|Mother|28211|4|One Parent: Female|$25,000 to $29,999|Yes: Active|No|Y|Yes||Self|General Community||RTBM|M|Multi-race (Black & White)||26|28211|Some College|Single|Finance|28210|0|5|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504345299|504347523|31|0|1|504397824|36|0|1|500846354|7|2|-2||4|1||-2||-2|0|10|||46|2|||1||421482027904269589|1981915209225039472
M1711|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|166|Green||2016-09-01|2016-09-22|NaT||||5.5||1|1|1|1|M|Black||9|No|Mother|28273|3|One Parent: Female|$35,000 to $39,999||||Yes||School|General Community||Match Support|M|White||41|28226|Bachelors Degree|Married|Business: Sales|28273|4|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504403567|504405809|31|0|1|504689704|1|0|1|500905927|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||5386346637278076349|4318803846885526429
M1712|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|601|Green||2013-10-18|2013-10-25|2015-06-18|Volunteer: Moved|Volunteer: Moved||19.7||1|1|1|1|F|Black||9|No|Mother|28208|1|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|F|White||26|28209|Bachelors Degree|Single|Retail: Sales|28209|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503589735|503591612|31|0|2|503488419|1|0|2|500720851|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1||3935539763241716148|3727920003273999020
M1713|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|90|Green||2016-11-14|2016-12-07|NaT||||3||1|1|2|2|M|White||9|No|Mother|28031|4|One Parent: Female|$15,000 to $19,999||||No||School|General Site||Match Support|M|Black||20|28035|||Student: College||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504909745|504912265|1|0|1|504634278|31|0|1|500927446|10|1|500000295|2128173570|2|1||-1||-1|0|4|||7464|9|||1||8034889377453131101|0
M1714|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1391|Green||2013-05-01|2013-05-16|NaT||||45.7||2|2|1|1|F|Black||9|No|Mother|28215|K|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||54|28211|Bachelors Degree|Separated|Retired||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|503062537|501090456|31|0|2|503455629|1|0|2|500695323|10|2|-2||2|1||-2||-2|0|10|||7462|13|||1||5741767063897867874|4753237757252407321
M1715|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|61|Green||2017-01-04|2017-01-05|NaT||||2||1|1|1|1|M|Black||9|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||16|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504976151|504978702|31|0|1|504722603|1|0|2|500938132|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1716|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|987|Green||2014-06-18|2014-06-24|NaT||||32.4||1|1|1|1|M|Multi-race (Black & Hispanic)||9|No|Mother|28215|1|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Hispanic||37|28202|Bachelors Degree|Single|Consultant|27607|1|0|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503774068|503776034|38|0|1|503866555|3|0|1|500767047|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1||4575902950186762737|0
M1717|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|169|Green|PERL 2014-2016|2016-09-07|2016-09-19|NaT||||5.6||1|1|1|1|F|Black||9|No|Mother|28216|3|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|Black||42|28105|Bachelors Degree|Married|Business|28277|0|2|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504604960|504607371|31|0|2|504374080|31|0|2|500906296|10|2|-2||2|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||46|2|||1|500014681|1653226628427425023|2876415545463317777
M1718|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|936|Green||2014-08-06|2014-08-14|NaT||||30.8||1|1|1|1|F|Black||9|No|GrandMother|28216|1|Grandparents|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||48|28269|Some College|Married|Finance: Banking|28262|0|0|Current/Previous Big|Relative|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|503866363|503838583|31|0|2|503946948|1|0|2|500771529|10|2|-2||2|1||-2|500000294|-2|0|10|||17160|11|||1||7679812394383646966|9060571453147419923
M1719|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|800|Green|PERL 2014-2016|2014-10-27|2014-11-04|2017-01-12|Volunteer: Time constraint|Volunteer: Time constraint||26.3||1|1|1|1|F|Black||9|No|Aunt|28208|1|Other Relative|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||54|28078|Associate Degree|Single|Medical|28025|10|7|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500020910|503862843|502431630|31|0|2|503926694|1|0|2|500788150|5|2|-2||4|1|500014681|-2|500000294, 500014681|-2|0|10|||7464|9|||1|500014681|3038247238543299436|0
M1720|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green||2015-10-16|2015-11-11|NaT||||15.8||1|1|1|1|F|Hispanic||9|No|Mother|28212|3|Two Parent|Less than $10,000||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504468558|504470831|3|0|2|504296388|1|0|2|500848725|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1721|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|678|Red||2013-07-26|2013-08-15|2015-06-24|Volunteer: Moved|Volunteer: Moved||22.3||1|1|1|1|M|Multi-race (Black & Asian)||9||Mother|28226|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|M|White||29|28208|Bachelors Degree|Single|Unknown|28202|0|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503476611|503478477|39|0|1|503495634|1|0|1|500704993|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1||4726905079488957916|776646640278297723
M1722|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|100|Yellow||2015-02-11|2015-02-23|2015-06-03|Volunteer: Time constraint|Volunteer: Time constraint||3.3||1|1|1|1|M|Black||9|No|Mother|28213|1|One Parent: Female|$20,000 to $24,999||||Yes|Radio|Media|General Community||RTBM|M|Black||28|28269|Bachelors Degree|Single|Business: Sales|28213|1|6|Kappa Alpha Psi|Fraternity/Sorority|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503856979|503858973|31|0|1|504170817|31|0|1|500813164|7|2|-2||4|2||-2||-2|55|1|||8693|14|||1||6627885846854295604|7795805164050330858
M1723|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|503|Green||2015-10-11|2015-10-21|NaT||||16.5||1|1|1|1|F|Black||9|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Black||17|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504449703|504178342|31|0|2|504302426|31|0|2|500846533|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1724|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|822|Green|PERL 2014-2016|2014-11-25|2014-11-28|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||27||1|1|1|1|F|Black||9|No|Mother|28208|2|One Parent: Female|$25,000 to $29,999||||No||School|General Community|PERL 2014-2016|Enrollment|F|Black||22|28208|Bachelors Degree|Single|Medical: Nurse|28278|0|7|Self|Self|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500018851|504106075|503933644|31|0|2|503995246|31|0|2|500799241|5|2|-2||4|1|500014681|-2|500014681|-2|0|4|||7464|9|||1|500014681|7089569121628268952|8626610080771140821
M1725|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|560|Green||2015-07-23|2015-08-25|NaT||||18.4||1|1|1|1|M|Black||9|No|Mother|28262|2|One Parent: Female|$30,000 to $34,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||40|28202|Bachelors Degree|Single|Self-Employed, Entrepreneur||7|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503967629|503969639|31|0|1|504276405|1|0|1|500834265|10|2|-2||2|1||-2||-2|34|2|||46|2|||1||6627885846854295604|6619197389800008587
M1726|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|364|Green||2016-03-03|2016-03-08|NaT||||12||1|1|1|1|F|Black||9|No|Mother|28208|3|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||24|28202|Bachelors Degree|Single|Business|28202|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|504445747|504448003|31|0|2|504321583|1|0|2|500882893|10|2|-2||3|1||-2||-2|34|2|||46|2|||1||6077912216232501082|3866301893856809726
M1727|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-12|2016-10-31|NaT||||4.2||1|1|1|1|M|Black||9|No|Mother|28212||One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|M|White||33|28202|PHD|Single|Real Estate: Realtor|28269|3|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504399529|504394964|31|0|1|504803637|1|0|1|500915028|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||6627885846854295604|3727915399477748546
M1728|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|127|Green||2016-10-12|2016-10-31|NaT||||4.2||1|1|1|1|M|Black||9|No|Mother|28212|3|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||32|28209||Single|Finance|28202|2|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504392725|504394964|31|0|1|504697126|1|0|1|500914996|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||6627885846854295604|3727915399477748546
M1729|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|214|Green||2016-01-22|2016-02-10|2016-09-11|Child: Changed school/site|Child: Changed school/site||7||1|1|4|4|F|White||9|No|Father|28027|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site|Cabarrus County|Match Support|F|Multi-race (Black & White)||23|28273|Some College|Single|Student: College|28227|0|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500012459|504579529|504581863|1|0|2|503853917|36|0|2|500874836|10|1|500000295|2128232374|4|1|500016374|-1|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7464|9|||1||3232906304025417619|0
M1730|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|174|Green||2015-10-28|2015-10-28|2016-04-19|Child/Family: Moved|Child/Family: Moved||5.7||1|1|2|2|M|Black||9|No|Mother|28205|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504443675|504445931|31|0|1|504310910|1|0|1|500853489|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1731|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|118|Green|Cabarrus County|2016-10-17|2016-11-09|NaT||||3.9||2|2|1|1|M|Black||9|No|Mother|28025|3|Other Relative|Less than $10,000|||Y|Yes||School|General Site|Cabarrus County|Match Support|M|White||17|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504605295|504607706|31|0|1|504875740|1|0|1|500916297|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|3324851395989241799|0
M1732|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|213|Green||2016-02-18|2016-02-29|2016-09-29|Volunteer: Time constraint|Volunteer: Time constraint||7||2|2|1|1|M|Black||9|No|Mother|28025|3|Other Relative|Less than $10,000|||Y|Yes||School|General Site|Cabarrus County|Match Support|M|White||17|28025|Some High School||Student: High School||0|0||High School Partner|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504605295|504607706|31|0|1|504629024|1|0|1|500880190|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||0|4|||1||3324851395989241799|0
M1733|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|257|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-06-16|2016-06-23|NaT||||8.4||1|1|1|1|F|Black||9|No|Mother|28215|3|One Parent: Female|$75,000 to $99,999||||Yes||School|General Community||Match Support|F|White||35|28215|Associate Degree|Divorced|Business|28215|0|8|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504507824|504510119|31|0|2|504575855|1|0|2|500896954|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1|500007920, 500011315, 500011316|6627885846854295604|4318803846885526429
M1734|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|345|Green||2014-10-29|2014-10-29|2015-10-09|Child: Changed school/site|Child: Changed school/site||11.3||1|1|2|2|F|White||9|No|Mother|28211|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504081854|504083883|1|0|2|503905493|1|0|2|500789754|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1735|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|473|Green||2015-11-16|2015-11-20|NaT||||15.5||1|1|1|1|M|Black||9|No|Mother|28212|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504478286|504480560|31|0|1|504297003|1|0|2|500860351|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1736|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|252|Green||2016-06-10|2016-06-28|NaT||||8.3||1|1|1|1|M|Black||9|No|Mother|28203|3|Two Parent|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||26|28202|Masters Degree|Single|Finance: Economist||0|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504601244|504603655|31|0|1|504577016|1|0|1|500896409|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|5|||7464|9|||1||8568001799025358453|904091744937704216
M1737|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|574|Green||2014-11-11|2014-11-17|2016-06-13|Volunteer: Moved|Volunteer: Moved||18.9||2|2|1|1|F|Hispanic||9|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||19|28278|Some High School|Single|Student: College||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504112150|504114144|3|0|2|503907569|1|0|2|500794590|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1738|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|2|2|F|Hispanic||9|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||18|28227|Some High School|Single|Student: College||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504112150|504114144|3|0|2|504296357|1|0|2|500928279|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1739|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|1257|Green||2013-09-25|2013-09-27|NaT||||41.3||1|1|2|2|M|Black||9|No|Mother|28078|3|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||47|28650|Bachelors Degree|Single|Personal Trainer/Coach||0|0|Michael Baisden|Media|Big|General Site|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500015820|503471487|503473349|31|0|1|502163847|31|0|1|500712990|10|1|500000295|2128173570|2|1||-1|500000294|-1|0|4|||11272|1|||1||8034889377453131101|0
M1740|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green||2016-11-30|2016-12-05|NaT||||3||1|1|1|1|F|Hispanic||9|No|Mother|28212|3|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||17|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504943196|504945747|3|0|2|504712668|1|0|2|500931723|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1741|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|91|Green||2016-11-16|2016-12-06|NaT||||3||1|1|1|1|M|Black||9|Yes|Mother|28226|3|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Site||Match Support|F|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504931624|504934175|31|0|1|504731990|1|0|2|500928283|10|1|500000296|2128173564|2|1||-1||-1|0|3|||0|4|||1||2762897743412756173|6604057783730669766
M1742|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|174|Green||2016-08-18|2016-09-14|NaT||||5.7||2|2|2|2|F|Black||9|No|Mother|28216|4|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||34|28078|Masters Degree|Single|Medical: Doctor, Provider|28001|0|2|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500013781|503454717|504995618|31|0|2|503323641|1|0|2|500903980|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||2979941694006626856|0
M1743|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|608|Green||2014-10-04|2014-10-08|2016-06-07|Volunteer: Moved|Volunteer: Moved||20||1|1|1|1|M|Hispanic||9|No|Mother|28212|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|M|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049330|504043821|3|0|1|503905491|1|0|1|500780594|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1744|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|139|Green||2016-09-21|2016-10-19|NaT||||4.6||1|1|1|1|M|Black||9|No|Mother|28262|2|One Parent: Female|$50,000 to $59,999||||No||School|General Community||Match Support|M|Black||35|28269|Masters Degree|Married|Business: Sales|29708|2|3|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504203765|504205876|31|0|1|504766376|31|0|1|500909175|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||4748|14|||1||7102230088759381237|3402014428779854546
M1745|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|106|Green||2016-11-04|2016-11-21|NaT||||3.5||1|1|2|2|F|Black||9|No|Mother|28208|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Hispanic||36|28210|Bachelors Degree|Married|Finance: Accountant|28203|4|0|BBBS National Site|Web Link|Big|General Site|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500015820|504886739|504889259|31|0|2|504000676|3|0|2|500924987|10|1|500000295|2128207319|2|1||-1|500014681|-1|0|4|||46|2|||1||3935539763241716148|0
M1746|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|270|Green||2016-05-02|2016-06-10|NaT||||8.9||1|1|2|2|F|Black||9|No|Mother|28031|3|Two Parent|$15,000 to $19,999|||Y|No||School|General Community||Match Support|F|White||48|28031|Bachelors Degree|Separated|Business: Marketing|28601|16|0|BBBS National Site|Web Link|Big|General Community|Amachi, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504577424|504579758|31|0|2|503698988|1|0|2|500891352|10|2|-2||2|1||-2|500000294, 500007920, 500011315, 500011316|-2|0|4|||46|2|||1||0|7137064858903755892
M1747|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|134|Green||2016-10-17|2016-10-24|NaT||||4.4||1|1|1|1|F|White||9|No|Aunt|28031|3|Other Relative|$50,000 to $59,999||||Yes||School|General Site||Match Support|F|White||55|28031|||Business||0|11|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504842848|504845350|1|0|2|504676684|1|0|2|500916575|10|1|500000295|2128173570|2|1||-1||-1|0|4|||18809|8|||1||8034889377453131101|5498785567357422131
M1748|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|105|Green|Cabarrus County|2016-11-04|2016-11-22|NaT||||3.4||1|1|6|6|F|Black||9|No|Mother|28083|4|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|Cabarrus County|Match Support|F|Black||38|28269|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500012459|504922812|504925332|31|0|2|500189256|31|0|2|500924982|10|1|500000295|2128232374|2|1|500016374|-1|500007920, 500011315, 500011316, 500016374|-1|0|4|||7464|9|1360|3|1|500016374|2043334928777030191|0
M1749|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|83|Green|Cabarrus County|2016-12-08|2016-12-14|NaT||||2.7||1|1|3|3|M|Black||9|No|Mother|28083|4|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|Cabarrus County|Match Support|M|Black||37|28273||Married|Business||0|0|ACN|Workplace Partner|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504936878|504925332|31|0|1|503216970|31|0|1|500934060|10|1|500000295|2128232374|2|1|500016374|-1|500016374|-1|0|4|||13581|3|||1|500016374|2043334928777030191|0
M1750|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|413|Green||2015-11-24|2016-01-19|NaT||||13.6||2|2|2|2|F|Black||9|No|Mother|28031|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||70|28031||Divorced|Consultant||0|0|Self|Self|Big|General Site|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500015820|504220461|504222575|31|0|2|503633204|1|0|2|500863240|10|1|500000295|2128173570|2|1||-1|500000294|-1|0|4|||7464|9|||1||8034889377453131101|0
M1751|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|265|Yellow||2015-02-27|2015-02-27|2015-11-19|Child/Family: Moved|Child/Family: Moved||8.7||2|2|1|1|F|Black||9|No|Mother|28031|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||63|28036|Masters Degree|Married|Business: Sales||3|6|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504220461|504222575|31|0|2|504029691|1|0|2|500816078|10|1|500000295|2128173570|4|2||-1||-1|0|4|||17159|12|||1||8034889377453131101|0
M1752|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|51|Green|Cabarrus County|2016-12-19|2017-01-15|NaT||||1.7||3|3|1|1|F|White||9|No|Mother|28027|2|Two Parent|Unknown||||Yes||School|General Community|Cabarrus County|Match Support|F|White||46|28027|High School Graduate|Married|Business: Sales|28078|2|2|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|503225825|503227613|1|0|2|504862689|1|0|2|500936501|10|2|500016307||2|1|500016374|-2|500016374|-2|0|4|||17159|12|||1|500016374|6810228174639243761|0
M1753|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|720|Red||2014-11-12|2014-11-19|2016-11-08|Volunteer: Time constraint|Volunteer: Time constraint||23.7||3|3|1|1|F|White||9|No|Mother|28027|2|Two Parent|Unknown||||Yes||School|General Community|Cabarrus County|Match Support|F|White||29|28138|Bachelors Degree|Single|Customer Service|28269|2|5|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500020753|503225825|503227613|1|0|2|503551624|1|0|2|500794940|10|2|-2||4|3|500016374|-2|500016374|-2|0|4|||7464|9|||1||6810228174639243761|0
M1754|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|362|Green||2016-03-04|2016-03-10|NaT||||11.9||1|1|1|1|M|Black||9|No|Mother|28213|3|One Parent: Female|$35,000 to $39,999||||Yes||School|General Community||Match Support|M|White||41|28078|Bachelors Degree|Married|Self-Employed, Entrepreneur|28031|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504262369|504264514|31|0|1|504538390|1|0|1|500883013|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||540227296891876425|2806833304218536184
M1755|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green|VOL - HSBigs|2016-11-17|2016-11-28|NaT||||3.3||1|1|1|1|M|Hispanic||9|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022908|504934152|504936703|3|0|1|504707562|1|0|1|500929179|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1|500014068|2762897743412756173|0
M1756|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|118|Green|Cabarrus County|2016-11-01|2016-11-09|NaT||||3.9||1|1|1|1|F|Multi-race (Black & White)||9|No|GrandMother|28025|4|Grandparents|Unknown|Yes: Active|No||Yes||School|General Site|Cabarrus County|Match Support|F|White||18|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504919512|504922026|36|0|2|504892783|1|0|2|500922382|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|1550830965009450729|0
M1757|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1150|Red|Cabarrus County|2013-09-06|2013-09-25|2016-11-18|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||37.8||1|1|3|3|F|Black||9|No|GrandMother|28083|K|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|F|Black||45|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500022817|503585543|503587420|31|0|2|500189320|31|0|2|500709465|10|2|500016307||4|3|500016374|-2|500016374|-2|34|2|||7464|9|||1|500016374|6810228174639243761|0
M1758|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|91|Green||2016-11-18|2016-12-06|NaT||||3||1|1|1|1|M|Hispanic||9|No|Father|28212|3|One Parent: Male|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|Hispanic||16|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504930090|504932641|3|0|1|504741770|3|0|2|500929343|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1759|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green|VOL - HSBigs|2016-11-16|2016-12-05|NaT||||3||1|1|1|1|F|Multi-race (Black & White)||9|No|Mother|28211|3|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504932947|504935498|36|0|2|504722595|1|0|2|500928481|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1|500014068|2762897743412756173|2127318745563037380
M1760|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|16|Green|Cabarrus County|2017-02-14|2017-02-19|NaT||||0.5||1|1|2|2|M|Black||9|No|Mother|28081|3|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||24|28081|Some High School|Single|Service: Hotel||4|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504902017|504904537|31|0|1|501028238|31|0|1|500946229|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||17159|12|||1|500016374|3142304990634129454|2544020271035850193
M1761|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-16|2016-11-30|NaT||||3.2||1|1|1|1|F|Hispanic||9|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||17|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504932921|504935472|3|0|2|504725071|1|0|2|500928475|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1762|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green||2016-11-18|2016-12-05|NaT||||3||1|1|1|1|F|Black||9|No|Mother|28212|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||16|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504932725|504935276|31|0|2|504719725|1|0|2|500929364|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1763|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|119|Green||2016-11-04|2016-11-08|NaT||||3.9||1|1|1|1|M|Black||9|No|Mother|28208|3|Two Parent|$10,000 to $14,999||||Yes||School|General Site||Match Support|M|White||28|28105|Bachelors Degree|Single|Business||3|9|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504886700|504889220|31|0|1|504777354|1|0|1|500924913|10|1|500000295|2128207319|2|1||-1||-1|0|4|||18809|8|||1||3935539763241716148|7451594515531114270
M1764|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|8|Green||2017-02-06|2017-02-27|NaT||||0.3||1|1|1|1|F|Black||9|No|Mother|28269|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Multi-race (Black & White)||21|28213|Some College|Single|Business: Sales|28211|0|9|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504673056|504675483|31|0|2|504845407|36|0|2|500944794|10|2|-2||2|1|500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||64486389764866818|7044657180546140448
M1765|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|795|Green|Amachi|2014-08-13|2014-08-29|2016-11-01|Volunteer: Time constraint|Volunteer: Time constraint||26.1||1|1|1|1|F|Black||9|Yes|Mother|28208|2|One Parent: Female|Less than $10,000||||Yes||Therapist/Counselor|General Community|Amachi|Enrollment|F|White||26|28209|Masters Degree|Single|Education: Teacher|28212|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|503953662|503955662|31|0|2|503952799|1|0|2|500772194|5|2|-2||4|1|500000294|-2||-2|0|5|||7496|10|||1|500000294|0|7044657180546140448
M1766|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green|VOL - HSBigs|2016-11-16|2016-11-28|NaT||||3.3||1|1|1|1|F|Black||9|No|Mother|28212|3|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Site||Match Support|F|White||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504934155|504936706|31|0|2|504708831|1|0|2|500928443|10|1|500000296|2128173564|2|1||-1||-1|0|3|||0|4|||1|500014068|2762897743412756173|0
M1767|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|405|Green||2016-01-14|2016-01-27|NaT||||13.3||1|1|1|1|M|White||9|No|Mother|28105|2|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504574836|504577170|1|0|1|504303283|1|0|2|500872025|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1768|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|519|Yellow|Amachi|2014-04-28|2014-04-30|2015-10-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.1||1|1|1|1|F|Black||9|Yes|Mother|28269|K|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||26|28212|Some College||Medical: Nurse||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500012459|503798419|503800396|31|0|2|502994003|31|0|2|500761356|10|2|-2||4|2|500000294|-2|500000294|-2|34|2|||7462|13|||1|500000294|967246839551912690|7795805164050330858
M1769|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|49|Green||2017-01-10|2017-01-17|NaT||||1.6||1|1|1|1|F|Black||9|No|GrandMother|28212|3|Grandparents|Unknown||||Yes||School|General Site||Match Support|F|White||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504970016|504972567|31|0|2|504708027|1|0|2|500939291|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1770|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|589|Green||2014-12-01|2014-12-10|2016-07-21|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||19.4||1|1|1|1|M|Black||9|No|Mother|28206|2|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||59|28078|Masters Degree|Married|Firefighter|28202|28|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500016270|503996764|503998741|31|0|1|503889103|31|0|1|500799922|10|1|500000295|2128173561|4|1||-1||-1|0|4|||7496|10|||1||7960300212314874874|0
M1771|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-16|2016-11-30|NaT||||3.2||1|1|1|1|F|Hispanic||9|No|Mother|28212|3|Two Parent|$20,000 to $24,999||||Yes||Relative|General Site||Match Support|F|White||16|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504933050|504935601|3|0|2|504707396|1|0|2|500928434|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M1772|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|372|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-17|2016-02-29|NaT||||12.2||1|1|1|1|M|Black||9|No|Mother|28214|2|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|White||23|28202|Bachelors Degree|Single|Consultant|28202|0|5|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500021785|504153377|504155427|31|0|1|504487777|1|0|1|500879869|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|500007920, 500011315, 500011316|7089569121628268952|1335047838269305508
M1773|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green|VOL - HSBigs|2016-11-16|2016-11-28|NaT||||3.3||1|1|1|1|M|Hispanic||9|No|Mother|28212|3|Two Parent|Unknown||||Yes||Relative|General Site||Match Support|M|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504932900|504935451|3|0|1|504718207|1|0|1|500928450|10|1|500000296|2128173564|2|1||-1||-1|0|3|||0|4|||1|500014068|2762897743412756173|0
M1774|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green||2016-11-18|2016-12-05|NaT||||3||1|1|1|1|M|Black||9|No|Mother|28222|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504933011|504935562|31|0|1|504718087|1|0|2|500929319|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1775|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|91|Green||2016-11-16|2016-12-06|NaT||||3||1|1|1|1|F|Black||9|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504931636|504934187|31|0|2|504722516|1|0|2|500928454|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1776|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|615|Green||2015-07-01|2015-07-01|NaT||||20.2||1|1|1|1|M|Black||9|No|Mother|28269|1|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|M|Black||28|28205|Bachelors Degree|Single|Finance|28202|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504219209|504221323|31|0|1|504301519|31|0|1|500831883|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||0|0
M1777|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|622|Green||2014-09-29|2014-09-30|2016-06-13|Volunteer: Moved|Volunteer: Moved||20.4||1|1|1|1|F|Black||9|No|Mother|28217|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504030927|504032945|31|0|2|503905447|1|0|2|500778749|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1778|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|363|Green|Cabarrus County|2016-03-03|2016-03-09|NaT||||11.9||1|1|1|1|M|White||9|No|Mother|28083|2|One Parent: Female|Less than $10,000||||Yes||School|General Site|Cabarrus County|Match Support|M|White||83|28081||Widowed|Retired||0|0|Self|Self|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500012459|504530646|504532978|1|0|1|504637067|1|0|1|500882896|10|1|500000295|2128232374|2|1|500016374|-1|500007920, 500011315, 500011316, 500016374|-1|0|4|||7464|9|||1|500016374|2043334928777030191|0
M1779|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|683|Green||2015-04-24|2015-04-24|NaT||||22.4||1|1|1|1|F|Multi-race (Black & Hispanic)||9|No|Mother|28269|1|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||30|28206|Masters Degree|Single|Human Services: Psychologist|28211|2|2|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504220029|504222143|38|0|2|504198281|1|0|2|500824763|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||5367149751093883357|7044657180546140448
M1780|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|61|Green||2016-12-06|2017-01-05|NaT||||2||1|1|1|1|F|White||9|No|Step-Father|28211|3|Two Parent|$20,000 to $24,999|||Y|Yes||School|General Site||Match Support|F|White||17|28211|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504965759|504968310|1|0|2|504718233|1|0|2|500933616|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1781|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|374|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-22|2016-02-27|NaT||||12.3||1|1|1|1|F|Black||9|Yes|Mother|28208|2|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|F|Black||35|28216|Masters Degree|Married|Medical||0|3|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504404998|504403590|31|0|2|504481744|31|0|2|500880569|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|500007920, 500011315, 500011316|0|4309014537710246316
M1782|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1350|Green||2013-06-25|2013-06-26|NaT||||44.4||1|1|1|1|F|Black||9||Mother|28216|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||29|28269|Bachelors Degree|Single|Medical: Nurse||1|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503286862|503261359|31|0|2|503386901|1|0|2|500701858|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||8568001799025358453|7044657180546140448
M1783|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|366|Yellow||2015-07-16|2015-07-28|2016-07-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12||1|1|2|2|M|Black||9|No|Mother|28215|1|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Enrollment|M|Hispanic||31|28209|High School Graduate|Single|Finance|28262|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|504039337|504041355|31|0|1|504011759|3|0|1|500833679|5|2|-2||4|2||-2||-2|0|4|||46|2|||1||5741767063897867874|7044657180546140448
M1784|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|287|Red||2014-05-19|2014-05-22|2015-03-05|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||9.4||2|2|2|2|M|Black||9|Yes|Mother|28204|3|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|White||42|28205|Bachelors Degree|Married|Arts, Entertainment, Sports|28205|14|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017777|503663973|503665933|31|0|1|503865770|1|0|1|500763734|10|2|-2||4|3||-2|500000294|-2|0|10|||17159|12|||1||6407809237813394802|0
M1785|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|135|Green||2016-04-13|2016-05-17|2016-09-29|Volunteer: Time constraint|Volunteer: Time constraint||4.4||2|2|1|1|M|Black||9|Yes|Mother|28204|3|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|White||25|28209|Bachelors Degree|Single|Finance|28277|0|9|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500021785|503663973|503665933|31|0|1|504568754|1|0|1|500888979|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||6407809237813394802|0
M1786|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green|VOL - HSBigs|2016-11-17|2016-12-05|NaT||||3||1|1|1|1|F|Black||9|No|Mother|28205|3|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|Black||17|28273|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504943089|504945640|31|0|2|504725175|31|0|2|500929169|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1|500014068|2762897743412756173|2084013234086765119
M1787|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|362|Green||2016-02-23|2016-03-10|NaT||||11.9||1|1|1|1|F|Black||9|No|Mother|28217|2|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||42|28210|Bachelors Degree|Single|Business|28262|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504425557|504427813|31|0|2|504124868|1|0|2|500880862|10|2|-2||3|1||-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1||8981704271528751143|482329911636883098
M1788|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|554|Green|PERL 2014-2016, Cabarrus County|2015-08-14|2015-08-31|NaT||||18.2||1|1|1|1|F|Black||9|No|Mother|28075|1|Two Parent|$10,000 to $14,999||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||26|28027|Bachelors Degree|Single|Medical|28025|0|8|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504298787|504301001|31|0|2|504325174|31|0|2|500836212|10|2|500016307||2|1|500014681, 500016374|-2|500016374|-2|0|4|||46|2|||1|500014681, 500016374|3380316005507597709|7044657180546140448
M1789|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|923|Green||2014-08-20|2014-08-27|NaT||||30.3||1|1|1|1|M|Black||9|No|Mother|28208|K|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||35|28217|Some College|Married|Law: Police Officer|28229|0|8|Man Up Campaign|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503739912|503702247|31|0|1|503929189|31|0|1|500772941|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1||2611337051335117774|7044657180546140448
M1790|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|90|Green||2016-12-06|2016-12-07|NaT||||3||1|1|1|1|F|Hispanic||9|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|Asian||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504965797|504968348|3|0|2|504719673|4|0|2|500933336|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1791|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|56|Green||2017-01-10|2017-01-10|NaT||||1.8||1|1|1|1|M|Black||9|Yes|Mother|28212|3|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||17|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504970025|504972576|31|0|1|504718076|1|0|2|500939301|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1792|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|491|Green||2013-10-07|2013-10-08|2015-02-11|Child: Changed school/site|Child: Changed school/site||16.1||1|1|1|1|F|Black||9|No|Mother|28217|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||19|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503637911|503639871|31|0|2|503507211|31|0|2|500716290|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1793|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|198|Green||2016-02-09|2016-02-26|2016-09-11|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||6.5||2|2|1|1|M|Black||9|No|Mother|28081|4|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site|Cabarrus County|Match Support|M|White||19|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Enrollment|0|1|1|0|277|60|598|500000170|500012459|504599974|504602385|31|0|1|504579851|1|0|1|500878393|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||6810228174639243761|0
M1794|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|118|Green|Cabarrus County|2016-11-01|2016-11-09|NaT||||3.9||2|2|1|1|M|Black||9|No|Mother|28081|4|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site|Cabarrus County|Match Support|M|White||15|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504599974|504602385|31|0|1|504905469|1|0|1|500922311|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|6810228174639243761|0
M1795|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|378|Green||2016-02-04|2016-02-23|NaT||||12.4||1|1|1|1|M|Black||9|No|Mother|28208|1|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Multi-Race (None of the above)||36|28226||Married|Business: Engineer||0|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|503978163|503980164|31|0|1|504510675|7|0|1|500877548|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||2611337051335117774|0
M1796|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|89|Green||2016-11-16|2016-12-08|NaT||||2.9||1|1|1|1|M|Black||9|No|Mother|28211|3|Two Parent|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504933006|504935557|31|0|1|504708229|1|0|2|500928425|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1797|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|539|Green||2015-09-01|2015-09-15|NaT||||17.7||1|1|1|1|M|Black||9|Yes|GrandMother|28269|1|Grandparents|Less than $10,000|||Y|Yes||School|General Community|Amachi|Match Support|M|White||32|28205|Bachelors Degree|Married|Real Estate: Realtor|28202|6|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504185266|503032503|31|0|1|504213307|1|0|1|500838024|10|2|-2||2|1|500000294|-2||-2|0|4|||17159|12|||1||8998367770661215127|7044657180546140448
M1798|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|809|Green||2014-12-03|2014-12-19|NaT||||26.6||1|1|1|1|M|Black||9|No|Mother|28215|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||34|28269|Bachelors Degree|Living w/ Significant Other|Tech: Sales, Mktg|28117|2|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503663417|503665377|31|0|1|504057497|1|0|1|500800835|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||6407809237813394802|0
M1799|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|616|Green||2014-10-04|2014-10-06|2016-06-13|Volunteer: Moved|Volunteer: Moved||20.2||2|2|1|1|M|Black||9|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||Relative|General Site||Match Support|M|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504033095|504035113|31|0|1|503900507|1|0|1|500780582|10|1|500000296|2128173564|4|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1800|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|M|Black||9|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||Relative|General Site||Match Support|M|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504033095|504035113|31|0|1|504708147|1|0|1|500928418|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M1801|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Pending Match|465|Red||2015-05-11|2015-05-22|2016-08-29|Volunteer: Time constraint|Volunteer: Time constraint||15.3||1|2|1|1|F|Hispanic||9|No|Mother|28212|1|One Parent: Female|$10,000 to $14,999||||Yes||Therapist/Counselor|General Community||Pending Match|F|Hispanic||32|28205|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28203|0|9|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017777|504254967|504257111|3|0|2|504209409|3|0|2|500826456|9|2|-2||4|3||-2|500000294|-2|0|5|||17159|12|||1||9080589164524051479|0
M1802|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|270|Green||2016-05-10|2016-06-10|NaT||||8.9||1|1|1|1|F|Black||9|No|Mother|28206|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||28|28203|Bachelors Degree|Living w/ Significant Other|Finance|28202|0|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504473041|504475315|31|0|2|504582115|1|0|2|500892533|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1||4952249713946979108|5228205320249384837
M1803|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1077|Green||2014-03-26|2014-03-26|NaT||||35.4||1|1|1|1|F|Black||9|Yes|GrandMother|28208|K|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||31|28269||Single|Unemployed||0|0|Recruitment Event|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503530548|503146148|31|0|2|503635342|31|0|2|500756727|10|2|500003586||2|1|500000294|-2||-2|0|10|||7458|9|||1||7679812394383646966|1786514887916898235
M1804|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|687|Green||2014-04-30|2014-05-12|2016-03-29|Child/Family: Time constraints|Child/Family: Time constraints||22.6||1|1|2|2|F|Black||9|No|Mother|28208|K|Two Parent|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||48|28031|Bachelors Degree|Separated|Business: Marketing|28601|16|0|BBBS National Site|Web Link|Big|General Community|Amachi, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500018851|503833932|503835911|31|0|2|503698988|1|0|2|500761753|5|2|-2||4|1||-2|500000294, 500007920, 500011315, 500011316|-2|34|2|||46|2|||1||2611337051335117774|3630529025150538848
M1805|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|167|Green||2015-10-16|2015-11-04|2016-04-19|Child/Family: Moved|Child/Family: Moved||5.5||1|1|1|1|F|Hispanic||9|No|Mother|28213|2|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500011349|504468548|503016895|3|0|2|504297196|1|0|2|500848754|10|1|500000296|2128173564|4|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1806|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|677|Green|Cabarrus County|2015-04-16|2015-04-30|NaT||||22.2||1|1|1|1|F|Black||9|No|Mother|28083|1|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|F|Multi-race (Asian & White)||33|28025|Associate Degree|Married|Business: Marketing|28269|10|0|Self|Self|Big|General Community|Amachi, Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504241299|504243414|31|0|2|504194344|37|0|2|500823537|10|2|500016307||2|1|500016374|-2|500000294, 500016374|-2|34|2|||7464|9|||1|500016374|2437132833506538679|1579263579908564057
M1807|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|120|Green||2016-10-25|2016-11-07|NaT||||3.9||1|1|1|1|F|Black||9|No|Mother|28212|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||32|28269|Masters Degree|Single|Finance|28202|10|1|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504727612|504730049|31|0|2|504822117|31|0|2|500919533|10|2|-2||2|1|500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||7284449467126735125|4127833823859005557
M1808|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|860|Green|PERL 2014-2016|2014-10-15|2014-10-29|NaT||||28.3||1|1|1|1|M|Black||9|No|Mother|28206|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Hispanic||30|28227|Bachelors Degree|Single|Retail: Sales|28105|8|0|Current/Previous Big|Relative|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500008321|503834833|503836805|31|0|1|503968276|3|0|1|500783899|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||17160|11|||1|500014681|421482027904269589|0
M1809|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-18|2016-12-02|NaT||||3.1||1|1|1|1|M|Hispanic||9|No|Father|28212|3|Two Parent|$25,000 to $29,999||||Yes||School|General Site||Match Support|F|White||17|28207|Some High School||Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504929993|504932544|3|0|1|504716201|1|0|2|500929358|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1810|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|544|Green||2015-08-31|2015-09-10|NaT||||17.9||1|1|1|1|M|Black||9|No|Mother|28213|2|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|M|Black||29|28215|Masters Degree|Living w/ Significant Other|Education: Teacher|28206|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503290655|503292479|31|0|1|504326647|31|0|1|500837772|10|2|-2||2|1||-2||-2|0|3|||17159|12|||1||392688197545050058|7380197113384848862
M1811|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|916|Green||2014-08-19|2014-09-03|NaT||||30.1||1|1|1|1|F|Multi-race (Black & Hispanic)||9|No|Mother|28212|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Education: Teacher|28078|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503955220|503838508|38|0|2|503874105|1|0|2|500772805|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||6627885846854295604|7044657180546140448
M1812|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1264|Green||2013-09-09|2013-09-20|NaT||||41.5||1|1|1|1|M|Black||9|No|Mother|28216|3|One Parent: Female|$45,000 to $49,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|Black||35|28216|Some College|Married|Tech: Engineer|28120|0|7|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503366783|503368628|31|0|1|503493458|31|0|1|500709610|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1||2456895876914964961|1202530717971184330
M1813|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|61|Green||2016-12-09|2017-01-05|NaT||||2||1|1|1|1|M|Black||9|No|Mother|28211|3|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504967850|504970401|31|0|1|504718021|1|0|2|500934497|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1814|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|61|Green||2016-12-09|2017-01-05|NaT||||2||1|1|1|1|M|White||9|No|Mother|28211|3|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||17|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504965771|504968322|1|0|1|504718182|1|0|2|500934482|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1815|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-17|2016-12-02|NaT||||3.1||1|1|1|1|M|Multi-race (Black & White)||9|No|Mother|28212|3|Two Parent|$15,000 to $19,999||||Yes||School|General Site||Match Support|M|White||17|28278|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504929976|504932527|36|0|1|504712694|1|0|1|500929156|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1816|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|496|Green||2015-10-16|2015-10-28|NaT||||16.3||1|1|1|1|F|Black||9|No|Mother|28212|2|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504441617|504443869|31|0|2|504296345|1|0|2|500848815|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1817|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|518|Green||2015-10-06|2015-10-06|NaT||||17||1|1|1|1|F|Hispanic||9|No|Mother|28212|2|One Parent: Female|$10,000 to $14,999||||No||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504443588|504444557|3|0|2|504308465|1|0|2|500844549|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1818|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|923|Green||2014-08-12|2014-08-27|NaT||||30.3||1|1|1|1|F|Hispanic||9|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||Relative|General Community||Match Support|F|Hispanic||25|28210|Bachelors Degree|Single|Business: Sales|28277|2|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503496397|503498265|3|0|2|503797696|3|0|2|500772113|10|2|-2||2|1||-2||-2|0|3|||7464|9|||1||2056258660718146620|0
M1819|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|377|Green||2014-10-07|2014-10-22|2015-11-03|Volunteer: Time constraint|Volunteer: Time constraint||12.4||2|2|1|1|M|Black||9|No|Mother|28210|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504029216|504031234|31|0|1|503916972|1|0|1|500781519|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1820|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|334|Green||2015-11-03|2015-11-04|2016-10-03|Child: Changed school/site|Child: Changed school/site||11||2|2|1|1|M|Black||9|No|Mother|28210|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28203|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500011349|504029216|504031234|31|0|1|504307988|1|0|1|500855718|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1821|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|569|Green||2014-11-17|2014-11-17|2016-06-08|Volunteer: Moved|Volunteer: Moved||18.7||1|1|1|1|M|Black||9|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||18|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504030970|504032988|31|0|1|503995921|1|0|2|500796543|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1822|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green|VOL - HSBigs|2016-11-18|2016-11-18|NaT||||3.6||1|1|1|1|F|Black||9|No|Mother|28212|3|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||16|28209|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504929983|504932534|31|0|2|504741735|1|0|2|500929339|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1|500014068|2762897743412756173|0
M1823|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|180|Green||2015-10-15|2015-10-22|2016-04-19|Child/Family: Moved|Child/Family: Moved||5.9||1|1|2|2|M|Hispanic||9|No|Mother|28212|2|Two Parent|Unknown||||Yes||School|General Site||Match Support|M|White||18|28209|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504449801|504452057|3|0|1|504296421|1|0|1|500848539|10|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1824|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|187|Green||2015-10-09|2015-10-21|2016-04-25|Child/Family: Moved|Child/Family: Moved||6.1||1|1|2|2|F|Black||9|No|Mother|28216|2|One Parent: Female|$10,000 to $14,999||||No||School|General Site||Match Support|F|Black||18|28173|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500020908|504443634|504445890|31|0|2|504297141|31|0|2|500846343|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1825|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|661|Green||2013-10-08|2013-10-15|2015-08-07|Volunteer: Moved|Volunteer: Moved||21.7||2|2|1|1|M|Black||9|No|Mother|28211||One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||21|28277|Some High School||Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503644251|503646211|31|0|1|503288713|1|0|1|500717195|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1826|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|503|Green||2015-10-09|2015-10-21|NaT||||16.5||2|2|1|1|M|Black||9|No|Mother|28211||One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|503644251|503646211|31|0|1|504375905|31|0|1|500846324|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1827|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-30|2016-11-30|NaT||||3.2||1|1|1|1|F|Black||9|Yes|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||16|28211|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504956436|504958987|31|0|2|504725140|1|0|2|500931755|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|6084148439133243542
M1828|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|400|Green||2016-01-14|2016-02-01|NaT||||13.1||1|1|2|2|F|Hispanic||9|No|Mother|28212|2|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504576297|504578631|3|0|2|504308458|1|0|2|500872020|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1829|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-17|2016-11-30|NaT||||3.2||1|1|1|1|F|Multi-race (Black & White)||9|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||16|28270|Some High School||Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504942885|504945436|36|0|2|504732009|1|0|2|500929167|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1830|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|637|Green||2013-10-08|2013-10-22|2015-07-21|Volunteer: Moved|Volunteer: Moved||20.9||2|2|1|1|M|Hispanic||9|Yes|Mother|28270|K|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|Match Support|M|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503629828|503631767|3|0|1|503497539|1|0|1|500717190|10|1|500000296|2128173564|4|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1831|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green||2015-10-09|2015-11-11|NaT||||15.8||2|2|1|1|M|Hispanic||9|Yes|Mother|28270|K|One Parent: Female|Unknown|||Y|Yes||School|General Site|Amachi|Match Support|M|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|503629828|503631767|3|0|1|504306008|1|0|1|500846397|10|1|500000296|2128173564|2|1|500000294|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1832|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|48|Green||2016-12-12|2017-01-18|NaT||||1.6||1|1|1|1|F|Black||9|No|Mother|28211|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500021785|504971582|504974133|31|0|2|504708804|1|0|2|500934991|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1833|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-18|2016-11-30|NaT||||3.2||1|1|1|1|M|White||9|No|Mother|28211|3|Two Parent|$30,000 to $34,999||||No||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504932937|504935488|1|0|1|504719691|1|0|2|500929360|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1834|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|707|Yellow|PERL 2014-2016|2015-03-16|2015-03-31|NaT||||23.2||1|1|1|1|M|Black||9|No|GrandMother|28206|3|Grandparents|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||30|28205|Bachelors Degree|Single|Journalist/Media|28202|2|10|Current/Previous Big|Other Big|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|503965808|503967818|31|0|1|504180840|1|0|1|500818934|10|2|-2||2|2|500014681|-2|500000294, 500014681|-2|0|5|||17159|12|||1|500014681|0|0
M1835|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|62|Green||2015-11-12|2015-11-13|2016-01-14|Child: Lost interest|Child: Lost interest||2||1|1|4|4|F|Black||9|No|Mother|28025|2|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|Multi-race (Black & White)||23|28273|Some College|Single|Student: College|28227|0|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500012459|504517488|504519789|31|0|2|503853917|36|0|2|500859286|10|1|500000295|2128212924|4|1||-1|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7464|9|||1||3232906304025417619|0
M1836|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1303|Green||2013-07-30|2013-08-12|NaT||||42.8||1|1|1|1|F|Black||9|Yes|Mother|28215|3|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||47|28269|Associate Degree|Single|Tech: Computer/Programmer|28269|21|0|Big For A Day|Special Event|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503558194|503560069|31|0|2|503527934|31|0|2|500705245|10|2|-2||2|1||-2||-2|0|10|||16422|8|||1||0|1786514887916898235
M1837|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|655|Green||2013-10-09|2013-10-21|2015-08-07|Volunteer: Moved|Volunteer: Moved||21.5||2|2|1|1|M|Black||9|No|Mother|28211|K|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||20|28269|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503661150|503663110|31|0|1|503603498|31|0|1|500717795|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1838|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|509|Green||2015-10-09|2015-10-15|NaT||||16.7||2|2|1|1|M|Black||9|No|Mother|28211|K|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Black||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|503661150|503663110|31|0|1|504297094|31|0|1|500846382|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1839|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|91|Green|VOL - HSBigs|2016-12-05|2016-12-06|NaT||||3||1|1|1|1|M|Black||8|No|Mother|28212|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|Black||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504960078|504962629|31|0|1|504707677|31|0|2|500933245|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1|500014068|2762897743412756173|0
M1840|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|273|Green|PERL 2014-2016|2014-12-02|2014-12-09|2015-09-08|Child/Family: Moved|Child/Family: Moved||9||1|1|2|2|F|Hispanic||8|No|Mother|28025||Other/Unknown|Unknown||||Yes||School|General Site|PERL 2014-2016|Match Support|F|White||31|28025||Married|Retail: Mgt|28025|5|0|Recruitment Event|Workplace Partner|Big|General Site|Cabarrus County, PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500012459|504106167|503675596|3|0|2|504026893|1|0|2|500800151|10|1|500000295|2128212924|4|1|500014681|-1|500014681, 500016374|-1|0|4|||7446|3|||1|500014681|3232906304025417619|0
M1841|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|518|Green||2015-10-06|2015-10-06|NaT||||17||1|1|1|1|F|Black||8|No|Mother|28212|2|Two Parent|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Asian||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504442292|504444548|31|0|2|504375946|4|0|2|500844547|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1842|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|400|Green|Cabarrus County|2016-01-25|2016-02-01|NaT||||13.1||1|1|1|1|F|Multi-race (Hispanic & White)||8|No|Mother|28025||One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|Multi-race (Black & White)||24|28027|Bachelors Degree|Single|Law: Police Officer|28078|1|3|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504533508|504535058|35|0|2|504443510|36|0|2|500875127|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|500016374|643003066716863548|2141487034287122220
M1843|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|984|Green|VOL - Mentoring Hispanic Youth|2014-06-16|2014-06-27|NaT||||32.3||1|1|1|1|F|Hispanic||8|No|Mother|28206|K|One Parent: Female|Unknown||||Yes|Spanish Radio|Media|General Community||Match Support|F|Hispanic||37|28206|Masters Degree|Single|Unknown|28223|1|0|Local Radio|Media|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020753|503575837|503577713|3|0|2|503825634|3|0|2|500766748|10|2|-2||2|1||-2|500014681|-2|7068|1|||7437|1|||1|500011312|392688197545050058|0
M1844|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|133|Red||2016-03-03|2016-03-31|2016-08-11|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.4||1|1|2|2|M|Black||8|No|Mother|28027|2|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|Black||58|28215|Some College|Divorced|Customer Service||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020753|504487104|504489379|31|0|1|502924751|31|0|1|500882883|10|2|-2||4|3|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|34|2|||7464|9|||1||3232906304025417619|2447619215802866303
M1845|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|47|Green||2017-01-18|2017-01-19|NaT||||1.5||1|1|1|1|F|Hispanic||8|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||16|28205|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504998024|505000584|3|0|2|504718378|1|0|2|500940767|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1846|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|47|Green||2017-01-18|2017-01-19|NaT||||1.5||1|1|1|1|F|Hispanic||8|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504998017|505000577|3|0|2|504714248|1|0|2|500940762|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1847|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1287|Green||2013-08-16|2013-08-28|NaT||||42.3||1|1|1|1|F|Black||8|No|Mother|28203|1|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||40|28204|Masters Degree|Single|Finance: Banking|28212|5|7|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503579909|502958068|31|0|2|503552956|1|0|2|500707000|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||7960300212314874874|0
M1848|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|872|Green||2014-10-14|2014-10-17|NaT||||28.6||1|1|1|1|F|Black||8|Yes|Mother|28211|K|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||26|28277|Bachelors Degree|Single|Business|28273|1|9|Local Print|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503798824|503800801|31|0|2|503895001|1|0|2|500783536|10|2|-2||2|1|500000294|-2||-2|0|10|||7439|1|||1||7807202941877299922|0
M1849|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|112|Green||2016-11-15|2016-11-15|NaT||||3.7||1|1|1|1|M|Black||8|No|Mother|28211|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|M|White||17|28211|Some High School||Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504930097|504932648|31|0|1|504707501|1|0|1|500927976|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1850|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|573|Green||2014-11-11|2014-11-18|2016-06-13|Volunteer: Moved|Volunteer: Moved||18.8||1|1|1|1|M|Black||8|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504103356|504105390|31|0|1|503896267|1|0|2|500794446|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1851|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|553|Green||2014-01-09|2014-01-30|2015-08-06|Child/Family: Moved|Child/Family: Moved||18.2||1|1|1|1|F|Black||8|No|Mother|28203|1|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||33|28277|Bachelors Degree|Single|Insurance|28277|3|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500015820|503554921|503556796|31|0|2|503556149|1|0|2|500742082|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1||6095563712459522926|0
M1852|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|922|Green||2014-08-12|2014-08-28|NaT||||30.3||2|2|1|1|F|Black||8|No|Mother|28216|2|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Asian||31|28202|Bachelors Degree|Single|Business: Sales|28217|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503654738|500740560|31|0|2|503853843|4|0|2|500772115|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1||3664007741235143067|0
M1853|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-17|2016-12-02|NaT||||3.1||1|1|1|1|M|Black||8|Yes|Mother|28227|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||17|28207|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504931611|504934162|31|0|1|504709361|1|0|2|500929164|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1854|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|341|Green||2015-09-29|2015-10-28|2016-10-03|Child: Changed school/site|Child: Changed school/site||11.2||1|1|2|2|M|Black||8|No|Mother|28212||One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500022905|504442313|504444569|31|0|1|504297082|1|0|1|500843033|10|1|500000296|2128173564|4|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1855|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-28|2016-12-02|NaT||||3.1||1|1|1|1|M|Black||8|No|Mother|28211|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504037433|504039451|31|0|1|504722559|1|0|2|500930970|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|862536831521836203
M1856|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|232|Red||2015-03-24|2015-04-14|2015-12-02|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.6||1|1|2|2|M|Black||8|No|Mother|28208|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|M|Multi-race (Black & White)||29|28216|Doctor of Medicine (MD)|Married|Retired||8|0|AA Task Force|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500013781|503856172|503858166|31|0|1|503961801|36|0|1|500820145|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|3|||9223|3|||1||2762897743412756173|6397220780367831607
M1857|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|644|Green||2013-10-29|2013-11-01|2015-08-07|Volunteer: Moved|Volunteer: Moved||21.2||2|2|1|1|M|Hispanic||8|No|Mother|28270|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503644282|503646242|3|0|1|503521705|1|0|2|500724454|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1858|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|508|Green||2015-10-15|2015-10-16|NaT||||16.7||2|2|1|1|M|Hispanic||8|No|Mother|28270|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|503644282|503646242|3|0|1|504301111|1|0|1|500848542|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1859|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|92|Green|Cabarrus County|2016-11-22|2016-12-05|NaT||||3||1|1|2|2|M|Black||8|Yes|Mother|28025|3|One Parent: Female|Less than $10,000|||Y|No|BBBS National Site|Web Link|General Community|Amachi, Cabarrus County|Match Support|M|Asian||27|28075|Bachelors Degree|Single|Finance: Banking|28202|3|0|Local Print|Media|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|503617871|503619748|31|0|1|503786945|4|0|1|500930374|10|2|500016307||2|1|500000294, 500016374|-2|500014681, 500016374|-2|34|2|||7439|1|||1|500016374|0|2763237020791144915
M1860|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|61|Green||2016-12-12|2017-01-05|NaT||||2||1|1|1|1|M|Hispanic||8|No|Mother|28212|3|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||16|28209|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504971614|504974165|3|0|1|504708240|1|0|2|500934860|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1861|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|48|Green||2017-01-18|2017-01-18|NaT||||1.6||1|1|1|1|M|Some Other Race||8|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|505001625|505004185|41|0|1|504716181|1|0|2|500940772|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1862|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|135|Green|Cabarrus County|2016-10-11|2016-10-23|NaT||||4.4||1|1|1|1|F|White||8|No|GrandMother|28025|3|Grandparents|$15,000 to $19,999||||Yes||Self|General Community|Cabarrus County|Match Support|F|White||51|28081|Associate Degree|Married|Medical: Nurse|28025|87|11|Local TV|Media|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504819428|504821927|1|0|2|504805078|1|0|2|500914390|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7438|1|||1|500016374|5064856656261650513|0
M1863|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|202|Yellow||2016-03-03|2016-03-11|2016-09-29|Volunteer: Time constraint|Volunteer: Time constraint||6.6||1|1|5|5|F|Black||8|No|GrandMother|28025|2|Grandparents|Less than $10,000|||Y|Yes||School|General Site|Cabarrus County|RTBM|F|White||44|28075|Bachelors Degree|Married|Tech: Computer/Programmer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500012459|504579544|504581878|31|0|2|502143796|1|0|2|500882802|7|1|500000295|2128212924|4|2|500016374|-1|500007920, 500011315, 500011316, 500016374|-1|0|4|||7496|10|||1||3232906304025417619|0
M1864|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|576|Green||2014-11-09|2014-11-10|2016-06-08|Volunteer: Moved|Volunteer: Moved||18.9||1|1|1|1|F|White||8|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504101750|504103784|1|0|2|503898526|1|0|2|500793661|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1865|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|205|Green||2015-08-07|2015-08-31|2016-03-23|Child/Family: Moved|Child/Family: Moved||6.7||1|1|1|1|M|Black||8|Yes|Mother|28216|2|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|White||28|28269|Bachelors Degree|Single|Finance: Banking|28025|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500017732|503805008|503806985|31|0|1|504322860|1|0|1|500835488|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||7284449467126735125|0
M1866|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|99|Green|VOL - HSBigs|2016-11-18|2016-11-28|NaT||||3.3||1|1|1|1|F|Hispanic||8|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||16|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504934159|504936710|3|0|2|504709318|1|0|2|500929367|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1|500014068|2762897743412756173|0
M1867|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|608|Green||2014-10-07|2014-10-14|2016-06-13|Volunteer: Moved|Volunteer: Moved||20||2|2|1|1|F|Black||8|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504029245|504031263|31|0|2|503907342|1|0|2|500781518|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1868|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||2|2|1|1|F|Black||8|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Black||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504029245|504031263|31|0|2|504719766|31|0|2|500929321|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1869|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|91|Green||2016-12-06|2016-12-06|NaT||||3||1|1|1|1|M|Black||8|No|Mother|28212|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|M|White||16|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504956449|504959000|31|0|1|504712902|1|0|1|500933319|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1870|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green||2016-12-05|2016-12-05|NaT||||3||1|1|1|1|F|Hispanic||8|No|Mother|28218|3|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504960064|504962615|3|0|2|504719639|1|0|2|500932930|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1871|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|665|Green||2013-10-08|2013-10-11|2015-08-07|Volunteer: Moved|Volunteer: Moved||21.8||2|2|1|1|F|Hispanic||8|No|Mother|28203|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28173||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503644208|503646168|3|0|2|503540957|1|0|2|500717203|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1872|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|348|Green||2015-10-09|2015-10-21|2016-10-03|Child: Changed school/site|Child: Changed school/site||11.4||2|2|2|2|F|Hispanic||8|No|Mother|28203|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|503644208|503646168|3|0|2|504301129|1|0|2|500846345|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1873|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|426|Green||2014-09-29|2014-09-30|2015-11-30|Child/Family: Moved|Child/Family: Moved||14||1|1|1|1|F|Black||8|No|Step-Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500020909|504033059|504035077|31|0|2|503898570|1|0|2|500778743|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1874|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||1|1|1|1|M|Hispanic||8|No|Mother|28211|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||16|28209|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504933160|504935711|3|0|1|504709325|1|0|2|500928440|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1875|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|77|Green|Cabarrus County|2016-12-06|2016-12-20|NaT||||2.5||1|1|1|1|F|Black||8|No|Mother|28083|3|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|Cabarrus County|Match Support|F|Black||19|28025|Some College|Single|Business|28025|0|1|Current/Previous Big|Other Big|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504966805|504969356|31|0|2|504843117|31|0|2|500933679|10|1|500000295|2128232374|2|1|500016374|-1|500016374|-1|0|4|||17159|12|||1|500016374|2043334928777030191|0
M1876|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|95|Green||2016-11-17|2016-12-02|NaT||||3.1||1|1|1|1|F|Hispanic||8|No|Mother|28212|3|Two Parent|Less than $10,000||||Yes||School|General Site||Match Support|F|White||16|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504933392|504935943|3|0|2|504707250|1|0|2|500929147|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1877|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|298|Green||2014-10-30|2014-11-21|2015-09-15|Child/Family: Moved|Child/Family: Moved||9.8||1|1|1|1|F|Multi-race (Black & White)||8|Yes|Aunt|28027||Two Parent|Unknown||||Yes||School|General Site||Match Support|F|Black||56|28027||Married|Retail: Mgt||0|3|Recruitment Event|Workplace Partner|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|1|0|1|0|277|60|598|500000170|500012459|504073275|504075304|36|0|2|504032411|31|0|2|500790059|10|1|500000295|2128212924|4|1||-1|500007920, 500011315, 500011316, 500016374|-1|0|4|||7446|3|||1||3232906304025417619|0
M1878|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|32|Green||2017-01-26|2017-02-03|NaT||||1.1||1|1|1|1|F|Hispanic||8|No|Mother|28212|3|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|Asian||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|505011025|505013585|3|0|2|504707532|4|0|2|500942145|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1879|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|419|Yellow||2014-05-06|2014-05-16|2015-07-09|Volunteer: Moved|Volunteer: Moved||13.8||2|2|1|1|F|Black||8|Yes|Mother|28216|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||33|28202|Masters Degree|Single|Consultant|28202|0|1|Man Up Campaign|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|503717075|503719040|31|0|2|503842851|1|0|2|500762275|10|2|-2||4|2||-2||-2|0|10|||17101|1|||1||1653226628427425023|0
M1880|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|477|Green||2015-11-02|2015-11-16|NaT||||15.7||2|2|1|1|F|Black||8|Yes|Mother|28216|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Business|28217|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503717075|503719040|31|0|2|504270682|1|0|2|500854847|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||1653226628427425023|0
M1881|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|198|Green||2016-03-11|2016-03-15|2016-09-29|Child/Family: Moved|Child/Family: Moved||6.5||1|1|2|2|F|Black||8|No|Mother|28025|2|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|Cabarrus County|Match Support|F|Hispanic||17|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504652697|504655124|31|0|2|504579805|3|0|2|500884397|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||9080589164524051479|0
M1882|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|213|Green||2016-02-23|2016-02-29|2016-09-29|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||7||2|2|1|1|F|Black||8|Yes|Mother|28027|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Site|Cabarrus County|Match Support|F|White||19|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504599957|504602368|31|0|2|504579744|1|0|2|500881126|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||6810228174639243761|0
M1883|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|118|Green|Cabarrus County|2016-10-17|2016-11-09|NaT||||3.9||2|2|1|1|F|Black||8|Yes|Mother|28027|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Site|Cabarrus County|Match Support|F|White||17|28027|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504599957|504602368|31|0|2|504871177|1|0|2|500916295|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||0|4|||1|500016374|6810228174639243761|0
M1884|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|315|Green|Cabarrus County|2016-04-05|2016-04-26|NaT||||10.3||1|1|1|1|M|Black||8|No|Mother|28027|2|One Parent: Female|$20,000 to $24,999|||Y|Yes||Therapist/Counselor|General Community|Cabarrus County|Match Support|M|White||28|28083|Some College|Married|Business||10|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504612286|504614697|31|0|1|504634827|1|0|1|500887835|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|5|||7464|9|||1|500016374|3664007741235143067|3409063327463232933
M1885|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|246|Green||2015-01-23|2015-01-29|2015-10-02|Volunteer: Time constraint|Volunteer: Time constraint||8.1||2|2|1|1|F|Black||8||Mother|28025||One Parent: Female|Unknown||||Yes||School|General Site|Cabarrus County|Match Support|F|White||19|28027|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500002335|504106116|504108150|31|0|2|504043276|1|0|2|500809861|10|1|500000296|2128173571|4|1|500016374|-1||-1|0|4|||0|4|||1||5208542183136337346|0
M1886|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|375|Green|Cabarrus County|2016-02-18|2016-02-26|NaT||||12.3||2|2|1|1|F|Black||8||Mother|28025||One Parent: Female|Unknown||||Yes||School|General Site|Cabarrus County|Match Support|F|White||18|28027|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504106116|504108150|31|0|2|504579862|1|0|2|500880037|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|5208542183136337346|0
M1887|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|374|Green||2014-09-29|2014-09-30|2015-10-09|Child: Changed school/site|Child: Changed school/site||12.3||1|1|2|2|M|Hispanic||8|No|Mother|28211|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28036|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504035892|504037910|3|0|1|503905466|1|0|1|500778750|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1888|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|357|Green||2014-11-11|2014-11-11|2015-11-03|Child: Changed school/site|Child: Changed school/site||11.7||1|1|3|3|M|Hispanic||8|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||19|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504095796|504097830|3|0|1|503905482|1|0|1|500794472|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1889|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|206|Green||2015-06-19|2015-07-17|2016-02-08|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||6.8||1|1|1|1|M|Black||8|No|Mother|28273|1|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|Black||54|28278|Some College|Married|Business: Sales|28205|2|8|Igniting Breakfast|Special Event|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500020990|503902854|503904854|31|0|1|504273752|31|0|1|500830786|5|2|-2||4|1||-2||-2|34|2|||17266|8|||1||7508998544817094399|6156547733130613405
M1890|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|368|Green||2014-10-04|2014-10-06|2015-10-09|Child: Changed school/site|Child: Changed school/site||12.1||1|1|2|2|M|Black||8|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504033104|504035122|31|0|1|503907262|1|0|1|500780583|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1891|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|401|Green||2016-01-12|2016-01-31|NaT||||13.2||1|1|1|1|M|Black||8|Yes|Mother|28215|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|M|White||30|28205|Bachelors Degree||Arts, Entertainment, Sports|28206|0|3|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504231851|504233090|31|0|1|503291779|1|0|1|500871254|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||6077912216232501082|7327400833679234452
M1892|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|98|Green||2016-11-18|2016-11-29|NaT||||3.2||1|1|1|1|M|Black||8|No|Father|28212|3|One Parent: Male|Unknown||||Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022908|504930076|504932627|31|0|1|504709344|1|0|2|500929337|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1893|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|505|Green||2015-10-06|2015-10-19|NaT||||16.6||1|1|1|1|F|Black||8|No|Mother|28203|2|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||24|28202|Masters Degree|Single|Education: Teacher|28208|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504388144|504390375|31|0|2|504365599|1|0|2|500844802|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||8568001799025358453|2876415545463317777
M1894|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|516|Green||2014-05-22|2014-05-31|2015-10-29|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17||1|1|1|1|M|Multi-race (Black & White)||8|No|Mother|28115|2|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|White||45|28031|Bachelors Degree|Married|Real Estate: Realtor|28031|20|0|Local Print|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503572810|503078467|36|0|1|503785317|1|0|1|500764166|5|2|-2||4|1||-2||-2|0|10|||7439|1|||1||7857548027029642592|8690133977366715726
M1895|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|322|Green||2016-03-14|2016-04-19|NaT||||10.6||1|1|1|1|F|Black||8|No|Mother|28217|1|One Parent: Female|$25,000 to $29,999|||Y|No||Self|General Community||Match Support|F|White||28|28210|Masters Degree|Single|Finance: Accountant|28210|0|3|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504532539|504534872|31|0|2|504467958|1|0|2|500884487|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||0|1136572582102976964
M1896|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|475|Green||2015-10-16|2015-10-28|2017-02-14|Volunteer: Health|Volunteer: Health||15.6||2|2|1|1|F|Black||8|No|Mother|28211|2|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Black||17|28262|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500022909|504468571|504065687|31|0|2|504301055|31|0|2|500848763|10|1|500000296|2128173564|4|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1897|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|21|Green|VOL - HSBigs|2017-02-14|2017-02-14|NaT||||0.7||2|2|1|1|F|Black||8|No|Mother|28211|2|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504468571|504065687|31|0|2|504707239|1|0|2|500946313|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|4|||0|4|||1|500014068|2762897743412756173|0
M1898|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|85|Green||2016-12-06|2016-12-12|NaT||||2.8||1|1|1|1|F|Black||8|No|Mother|28217|3|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||22|28117||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504886770|504889290|31|0|2|504771529|1|0|2|500933349|10|1|500000295|2128207319|2|1||-1||-1|0|4|||46|2|||1||3935539763241716148|0
M1899|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|130|Green||2016-10-07|2016-10-28|NaT||||4.3||1|1|2|2|M|Multi-Race (None of the above)||8|No|Mother|28031|3|Two Parent|$30,000 to $34,999||||No||School|General Site||Match Support|M|Black||21|28035|Some College|Single|Student: College||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504883829|504886349|7|0|1|504629735|31|0|1|500913774|10|1|500000295|2128173570|2|1||-1||-1|0|4|||7464|9|||1||8034889377453131101|7489588860826267930
M1900|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|599|Green||2015-06-18|2015-07-17|NaT||||19.7||1|1|1|1|M|Black||8|No|Mother|28202|1|One Parent: Female|$25,000 to $29,999||||Yes||School|General Community||Match Support|M|White||25|28210|Bachelors Degree|Single|Business: Sales|29172|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503804124|503712061|31|0|1|504284484|1|0|1|500830694|10|2|-2||2|1||-2||-2|0|4|||17159|12|||1||6368218764956286027|5056473444237941296
M1901|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|111|Green|Cabarrus County|2016-11-16|2016-11-16|NaT||||3.6||1|1|1|1|F|White||8|No|Mother|28081|3|One Parent: Female|Less than $10,000||||Yes||Relative|General Community|Cabarrus County|Match Support|F|White||24|28027|Bachelors Degree|Single|Business|28205|0|3|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500020753|504915869|504864541|1|0|2|504933506|1|0|2|500928289|10|2|-2||2|1|500016374|-2|500016374|-2|0|3|||7464|9|||1|500016374|6810228174639243761|2036270106764562772
M1902|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|189|Green||2016-08-22|2016-08-30|NaT||||6.2||1|1|1|1|M|Black||8|No|Mother|28208|2|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||24|28209|Bachelors Degree|Single|Finance: Accountant|28209|0|1|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504348389|504350613|31|0|1|504667599|1|0|1|500904262|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||3038247238543299436|7795805164050330858
M1903|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|401|Green||2016-01-08|2016-01-31|NaT||||13.2||1|1|2|2|F|Black||8|Yes|Mother|28262|2|One Parent: Female|$25,000 to $29,999|||Y|Yes||Relative|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504538972|504402454|31|0|2|502171015|31|0|2|500870863|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|3|||7496|10|||1||2417657944362725638|6156547733130613405
M1904|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|224|Green||2016-06-02|2016-06-16|2017-01-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.4||1|1|2|2|M|Black||8|Yes|Mother|28262|2|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|Multi-race (Black & White)||29|28216|Doctor of Medicine (MD)|Married|Retired||8|0|AA Task Force|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500021785|504400213|504402454|31|0|1|503961801|36|0|1|500895512|5|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|34|2|||9223|3|||1||2417657944362725638|6156547733130613405
M1905|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|393|Green||2014-10-29|2014-11-03|2015-12-01|Child/Family: Moved|Child/Family: Moved||12.9||1|1|1|1|F|Black||8|Yes|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504081829|504083858|31|0|2|503916445|1|0|2|500789776|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1906|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|280|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-23|2016-05-31|NaT||||9.2||1|1|1|1|M|Black||8|No|Mother|28213|1|One Parent: Female|$40,000 to $44,999||||No||School|General Community||Match Support|M|White||27|28203|Bachelors Degree||Transport: Driver|28105|2|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504155409|504157461|31|0|1|504606544|1|0|1|500894080|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|500007920, 500011315, 500011316|0|5439372922340750169
M1907|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|563|Green||2014-11-04|2014-11-18|2016-06-03|Volunteer: Moved|Volunteer: Moved||18.5||1|1|1|1|M|Asian||8|No|Mother|28212||One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504041991|504044009|4|0|1|503898591|1|0|2|500791891|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1908|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|109|Green||2016-11-18|2016-11-18|NaT||||3.6||1|1|1|1|M|Black||8|No|Mother|28212|3|One Parent: Female|Less than $10,000||||No||School|General Site||Match Support|F|White||17|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504933110|504935661|31|0|1|504719709|1|0|2|500929340|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1909|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|622|Green||2014-09-29|2014-09-30|2016-06-13|Volunteer: Moved|Volunteer: Moved||20.4||2|2|1|1|F|Hispanic||8|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|Asian||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504033052|504035070|3|0|2|503896236|4|0|2|500778748|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1910|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|F|Hispanic||8|No|Mother|28212|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504033052|504035070|3|0|2|504732663|1|0|2|500928447|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1911|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|97|Green||2016-11-30|2016-11-30|NaT||||3.2||1|1|1|1|F|Black||8|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999||||Yes||Relative|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504956421|504958972|31|0|2|504727760|1|0|2|500931748|10|1|500000296|2128173564|2|1||-1||-1|0|3|||0|4|||1||2762897743412756173|0
M1912|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|401|Green||2015-07-26|2015-07-26|2016-08-30|Child/Family: Moved|Child/Family: Moved||13.2||1|1|1|1|F|Black||8|No|Mother|28214|1|One Parent: Female|$45,000 to $49,999||||Yes||School|General Community||Match Support|F|White||25|28269|Bachelors Degree|Single|Law|28277|0|7|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|504272839|504275039|31|0|2|504114967|1|0|2|500834459|10|2|-2||4|1||-2||-2|0|4|||46|2|||1||0|2806833304218536184
M1913|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|119|Green|Cabarrus County|2016-11-04|2016-11-08|NaT||||3.9||2|2|2|2|F|Black||8|No|Mother|28025|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Site|Cabarrus County|Match Support|F|Hispanic||18|28027|Some High School||Student: College||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504629014|504631425|31|0|2|504619516|3|0|2|500924799|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|6898335769881586649|0
M1914|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|235|Green||2016-02-18|2016-03-03|2016-10-24|Child: Changed school/site|Child: Changed school/site||7.7||2|2|2|2|F|Black||8|No|Mother|28025|2|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Site|Cabarrus County|Match Support|F|Hispanic||18|28027|Some High School||Student: College||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504629014|504631425|31|0|2|504619516|3|0|2|500880074|10|1|500000296|2128173571|4|1|500016374|-1|500016374|-1|0|4|||7464|9|||1||6898335769881586649|0
M1915|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|61|Green||2016-12-07|2017-01-05|NaT||||2||1|1|1|1|M|Asian||8|No|Mother|28211|3|Two Parent|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||17|28226||Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504967881|504970432|4|0|1|504707461|1|0|2|500933957|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1916|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|31|Green|Cabarrus County|2017-01-27|2017-02-04|NaT||||1||1|1|1|1|F|Black||8|No|Mother|28027|2|One Parent: Female|$30,000 to $34,999||||No||Therapist/Counselor|General Community|Cabarrus County|Match Support|F|White||35|28269|Bachelors Degree|Married|Business: Sales|30097|9|3|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504952245|504954796|31|0|2|504757125|1|0|2|500942600|10|2|500016307||2|1|500016374|-2|500016374|-2|0|5|||7464|9|||1|500016374|3575183301237417432|4698448699835736001
M1917|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|21|Green||2017-02-07|2017-02-14|NaT||||0.7||1|1|1|1|F|Black||8|No|Mother|28212|3|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|505022089|505024657|31|0|2|504741631|1|0|2|500945080|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1918|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|637|Green||2013-10-29|2013-11-08|2015-08-07|Volunteer: Moved|Volunteer: Moved||20.9||2|2|1|1|F|Hispanic||8|No|Mother|28105|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|503661106|503663066|3|0|2|503608284|1|0|2|500724456|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1919|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|348|Green||2015-10-09|2015-10-21|2016-10-03|Child: Changed school/site|Child: Changed school/site||11.4||2|2|2|2|F|Hispanic||8|No|Mother|28105|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500022905|503661106|503663066|3|0|2|504303240|1|0|2|500846360|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1920|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|85|Green|Cabarrus County|2016-11-22|2016-12-12|NaT||||2.8||1|1|1|1|F|Black||8|No|Mother|28027|3|One Parent: Female|$15,000 to $19,999||||Yes||School|General Community|Cabarrus County|Match Support|F|White||51|28027|Masters Degree|Married|Business|28213|1|10|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504937124|504939686|31|0|2|504828127|1|0|2|500930334|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||17159|12|||1|500016374|1550830965009450729|0
M1921|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|488|Green||2015-10-20|2015-11-05|NaT||||16||1|1|1|1|M|Black||8|No|Mother|28269|K|One Parent: Female|$30,000 to $34,999||||Yes||School|General Community||Match Support|M|White||27|28204|Bachelors Degree|Married|Business: Mgt, Admin|28117|0|6|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504275417|504277617|31|0|1|504249590|1|0|1|500849815|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||7458247995093008174|4148565630505427365
M1922|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|397|Red||2015-02-10|2015-03-18|2016-04-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13||1|1|1|1|M|Multi-race (Black & Hispanic)||8|No|Mother|28105|K|One Parent: Female|$25,000 to $29,999|||Y|Yes|Radio|Media|General Community|VOL - Mentoring Hispanic Youth|Enrollment|M|White||30|28270|Some College|Single|Business: Marketing||5|0|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503781255|503783232|38|0|1|504179316|1|0|1|500813063|5|2|-2||4|3|500011312|-2||-2|55|1|||7438|1|||1||7134583514356134698|9044147131226222704
M1923|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2017-01-17|2017-01-30|NaT||||1.2||1|1|1|1|F|Black||8|No|Mother|28208|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||54|28273|Bachelors Degree|Single|Tech: Research/Design|6082|7|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504917122|504919642|31|0|2|504453155|31|0|2|500940412|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1||3935539763241716148|7044657180546140448
M1924|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|820|Green||2014-11-19|2014-12-08|NaT||||26.9||1|1|1|1|F|Black||8|Yes|Mother|28262|K|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|White||40|28205|Bachelors Degree|Divorced|Law|28204|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|503993975|503969639|31|0|2|503947272|1|0|2|500797389|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1||6627885846854295604|6619197389800008587
M1925|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|351|Green||2014-11-09|2014-11-10|2015-10-27|Child: Changed school/site|Child: Changed school/site||11.5||1|1|2|2|M|Black||8|Yes|Mother|28232|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28207|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504095814|504097848|31|0|1|503901733|1|0|2|500793662|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1926|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2017-01-12|2017-01-30|NaT||||1.2||1|1|1|1|M|Black||8|Yes|Mother|28217|1|One Parent: Female|$30,000 to $34,999||||No||School|General Community||Match Support|M|White||25|28209|Bachelors Degree|Single|Finance: Accountant|28205|3|3|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504456510|504458770|31|0|1|504829731|1|0|1|500939755|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||0|5597049740348738
M1927|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|139|Green||2016-09-21|2016-10-19|NaT||||4.6||1|1|1|1|M|Black||8|No|Aunt|28208||Other Relative|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||34|28205|Bachelors Degree|Separated|Business: Sales|28273|3|1|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|503862846|502431630|31|0|1|504765492|1|0|1|500909169|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||0|0
M1928|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|334|Green||2016-03-09|2016-04-07|NaT||||11||1|1|1|1|F|Black||8|No|Mother|28262|1|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||43|28117|Bachelors Degree|Married|Insurance|2114|14|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020752|504357786|504360012|31|0|2|504163106|1|0|2|500883845|10|2|-2||3|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1||7102230088759381237|5081726734274569781
M1929|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|569|Green||2014-11-04|2014-11-17|2016-06-08|Volunteer: Moved|Volunteer: Moved||18.7||1|1|1|1|M|Black||8|Yes|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504041716|504043734|31|0|1|503916375|1|0|2|500791873|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1930|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|196|Green||2016-04-01|2016-04-11|2016-10-24|Child: Changed school/site|Child: Changed school/site||6.4||1|1|2|2|M|Hispanic||8|No|Mother|28078|K|One Parent: Female|Unknown||||Yes||School|General Site|Amachi|Match Support|M|Black||20|28035|||Student: College||0|0|Self|Self|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500015820|504579602|504581936|3|0|1|504634278|31|0|1|500887470|10|1|500000295|2128173570|4|1|500000294|-1||-1|0|4|||7464|9|||1||8034889377453131101|0
M1931|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|832|Green|Cabarrus County|2014-10-22|2014-11-26|NaT||||27.3||1|1|2|2|F|Black||8|No|Mother|28083|2|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||69|28027||Married|Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|504069856|504071884|31|0|2|502591360|31|0|2|500786507|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|0|0
M1932|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|200|Green|Cabarrus County|2016-08-11|2016-08-19|NaT||||6.6||1|1|1|1|M|Multi-race (Hispanic & White)||8|No|GrandMother|28027|2|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Site|Cabarrus County|Match Support|M|White||36|28027||Married|Medical: Doctor, Provider|28027|0|6|Recruitment Event|Neighbor/Friend|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504026699|504028717|35|0|1|504659125|1|0|1|500903059|10|1|500000295|2128212924|2|1|500016374|-1|500016374|-1|0|4|||7459|10|||1|500016374|3232906304025417619|0
M1933|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|515|Green||2015-10-09|2015-10-09|NaT||||16.9||1|1|1|1|F|Black||8|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504449794|504452050|31|0|2|504303177|1|0|2|500846140|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1934|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|475|Green||2015-11-16|2015-11-18|NaT||||15.6||1|1|1|1|M|Black||8|No|Mother|28212|1|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site||Match Support|F|White||18|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504447302|504444540|31|0|1|504307845|1|0|2|500860347|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1935|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|731|Red|Cabarrus County|2014-11-10|2014-11-21|2016-11-21|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||24||1|1|1|1|F|Black||8|Yes|GrandMother|28083||One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||25|28081||Single|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Enrollment|1|0|1|0|277|60|598|500000170|500022817|504096330|503587420|31|0|2|503992956|1|0|2|500794009|10|2|500016307||4|3|500000294, 500016374|-2|500016374|-2|0|10|||46|2|||1|500016374|6810228174639243761|0
M1936|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|731|Red|Cabarrus County|2014-10-30|2014-11-21|2016-11-21|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||24||1|1|1|1|F|Black||8|Yes|GrandMother|28083||One Parent: Female|Unknown|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||28|28027|Masters Degree|Single|Human Services: Social Worker|28202|1|1|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500022817|504096289|503587420|31|0|2|503776419|31|0|2|500790461|10|2|500016307||4|3|500016374|-2|500014681, 500016374|-2|0|10|||7464|9|||1|500016374|6810228174639243761|0
M1937|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|866|Green||2014-10-15|2014-10-23|NaT||||28.5||1|1|1|1|F|Black||8|No|Mother|28213|K|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||27|28269|Some College|Single|Business|28269|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|504044312|504046330|31|0|2|503862152|31|0|2|500783874|10|2|-2||2|1||-2||-2|0|10|||46|2|||1||7458247995093008174|6368850787260662385
M1938|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|361|Green||2015-10-09|2015-10-09|2016-10-04|Child: Changed school/site|Child: Changed school/site||11.9||1|1|1|1|M|Black||8|Yes|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|M|Black||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|RTBM|0|1|1|0|277|60|598|500000170|500011349|504029267|504031285|31|0|1|504375960|31|0|1|500846132|10|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||7554307376683929204|0
M1939|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|365|Green|PERL 2014-2016, Cabarrus County|2016-02-29|2016-03-07|NaT||||12||1|1|1|1|M|Hispanic||8|No|Foster Parent|28078|1|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||50|28036||Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504433829|504436084|3|0|1|504470539|1|0|1|500882069|10|2|500016307||2|1|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|5|||46|2|||1|500014681, 500016374|0|7470110347975227693
M1940|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|497|Green||2015-10-09|2015-10-27|NaT||||16.3||1|1|1|1|F|Hispanic||8|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||18|28211|High School Graduate|Single|Student: College||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504443697|504443839|3|0|2|504307612|1|0|2|500846368|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1941|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|189|Green||2016-08-22|2016-08-30|NaT||||6.2||1|1|1|1|M|Black||8|No|Mother|28262|K|One Parent: Female|$35,000 to $39,999|||Y|No||Self|General Community||Match Support|M|White||24|28202|Bachelors Degree|Single|Finance: Banking||0|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504180621|504182730|31|0|1|504624656|1|0|1|500904258|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1||6933349951274183958|2029142410245134798
M1942|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|875|Green||2014-06-12|2014-06-27|2016-11-18|Volunteer: Moved|Volunteer: Moved||28.7||1|1|1|1|F|Black||8|No|Mother|28212|2|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||RTBM|F|Black||63|28213||Single|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|503774486|503776463|31|0|2|503792812|31|0|2|500766439|7|2|-2||4|1||-2||-2|34|2|||7464|9|||1||314687390558932914|4127833823859005557
M1943|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|97|Green||2014-10-07|2014-10-21|2015-01-26|Child/Family: Moved|Child/Family: Moved||3.2||1|1|2|2|F|Hispanic||8|Yes|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||18|28222|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500019116|504049133|504051157|3|0|2|503907282|1|0|2|500781527|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1944|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|175|Green||2014-11-09|2014-11-17|2015-05-11|Child/Family: Moved|Child/Family: Moved||5.7||1|1|2|2|F|White||8|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28209||Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504095817|504097851|1|0|2|503995722|1|0|2|500793665|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1945|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|141|Green||2016-10-07|2016-10-17|NaT||||4.6||1|1|1|1|M|Black||8|No|Mother|28031|1|Two Parent|$30,000 to $34,999||||No||School|General Site||Match Support|M|White||37|28273|Bachelors Degree|Married|Tech: Management|28031|4|0|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504834879|504837381|31|0|1|504666284|1|0|1|500913775|10|1|500000295|2128173570|2|1||-1||-1|0|4|||18809|8|||1||8034889377453131101|0
M1946|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|173|Green||2016-09-02|2016-09-15|NaT||||5.7||1|1|1|1|M|Black||7|No|Mother|28208|1|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||27|28214|Masters Degree|Single|Business: Marketing|28208|1|0|Current/Previous Big|Relative|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504303891|504306109|31|0|1|504553488|1|0|1|500906091|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||17160|11|||1||0|7044657180546140448
M1947|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|2|2|M|White||7|No|Mother|28212|K|Two Parent|$50,000 to $59,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Multi-Race (None of the above)||18|29708|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504524465|504526796|1|0|1|504438216|7|0|2|500929201|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1948|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|314|Green|VOL - HSBigs|2015-11-19|2015-12-01|2016-10-10|Child: Changed school/site|Child: Changed school/site||10.3||2|2|2|2|M|White||7|No|Mother|28212|K|Two Parent|$50,000 to $59,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Multi-Race (None of the above)||18|29708|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500022905|504524465|504526796|1|0|1|504438216|7|0|2|500861403|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1|500014068|2762897743412756173|0
M1949|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|574|Green||2014-11-11|2014-11-17|2016-06-13|Volunteer: Moved|Volunteer: Moved||18.9||1|1|1|1|M|Hispanic||7|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|M|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504041803|504043821|3|0|1|503897667|1|0|1|500794453|7|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1950|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|90|Green||2016-12-02|2016-12-07|NaT||||3||1|1|1|1|F|Multi-race (Black & White)||7|No|Mother|28031|2|One Parent: Female|$30,000 to $34,999||||No||Self|General Site||Match Support|F|White||57|28205|High School Graduate|Single|Business: Mgt, Admin|28031|2|5|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504699174|504701602|36|0|2|504744195|1|0|2|500932604|10|1|500000295|2128173570|2|1||-1||-1|0|10|||18809|8|||1||8034889377453131101|4787903274998424796
M1951|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|686|Green||2015-04-15|2015-04-21|NaT||||22.5||1|1|1|1|F|Black||7|No|Mother|28213|1|One Parent: Female|$15,000 to $19,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||29|28211|Bachelors Degree|Single|Child/Day Care Worker||4|6|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503960671|503962680|31|0|2|504107327|1|0|2|500823484|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1||4013586283864837776|6084148439133243542
M1952|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|497|Green||2015-10-09|2015-10-27|NaT||||16.3||1|1|1|1|F|Hispanic||7|No|Mother|28212|1|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||18|28204|Some High School|Single|Student: College||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504447323|504449579|3|0|2|504303681|1|0|2|500846373|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1953|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|343|Green|Amachi|2016-03-15|2016-03-29|NaT||||11.3||1|1|2|2|M|Black||7|Yes|Mother|28208|K|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|Black||35|28273|Some College|Married|Business: Marketing|28203|1|1|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504405002|504403590|31|0|1|504241664|31|0|1|500884837|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|500000294|0|4309014537710246316
M1954|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|369|Green||2015-10-23|2015-10-30|2016-11-02|Volunteer: Time constraint|Volunteer: Time constraint||12.1||1|1|1|1|M|Black||7|Yes|Mother|28214|2|One Parent: Female|$35,000 to $39,999|||Y|Yes||School|General Community|Amachi|Enrollment|M|White||24|28203|Bachelors Degree|Single|Education|28203|0|2|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500018851|504182796|504184905|31|0|1|504378001|1|0|1|500851470|5|2|-2||4|1|500000294|-2|500000294|-2|0|4|||17159|12|||1||0|484306037765318169
M1955|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|228|Green||2015-10-16|2015-10-29|2016-06-13|Volunteer: Moved|Volunteer: Moved||7.5||1|1|1|1|F|Hispanic||7|No|Mother|28211|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||RTBM|F|White||18|28277|Some High School|Single|Student: College||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504112110|504114144|3|0|2|504409289|1|0|2|500848823|7|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1956|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2016-12-01|2017-01-30|NaT||||1.2||1|1|1|1|M|Black||7|No|Mother|28211|1|One Parent: Female|$30,000 to $34,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||25|28208|Bachelors Degree|Single|Business||1|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504682143|504684571|31|0|1|504313521|31|0|1|500932114|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1||967246839551912690|8408514790530965815
M1957|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|78|Green|Cabarrus County|2016-12-15|2016-12-19|NaT||||2.6||1|1|2|2|M|Black||7|No|Mother|28025|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||54|28025||Married|Clergy|28025|23|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504690665|504693093|31|0|1|502240986|31|0|1|500935855|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7671|13|||1|500016374|5208542183136337346|7044657180546140448
M1958|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|24|Green|Cabarrus County|2017-02-10|2017-02-11|NaT||||0.8||1|1|1|1|F|Multi-race (Hispanic & White)||7|No|Mother|28025|2|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|White||58|28025||Married|Business: Sales|28025|0|6|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504982340|504984889|35|0|2|504755956|1|0|2|500945687|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|500016374|3575183301237417432|0
M1959|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|76|Green||2016-12-01|2016-12-21|NaT||||2.5||1|1|1|1|M|Black||7|No|Mother|28208|1|One Parent: Female|$40,000 to $44,999||||Yes||School|General Community||Match Support|M|White||25|28203|Bachelors Degree|Single|Medical|85286|1|1|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504532089|504534422|31|0|1|504631918|1|0|1|500932298|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||976372749760822282|786532283575222488
M1960|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|118|Green|Cabarrus County|2016-11-02|2016-11-09|NaT||||3.9||1|1|1|1|F|Multi-race (Black & White)||7|No|GrandMother|28025|1|Grandparents|Unknown|Yes: Active|No||Yes||School|General Site|Cabarrus County|Match Support|F|White||17|28031|Some College|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504919506|504922026|36|0|2|504871597|1|0|2|500922780|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|1550830965009450729|0
M1961|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|300|Green||2015-11-19|2015-12-08|2016-10-03|Child: Changed school/site|Child: Changed school/site||9.9||1|1|3|3|F|Black||7|Yes|Mother|28212|1|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||18|28207|Some College|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504447304|504449560|31|0|2|504306107|1|0|2|500861429|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1962|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|344|Green||2014-11-09|2014-11-17|2015-10-27|Volunteer: Moved|Volunteer: Moved||11.3||2|2|1|1|M|Black||7|No|Mother|28211|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||20|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504101661|503631791|31|0|1|503925846|1|0|2|500793664|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1963|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|497|Green||2015-10-27|2015-10-27|NaT||||16.3||2|2|1|1|M|Black||7|No|Mother|28211|1|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||17|28209|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504101661|503631791|31|0|1|504302447|1|0|2|500852944|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1964|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|611|Green||2014-10-04|2014-10-06|2016-06-08|Volunteer: Moved|Volunteer: Moved||20.1||2|2|1|1|F|Black||7|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||19|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500011349|504049279|504051303|31|0|2|503898540|1|0|2|500780585|10|1|500000296|2128173564|4|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1965|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|F|Black||7|No|Mother|28212|K|One Parent: Female|Unknown|||Y|Yes||School|General Site||Match Support|F|White||16|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504049279|504051303|31|0|2|504741711|1|0|2|500928277|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1966|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|228|Green||2015-10-23|2015-10-29|2016-06-13|Volunteer: Moved|Volunteer: Moved||7.5||2|2|1|1|M|Hispanic||7|No|Father|28212|K|Two Parent|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||19|28277|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504478304|504178353|3|0|1|504443741|1|0|2|500851650|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1967|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|M|Hispanic||7|No|Father|28212|K|Two Parent|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504478304|504178353|3|0|1|504721191|1|0|2|500928490|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1968|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|495|Green||2015-10-29|2015-10-29|NaT||||16.3||1|1|1|1|F|Hispanic||7|Yes|Mother|28212|3|Two Parent|Less than $10,000||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28210|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504495891|504498176|3|0|2|504306089|1|0|2|500853677|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1969|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|355|Green||2016-03-09|2016-03-17|NaT||||11.7||1|1|1|1|F|Black||7|No|Mother|28208|1|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||27|28262|Masters Degree|Single|Medical: Admin|28210|0|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|503978167|503980164|31|0|2|504529749|31|0|2|500883846|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||2611337051335117774|0
M1970|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|184|Red||2015-03-11|2015-03-25|2015-09-25|Child/Family: Moved|Child/Family: Moved||6||1|1|1|1|F|Black||7|No|Mother|28206|K|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||30|28205|Bachelors Degree|Single|Arts, Entertainment, Sports|10011|2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500020752|504168599|504170705|31|0|2|504166556|1|0|2|500818071|10|2|-2||4|3||-2|500000294|-2|0|4|||46|2|||1||4863631750424600365|7044657180546140448
M1971|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|214|Green||2015-11-11|2015-11-11|2016-06-12|Volunteer: Moved|Volunteer: Moved||7||1|1|1|1|F|Black||7|No|Mother|28212|1|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|RTBM|F|Black||19|28203|Some High School||Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504505830|504508125|31|0|2|504419128|31|0|2|500858754|7|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1972|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|7|Green||2017-02-15|2017-02-28|NaT||||0.2||1|1|1|1|F|Multi-race (Black & Hispanic)||7|No|Mother|28212|1|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|Some Other Race||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|505026952|505029522|38|0|2|504725007|41|0|2|500946603|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1973|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|218|Green||2015-10-29|2015-10-29|2016-06-03|Volunteer: Moved|Volunteer: Moved||7.2||1|1|1|1|F|Hispanic||7|No|Mother|28212|1|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Site|VOL - HSBigs|RTBM|F|White||18|28226|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504495791|504444557|3|0|2|504452192|1|0|2|500853910|7|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M1974|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|687|Green|Cabarrus County|2015-04-13|2015-04-20|NaT||||22.6||1|1|1|1|F|Black||7|No|Mother|28083||One Parent: Female|$25,000 to $29,999|||Y|No||Self|General Community|Cabarrus County|Match Support|F|White||54|28081|Some College|Married|Finance: Banking|28026|13|5|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504075474|502762654|31|0|2|503792949|1|0|2|500822904|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374|0|4058276550489173605
M1975|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|311|Green|VOL - PreMatch, VOL - Mentoring Hispanic Youth, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-04-21|2016-04-30|NaT||||10.2||1|1|1|1|M|Hispanic||7|No|Mother|28205|K|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|Hispanic||37|28205|Bachelors Degree|Single|Tech: Engineer|28255|7|10|Community Engagement|Special Event|Big|General Community|VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504636958|504639369|3|0|1|504549037|3|0|1|500889969|10|2|-2||2|1||-2|500007920, 500011312, 500011315, 500011316|-2|0|4|||18809|8|||1|500007920, 500011312, 500011315, 500011316|4875067736105190023|0
M1976|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|148|Green||2016-09-16|2016-10-10|NaT||||4.9||1|1|1|1|M|Black||7|No|GrandMother|28212|K|One Parent: Female|$10,000 to $14,999|||Y|No||School|General Community||Match Support|M|White||25|28203|Bachelors Degree|Single|Finance: Accountant|28277|1|1|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504592686|504595050|31|0|1|504594988|1|0|1|500908171|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||0|0
M1977|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|90|Green||2016-12-02|2016-12-07|NaT||||3||1|1|1|1|F|Black||7|No|Mother|28031|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||45|28031|Bachelors Degree|Divorced|Business: Human Resources|28031|2|11|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504951117|504953668|31|0|2|504671040|1|0|2|500932594|10|1|500000295|2128173570|2|1||-1||-1|0|4|||18809|8|||1||8034889377453131101|0
M1978|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|36|Green||2017-01-23|2017-01-30|NaT||||1.2||1|1|1|1|M|Black||7|No|Mother|28214||One Parent: Female|$20,000 to $24,999||||Yes||Relative|General Community||Match Support|M|Black||40|28269|Bachelors Degree|Married|Consultant|28277|11|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504188050|504190159|31|0|1|504845940|31|0|1|500941540|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|3|||46|2|||1||9080589164524051479|458259588635328527
M1979|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|15|Green||2017-02-20|2017-02-20|NaT||||0.5||1|1|1|1|M|Hispanic||7|No|Mother|28212|1|Two Parent|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||16|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504998019|505000579|3|0|1|504739301|1|0|2|500947203|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1980|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|24|Green||2017-01-17|2017-02-06|2017-03-02|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||0.8||1|1|1|1|F|Black||7|No|Mother|28208|1|One Parent: Female|$25,000 to $29,999||||No||Self|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|F|White||27|28203|Masters Degree|Single|Education: Teacher|28216|2|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504915468|504917988|31|0|2|504349057|1|0|2|500940444|5|2|-2||4|1|500007920, 500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1||0|6156547733130613405
M1981|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|502|Green||2015-10-16|2015-10-22|NaT||||16.5||1|1|1|1|F|Native Hawaiian or Other Pacific Islander||7|No|Mother|28213|1|Two Parent|$30,000 to $34,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504461758|504464016|5|0|2|504468576|1|0|2|500848828|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1982|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|210|Green||2015-11-11|2015-11-11|2016-06-08|Volunteer: Moved|Volunteer: Moved||6.9||2|2|1|1|M|Black||7|No|Mother|28212|K|Two Parent|Less than $10,000|||Y|Yes||School|General Site|VOL - HSBigs|Match Support|M|Black||19|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504496553|504498838|31|0|1|504419043|31|0|1|500858609|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1983|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|M|Black||7|No|Mother|28212|K|Two Parent|Less than $10,000|||Y|Yes||School|General Site|VOL - HSBigs|Match Support|M|Multi-race (Asian & White)||16|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504496553|504498838|31|0|1|504723806|37|0|1|500929222|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1984|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|372|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-02-19|2016-02-29|NaT||||12.2||1|1|1|1|F|Black||7|No|Mother|28211|K|One Parent: Female|$25,000 to $29,999|Yes: Active|No|Y|Yes||Self|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Business|28270|10|8|AA Task Force|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504345301|504347523|31|0|2|504373845|1|0|2|500880266|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||6247|12|||1|500007920, 500011315, 500011316|421482027904269589|1981915209225039472
M1985|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|14|Green||2017-02-09|2017-02-21|NaT||||0.5||1|1|1|1|F|Black||7|No|GrandMother|28208|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Amachi|Match Support|F|White||36|28202|Bachelors Degree|Married|Business: Mgt, Admin|28204|1|8|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504622170|504624581|31|0|2|504802975|1|0|2|500945483|10|2|-2||2|1|500000294|-2||-2|0|4|||17159|12|||1||8568001799025358453|0
M1986|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|2|2|M|Black||7|Yes|Mother|28212|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|F|White||17|28210|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504495730|504044051|31|0|1|504428689|1|0|2|500929211|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1987|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|316|Green||2015-11-02|2015-11-18|2016-09-29|Child: Changed school/site|Child: Changed school/site||10.4||2|2|2|2|M|Black||7|Yes|Mother|28212|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|F|White||17|28210|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500022905|504495730|504044051|31|0|1|504428689|1|0|2|500855269|10|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1988|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|228|Green||2015-10-23|2015-10-29|2016-06-13|Volunteer: Moved|Volunteer: Moved||7.5||2|2|1|1|F|Black||7|No|Mother|28212|1|Two Parent|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||19|28226|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504478319|504480593|31|0|2|504419161|1|0|2|500851614|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1989|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|F|Black||7|No|Mother|28212|1|Two Parent|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504478319|504480593|31|0|2|504723859|1|0|2|500928462|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M1990|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|35|Green||2017-01-20|2017-01-31|NaT||||1.1||1|1|2|2|M|Hispanic||7|No|Mother|28212|1|Two Parent|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||17|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504997997|505000557|3|0|1|504729038|1|0|2|500941217|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1991|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|12|Green||2017-02-06|2017-02-23|NaT||||0.4||1|1|1|1|F|Black||7|Yes|Mother|28208|K|One Parent: Female|$15,000 to $19,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||30|28209|Bachelors Degree|Single|Medical|27410|6|10|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500008321|504617761|504620172|31|0|2|504911953|1|0|2|500944724|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|5|||7464|9|||1||0|7683788406654221511
M1992|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|66|Green||2015-11-02|2015-11-03|2016-01-08|Child/Family: Moved|Child/Family: Moved||2.2||1|1|2|2|M|Black||7|No|Mother|28212|K|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Black||18|28104|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504478033|504480307|31|0|1|504442352|31|0|2|500855268|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1993|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|33|Green||2017-01-25|2017-02-02|NaT||||1.1||1|1|1|1|M|Black||7|No|Mother|28031|1|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|M|Multi-race (Black & Hispanic)||20|28035||Single|Student: College||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504956464|504959015|31|0|1|504901170|38|0|1|500941974|10|1|500000295|2128173570|2|1||-1||-1|0|4|||7464|9|||1||8034889377453131101|0
M1994|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|156|Green||2016-01-08|2016-01-08|2016-06-12|Volunteer: Moved|Volunteer: Moved||5.1||2|2|2|2|F|Black||7|No|Mother|28212|K|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|Black||18|28104|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504571845|504574179|31|0|2|504442352|31|0|2|500870842|10|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1995|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|91|Green||2016-12-06|2016-12-06|NaT||||3||2|2|1|1|F|Black||7|No|Mother|28212|K|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||17|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022908|504571845|504574179|31|0|2|504731823|1|0|2|500933545|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1996|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|50|Green||2017-01-09|2017-01-16|NaT||||1.6||1|1|1|1|F|Black||7|No|Mother|28208|1|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||27|28210|Bachelors Degree|Single|Education|28203|0|0|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504970056|504972603|31|0|2|504764294|1|0|2|500939113|10|1|500000295|2128207319|2|1||-1||-1|0|4|||46|2|||1||3935539763241716148|0
M1997|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|214|Green||2015-11-11|2015-11-11|2016-06-12|Volunteer: Moved|Volunteer: Moved||7||2|2|1|1|F|Hispanic||7|Yes|Mother|28212|K|Two Parent|$20,000 to $24,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504505823|504508118|3|0|2|504416646|1|0|2|500858665|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1998|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|F|Hispanic||7|Yes|Mother|28212|K|Two Parent|$20,000 to $24,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022908|504505823|504508118|3|0|2|504741636|1|0|2|500929207|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M1999|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|203|Green||2015-11-23|2015-11-23|2016-06-13|Volunteer: Moved|Volunteer: Moved||6.7||2|2|1|1|F|Hispanic||7|No|Mother|28212|K|Two Parent|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||18|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504525282|504527614|3|0|2|504452202|1|0|2|500862563|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2000|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|F|Hispanic||7|No|Mother|28212|K|Two Parent|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||16|28104|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504525282|504527614|3|0|2|504732675|1|0|2|500929171|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2001|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|323|Green||2015-11-11|2015-11-11|2016-09-29|Child: Changed school/site|Child: Changed school/site||10.6||1|1|2|2|M|Hispanic||7|Yes|Mother|28203|K|Grandparents|$10,000 to $14,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|White||18|28226|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504502423|504504712|3|0|1|504452221|1|0|2|500858853|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2002|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|227|Green||2015-10-23|2015-10-29|2016-06-12|Volunteer: Moved|Volunteer: Moved||7.5||2|2|1|1|F|Hispanic||7|No|Mother|28211|K|Two Parent|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||19|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504461688|504463946|3|0|2|504442316|1|0|2|500851491|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2003|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|F|Hispanic||7|No|Mother|28211|K|Two Parent|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504461688|504463946|3|0|2|504723876|1|0|2|500928459|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2004|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|35|Green||2017-01-17|2017-01-31|NaT||||1.1||1|1|1|1|F|Hispanic||7|No|Mother|28212|1|Two Parent|$15,000 to $19,999||||Yes||School|General Site||Match Support|F|White||16|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504998028|505000588|3|0|2|504731856|1|0|2|500940358|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2005|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|336|Green||2016-03-01|2016-04-05|NaT||||11||1|1|1|1|M|Black||7|No|Mother|28273|K|One Parent: Female|$45,000 to $49,999|||Y|Yes||School|General Community||Match Support|M|White||25|28210|Bachelors Degree|Single|Finance|28211|10|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504276350|504278550|31|0|1|504273397|1|0|1|500882201|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||6202343250032725030|1176389127668227778
M2006|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|42|Green||2016-12-08|2017-01-24|NaT||||1.4||1|1|1|1|F|Black||7|No|Mother|28208|1|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site||Match Support|F|White||27|28209|Bachelors Degree|Single|Business: Sales|28203|2|6|Current/Previous Big|Other Big|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504960292|504962843|31|0|2|504714143|1|0|2|500934310|10|1|500000295|2128207319|2|1||-1||-1|0|4|||17159|12|||1||3935539763241716148|0
M2007|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|366|Green||2015-05-19|2015-05-19|2016-05-19|Volunteer: Time constraint|Volunteer: Time constraint||12||1|1|1|1|M|Black||7|No|Mother|28212||One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community|Amachi|Enrollment|M|White||46|28031|High School Graduate|Married|Business: Sales|28219|1|0|Relative|Relative|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500018851|504211341|504207614|31|0|1|504224356|1|0|1|500827550|5|2|-2||4|1|500000294|-2|500000294|-2|0|4|||17161|11|||1||392688197545050058|7500593753197857009
M2008|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|90|Green||2016-12-02|2016-12-07|NaT||||3||1|1|1|1|M|White||7|No|Father|28031|1|One Parent: Male|$30,000 to $34,999||||No||School|General Site||Match Support|F|Black||43|28083|PHD|Married|Business|28031|1|6|Community Engagement|Special Event|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504960210|504962761|1|0|1|504666420|31|0|2|500932599|10|1|500000295|2128173570|2|1||-1||-1|0|4|||18809|8|||1||8034889377453131101|0
M2009|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|402|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-01-20|2016-01-30|NaT||||13.2||1|1|1|1|F|Black||7|No|Mother|28075|K|Two Parent|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||36|28036|Bachelors Degree|Married|Self-Employed, Entrepreneur|28036|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504453477|504455735|31|0|2|503803589|1|0|2|500873679|10|2|-2||2|1||-2||-2|0|5|||7464|9|||1|500007920, 500011315, 500011316|6627885846854295604|2141487034287122220
M2010|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|227|Green||2015-10-23|2015-10-29|2016-06-12|Volunteer: Moved|Volunteer: Moved||7.5||1|1|1|1|M|White||7|No|Mother|28212|K|One Parent: Female|$20,000 to $24,999||||Yes||School|General Site|VOL - HSBigs|RTBM|M|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504478083|504480357|1|0|1|504438031|1|0|1|500851581|7|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2011|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|210|Green||2015-11-11|2015-11-11|2016-06-08|Volunteer: Moved|Volunteer: Moved||6.9||2|2|1|1|M|Black||7|No|Father|28212|K|Two Parent|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Black||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504505846|504508141|31|0|1|504438050|31|0|2|500858673|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2012|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|M|Black||7|No|Father|28212|K|Two Parent|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504505846|504508141|31|0|1|504723759|1|0|2|500929196|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2013|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|119|Green|Cabarrus County|2016-10-31|2016-11-08|NaT||||3.9||1|1|1|1|F|Hispanic||7|No|Mother|28027|1|One Parent: Female|Unknown||||Yes||School|General Site|Cabarrus County|Match Support|F|Hispanic||17|28217|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504918273|504920793|3|0|2|504871256|3|0|2|500921842|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||0|4|||1|500016374|1550830965009450729|0
M2014|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|292|Green||2016-05-03|2016-05-19|NaT||||9.6||1|1|1|1|F|Black||7|No|Mother|28212||One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|Black||25|28277|Bachelors Degree|Single|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504260164|504262304|31|0|2|504523141|31|0|2|500891594|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||0|4802885652788112046
M2015|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|88|Green||2016-12-06|2016-12-09|NaT||||2.9||1|1|1|1|F|Asian||7|No|Father|28211|1|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||17|28270|Some College||Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504963048|504965599|4|0|2|504724989|1|0|2|500933550|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|2837068013653064810
M2016|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|476|Green|Cabarrus County|2015-10-30|2015-11-17|NaT||||15.6||1|1|2|2|F|Black||7|No|Mother|28083||One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|F|Black||30|28027|Masters Degree|Married|Unemployed|28027|2|5|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504241295|504243414|31|0|2|503542037|31|0|2|500854635|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|34|2|||7464|9|||1|500016374|0|1579263579908564057
M2017|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|88|Green||2016-12-07|2016-12-09|NaT||||2.9||1|1|1|1|M|White||7|No|Mother|28211|1|One Parent: Female|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|Black||17|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504965733|504968284|1|0|1|504739346|31|0|2|500933977|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2018|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|222|Green||2015-11-02|2015-11-03|2016-06-12|Volunteer: Moved|Volunteer: Moved||7.3||2|2|1|1|M|Hispanic||7|No|Mother|28212|K|Two Parent|$10,000 to $14,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|Multi-race (Hispanic & White)||19|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500011349|504496656|504498942|3|0|1|504419085|35|0|2|500855270|10|1|500000296|2128173564|4|1|500014068|-1||-1|0|3|||0|4|||1||2762897743412756173|0
M2019|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|M|Hispanic||7|No|Mother|28212|K|Two Parent|$10,000 to $14,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|White||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504496656|504498942|3|0|1|504723816|1|0|1|500929217|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|3|||0|4|||1||2762897743412756173|0
M2020|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|214|Green||2015-11-11|2015-11-11|2016-06-12|Volunteer: Moved|Volunteer: Moved||7||2|2|1|1|F|Black||7|No|Mother|28212|K|Two Parent|$10,000 to $14,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|Black||19|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504502456|504504745|31|0|2|504428583|31|0|2|500858790|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2021|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|F|Black||7|No|Mother|28212|K|Two Parent|$10,000 to $14,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|Black||17|28203|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504502456|504504745|31|0|2|504739362|31|0|2|500929186|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|3|||0|4|||1||2762897743412756173|0
M2022|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|227|Green||2015-10-23|2015-10-29|2016-06-12|Volunteer: Moved|Volunteer: Moved||7.5||2|2|1|1|M|Hispanic||7|No|Mother|28211|K|Two Parent|$30,000 to $34,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|Some Other Race||19|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504478022|504480296|3|0|1|504428560|41|0|1|500851592|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2023|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|2|2|M|Hispanic||7|No|Mother|28211|K|Two Parent|$30,000 to $34,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|White||18|28226|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022908|504478022|504480296|3|0|1|504452221|1|0|2|500929203|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2024|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|190|Green||2015-12-03|2015-12-17|2016-06-24|Volunteer: Time constraint|Volunteer: Time constraint||6.2||1|1|1|1|M|White||6|Yes|GrandMother|28083|K|Grandparents|$20,000 to $24,999||||Yes||School|General Site|Cabarrus County|RTBM|F|Some Other Race||48|28083|Bachelors Degree|Married|Medical|27103|0|1|BBBS National Site|Web Link|Big|General Site|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|504530664|504532996|1|0|1|504363589|41|0|2|500864986|7|1|500000295|2128232374|4|1|500016374|-1|500016374|-1|0|4|||46|2|||1||2043334928777030191|0
M2025|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|32|Green||2015-10-23|2015-10-29|2015-11-30|Child/Family: Moved|Child/Family: Moved||1.1||1|1|2|2|M|Multi-race (Black & Hispanic)||6|No|Mother|28212|K|One Parent: Female|$10,000 to $14,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|White||19|28211|Some High School||Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500020909|504461329|504463587|38|0|1|504442387|1|0|1|500851488|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2026|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|481|Green|Cabarrus County|2015-11-10|2015-11-12|NaT||||15.8||1|1|1|1|M|Black||6|No|Mother|28081|K|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28025|Bachelors Degree|Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504366634|502790820|31|0|1|504346767|1|0|1|500858202|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||17159|12|||1|500016374|0|7044657180546140448
M2027|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|28|Green||2017-02-07|2017-02-07|NaT||||0.9||1|1|1|1|M|Hispanic||6|No|Mother|28211||One Parent: Female|Unknown||||Yes||School|General Site||Match Support|M|Some Other Race||17|28173|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|505004269|505006829|3|0|1|504729049|41|0|1|500945017|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2028|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|228|Green||2015-10-23|2015-10-29|2016-06-13|Volunteer: Moved|Volunteer: Moved||7.5||1|1|1|1|M|Black||6|Yes|Mother|28212|K|One Parent: Female|Less than $10,000||||Yes||Relative|General Site|VOL - HSBigs|RTBM|M|Black||19|28206|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504461792|504031285|31|0|1|504418898|31|0|1|500851564|7|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2029|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|35|Green||2017-01-18|2017-01-31|NaT||||1.1||1|1|1|1|F|Hispanic||6|No|Mother|28211|1|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|White||16|28270|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504997973|505000533|3|0|2|504729023|1|0|2|500940765|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2030|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|394|Red|Cabarrus County|2015-10-21|2015-10-21|2016-11-18|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||12.9||1|1|4|4|F|Black||6|No|GrandMother|28083|K|One Parent: Female|$30,000 to $34,999||||Yes||School|General Community|Cabarrus County|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500022817|504439153|503587420|31|0|2|500189709|31|0|2|500850116|10|2|500016307||4|3|500016374|-2|500000294, 500016374|-2|0|4|||2230|7|||1|500016374|6810228174639243761|0
M2031|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|54|Green||2017-01-03|2017-01-12|NaT||||1.8||1|1|1|1|F|Black||6|No|Mother|28208|1|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Site||Match Support|F|White||53|28226||Widowed|Homemaker||0|0|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504960282|504962833|31|0|2|504833597|1|0|2|500937903|10|1|500000295|2128207319|2|1||-1||-1|0|4|||46|2|||1||3935539763241716148|0
M2032|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|463|Green||2015-11-17|2015-11-30|NaT||||15.2||1|1|2|2|F|Multi-race (Black & White)||6|No|Mother|28269|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Amachi|Match Support|F|Black||46|28216|Bachelors Degree|Single|Business: Marketing|28036|0|3|Self|Self|Big|General Community|VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|504360025|504222143|36|0|2|503844843|31|0|2|500860778|10|2|-2||2|1|500000294|-2|500007920, 500011312, 500011315, 500011316|-2|0|4|||7464|9|||1||0|7044657180546140448
M2033|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|191|Green||2015-11-30|2015-11-30|2016-06-08|Volunteer: Moved|Volunteer: Moved||6.3||2|2|2|2|M|Black||6|No|Mother|28212|K|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|M|White||19|28211|Some High School||Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504524429|504526760|31|0|1|504442387|1|0|1|500863715|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2034|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|64|Green||2016-11-17|2016-11-17|2017-01-20|Child: Changed school/site|Child: Changed school/site||2.1||2|2|2|2|M|Black||6|No|Mother|28212|K|One Parent: Female|$15,000 to $19,999||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504524429|504526760|31|0|1|504729038|1|0|2|500929220|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2035|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|227|Green||2015-10-23|2015-10-29|2016-06-12|Volunteer: Moved|Volunteer: Moved||7.5||2|2|1|1|F|Hispanic||6|No|Mother|28212|K|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||19|28209|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504441583|504443839|3|0|2|504441249|1|0|2|500851492|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2036|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|F|Hispanic||6|No|Mother|28212|K|One Parent: Female|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28202|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504441583|504443839|3|0|2|504739276|1|0|2|500929181|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2037|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|227|Green||2015-10-23|2015-10-29|2016-06-12|Volunteer: Moved|Volunteer: Moved||7.5||2|2|1|1|M|Multi-race (Black & White)||6|No|Mother|28212|K|One Parent: Female|Less than $10,000||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|Black||18|28213|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504461293|504463551|36|0|1|504452241|31|0|1|500851487|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2038|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|M|Multi-race (Black & White)||6|No|Mother|28212|K|One Parent: Female|Less than $10,000||||Yes||Relative|General Site|VOL - HSBigs|Match Support|M|White||17|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022908|504461293|504463551|36|0|1|504721236|1|0|1|500928486|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|3|||0|4|||1||2762897743412756173|0
M2039|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|208|Green||2015-11-11|2015-11-18|2016-06-13|Volunteer: Moved|Volunteer: Moved||6.8||2|2|1|1|F|Hispanic||6|No|Mother|28212|K|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|White||18|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504502404|504504693|3|0|2|504418950|1|0|2|500858866|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2040|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|F|Hispanic||6|No|Mother|28212|K|One Parent: Female|$30,000 to $34,999||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|White||18|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504502404|504504693|3|0|2|504732709|1|0|2|500929215|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2041|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|202|Green||2015-11-23|2015-11-23|2016-06-12|Volunteer: Moved|Volunteer: Moved||6.6||2|2|1|1|M|Hispanic||6|No|Mother|28212|K|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||19|28277|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504530464|504532796|3|0|1|504428766|1|0|2|500862566|10|1|500000296|2128173564|4|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2042|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|110|Green||2016-11-17|2016-11-17|NaT||||3.6||2|2|1|1|M|Hispanic||6|No|Mother|28212|K|Two Parent|Unknown||||Yes||School|General Site||Match Support|F|White||16|28203|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504530464|504532796|3|0|1|504739376|1|0|2|500929190|10|1|500000296|2128173564|2|1||-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2043|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|206|Green||2015-11-19|2015-11-19|2016-06-12|Volunteer: Moved|Volunteer: Moved||6.8||2|2|1|1|F|Hispanic||6|No|Mother|28212|K|Two Parent|Less than $10,000|||Y|Yes||School|General Site|VOL - HSBigs|Match Support|F|White||19|28226|High School Graduate|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504524449|504526780|3|0|2|504442325|1|0|2|500861407|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2044|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|89|Green|VOL - HSBigs|2016-12-07|2016-12-08|NaT||||2.9||2|2|1|1|F|Hispanic||6|No|Mother|28212|K|Two Parent|Less than $10,000|||Y|Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28277|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500022909|504524449|504526780|3|0|2|504934167|1|0|2|500933981|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||7464|9|||1|500014068|2762897743412756173|0
M2045|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|397|Green|Cabarrus County|2016-01-25|2016-02-04|NaT||||13||1|1|1|1|F|Multi-race (Black & White)||6|No|Mother|28025|K|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Cabarrus County|Match Support|F|White||36|28025|Some College|Divorced|Finance: Banking|28262|0|5|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504533461|504535058|36|0|2|504565015|1|0|2|500875147|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||17159|12|||1|500016374|9080589164524051479|2141487034287122220
M2046|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|88|Green||2016-12-07|2016-12-09|NaT||||2.9||1|1|1|1|M|White||6|No|Mother|28212|1|Two Parent|$30,000 to $34,999||||Yes||School|General Site||Match Support|F|White||17|28277|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504965745|504968296|1|0|1|504721170|1|0|2|500933971|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2047|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|35|Green||2017-01-18|2017-01-31|NaT||||1.1||1|1|1|1|M|Hispanic||6|No|Mother|28211|1|Two Parent|$10,000 to $14,999||||Yes||School|General Site||Match Support|F|Black||17|28214|Some High School||Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500016270|504997959|505000519|3|0|1|504741689|31|0|2|500940763|10|1|500000296|2128173564|2|1||-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2048|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|39|Green||2017-01-10|2017-01-27|NaT||||1.3||1|1|1|1|M|Black||6|No|Mother|28227|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Black||29|28262|Masters Degree|Single|Education: Teacher||0|3|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020753|504415884|504418136|31|0|1|504930194|31|0|1|500939321|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7462|13|||1||5388127382485844452|1653590244760837916
M2049|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|194|Green||2015-11-19|2015-12-01|2016-06-12|Volunteer: Moved|Volunteer: Moved||6.4||1|1|1|1|M|Black||6|Yes|Mother|28215|K|One Parent: Female|$10,000 to $14,999||||Yes||School|General Site|VOL - HSBigs|RTBM|F|White||18|28210|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504524390|504445917|31|0|1|504438266|1|0|2|500861424|7|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2050|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|479|Green|Cabarrus County|2015-11-06|2015-11-14|NaT||||15.7||1|1|3|3|M|Black||6|No|Mother|28075|K|One Parent: Female|$60,000 to $74,999||||Yes||School|General Community|Cabarrus County|Match Support|M|Black||52|28025||Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504442355|504444611|31|0|1|500790181|31|0|1|500857210|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||7464|9|||1|500016374|3380316005507597709|2602987289799151214
M2051|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|RTBM|210|Green||2015-11-11|2015-11-11|2016-06-08|Volunteer: Moved|Volunteer: Moved||6.9||1|1|1|1|F|White||6|No|Mother|28212|K|Two Parent|$45,000 to $49,999||||No||School|General Site|VOL - HSBigs|RTBM|F|Multi-race (Black & White)||18|28105|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504502465|504504754|1|0|2|504438196|36|0|2|500858657|7|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2052|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|135|Green|Cabarrus County|2016-10-11|2016-10-23|NaT||||4.4||1|1|1|1|F|White||6|No|GrandMother|28025|1|Grandparents|$15,000 to $19,999||||Yes||Self|General Community|Cabarrus County|Match Support|F|White||46|28081|Associate Degree|Married|Law: Paralegal|28207|2|6|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504819441|504821927|1|0|2|504805076|1|0|2|500914392|10|2|500016307||2|1|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||17159|12|||1|500016374|5064856656261650513|0
M2053|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|482|Green||2015-11-11|2015-11-11|NaT||||15.8||1|1|1|1|F|Hispanic||6|No|Mother|28212|1|One Parent: Female|Unknown||||Yes||Relative|General Site|VOL - HSBigs|Match Support|F|White||18|28226|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|0|1|277|60|598|500000170|500022909|504502442|504504731|3|0|2|504428719|1|0|2|500858805|10|1|500000296|2128173564|2|1|500014068|-1|500014068|-1|0|3|||0|4|||1||2762897743412756173|0
M2054|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|119|Green|Cabarrus County|2016-11-02|2016-11-08|NaT||||3.9||1|1|1|1|F|Multi-race (Black & White)||6|No|Mother|28025|1|One Parent: Female|Less than $10,000||||Yes||School|General Site|Cabarrus County|Match Support|F|White||17|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504918305|504920825|36|0|2|504875774|1|0|2|500922787|10|1|500000296|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|5208542183136337346|0
M2055|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|209|Green||2016-07-29|2016-08-10|NaT||||6.9||1|1|1|1|M|White||6|No|Mother|28205|K|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||33|28205|Masters Degree|Single|Business|28203|3|0|Other|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504620049|504207619|1|0|1|504659863|1|0|1|500901159|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7671|13|||1||8998367770661215127|610388910998118020
M2056|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|88|Green||2016-12-06|2016-12-09|NaT||||2.9||1|1|1|1|M|Hispanic||6|No|Mother|28207|K|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site||Match Support|M|Some Other Race||26|28078|Bachelors Degree|Single|Consultant|28281|2|11|BBBS National Site|Web Link|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504899050|504901570|3|0|1|504850064|41|0|1|500933350|10|1|500000295|2128207319|2|1||-1||-1|0|4|||46|2|||1||3935539763241716148|0
M2057|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|63|Green||2016-12-12|2017-01-03|NaT||||2.1||1|1|1|1|F|Black||5|No|Mother|28217|K|One Parent: Female|Less than $10,000||||Yes||School|General Site||Match Support|F|White||31|28205|Masters Degree|Living w/ Significant Other|Tech: Management|28281|1|0|Wells Fargo|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500015820|504951130|504953681|31|0|2|504806060|1|0|2|500934868|10|1|500000295|2128207319|2|1||-1||-1|0|4|||18266|3|||1||3935539763241716148|0
M2058|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|92|Green|Cabarrus County|2016-12-05|2016-12-05|NaT||||3||1|1|1|1|M|Black||5|No|Mother|28027|K|Two Parent|Less than $10,000||||Yes||School|General Site|Cabarrus County|Match Support|M|White||18|28025|Some High School|Single|Student: High School||0|0|Self|Self|Big|General Site|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500012459|504918090|504920610|31|0|1|504883844|1|0|1|500933119|10|1|500000295|2128173571|2|1|500016374|-1|500016374|-1|0|4|||7464|9|||1|500016374|6810228174639243761|0
M2059|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|223|Green||2015-10-23|2015-10-29|2016-06-08|Volunteer: Moved|Volunteer: Moved||7.3||2|2|1|1|F|Hispanic||2|No|Mother|28212|K|Two Parent|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|Hispanic||18|28273|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site|VOL - HSBigs|Match Support|0|1|1|0|277|60|598|500000170|500011349|504461307|504463565|3|0|2|504452261|3|0|2|500851489|10|1|500000296|2128173564|4|1|500014068|-1|500014068|-1|0|4|||0|4|||1||2762897743412756173|0
M2060|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|111|Green||2016-11-16|2016-11-16|NaT||||3.6||2|2|1|1|F|Hispanic||2|No|Mother|28212|K|Two Parent|Unknown||||Yes||School|General Site|VOL - HSBigs|Match Support|F|White||17|28211|Some High School|Single|Student: High School||0|0||High School Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500016270|504461307|504463565|3|0|2|504725042|1|0|2|500928282|10|1|500000296|2128173564|2|1|500014068|-1||-1|0|4|||0|4|||1||2762897743412756173|0
M2061|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1532|Red||2012-06-07|2012-06-19|2016-08-29|Child: Graduated|Child: Graduated||50.3||1|1|2|2|M|Hispanic|Mexican|18|No|Mother|28215|7|One Parent: Female|Less than $10,000|||Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502527168|502527621|3|10|1|501646021|3|0|1|500618440|10|2|-2||4|3|500005291|-2||-2|2203|12|||7464|9|||1||0|0
M2062|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1225|Green||2013-10-24|2013-10-29|NaT||||40.2||2|2|1|1|M|Hispanic|Mexican|16|No|Mother|28213|9|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Hispanic||29|28214|Bachelors Degree|Single|Self-Employed, Entrepreneur|28214|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|502374716|502375154|3|10|1|503560077|3|0|1|500723012|10|2|-2||2|1||-2||-2|0|4|||46|2|||1||0|0
M2063|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|510|Red|VOL - Mentoring Hispanic Youth|2013-12-12|2013-12-20|2015-05-14|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||16.8||1|1|1|1|F|Hispanic|Mexican|16|No|Mother|28208|6|Two Parent|Unknown|||Y|Yes|Spanish Radio|Media|General Community||Match Support|F|White||35|28214|Bachelors Degree|Single|Transport: Flight Attendant|85034|0|3|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500017777|503490571|503492439|3|10|2|503645850|1|0|2|500738556|10|2|-2||4|3||-2|500000294|-2|7068|1|||7464|9|||1|500011312|9076057728106637014|0
M2064|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1240|Green||2012-03-30|2012-05-24|2015-10-16|Volunteer: Moved|Volunteer: Moved||40.7||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28205|4|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||28|27235|Bachelors Degree||Business: Engineer||1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502874566|502875969|3|10|2|502894480|1|0|2|500607372|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1||9080589164524051479|0
M2065|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|868|Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2014-10-15|2014-10-21|NaT||||28.5||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28212|5|Two Parent|Unknown|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||30|28226||Single|Unemployed||0|0|Relative|Relative|Big|General Community|PERL 2014-2016|Match Support|1|0|0|1|277|60|598|500000170|500020753|503895506|503897502|3|10|2|504026849|3|0|2|500784082|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17161|11|||1|500011312, 500014681|2056258660718146620|0
M2066|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1042|Green|VOL - Mentoring Hispanic Youth|2014-04-28|2014-04-30|NaT||||34.2||1|1|1|1|F|Hispanic|Mexican|13|No|Mother|28205|5|One Parent: Female|Unknown|||Y|Yes|BBBS National Site|Web Link|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||44|28213|Bachelors Degree|Married|Medical|28216|2|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|503706992|503708958|3|10|2|503709061|1|0|2|500761338|10|2|-2||2|1|500011312|-2||-2|34|2|||7464|9|||1|500011312|0|7044657180546140448
M2067|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|568|Green||2013-10-17|2014-02-17|2015-09-08|Child/Family: Moved|Child/Family: Moved||18.7||1|1|5|5|F|Hispanic|Mexican|12|No|Mother|28025||Other/Unknown|Unknown||||Yes||School|General Site||Match Support|F|White||44|28075|Bachelors Degree|Married|Tech: Computer/Programmer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|1|0|1|0|277|60|598|500000170|500012459|503673635|503675596|3|10|2|502143796|1|0|2|500720476|10|1|500000295|2128212924|4|1||-1|500007920, 500011315, 500011316, 500016374|-1|0|4|||7496|10|||1||3232906304025417619|0
M2068|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Completed|Match Support|862|Green|VOL - Mentoring Hispanic Youth|2014-02-03|2014-02-19|2016-06-30|Child: Graduated|Child: Graduated||28.3||1|1|1|1|F|Hispanic|Mexican|12|No|Mother|28217|5|One Parent: Female|Unknown||||Yes||School|General Site||Match Support|F|White||28|28277|Bachelors Degree|Single|Medical: Nurse|28203|1|6|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500013781|503779460|503781437|3|10|2|503659745|1|0|2|500746618|10|1|500000295|2128173557|4|1||-1||-1|0|4|||7464|9|||1|500011312|8981704271528751143|0
M2069|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|S|Active|Match Support|882|Green|mentor2.0, mentor2.0 2014|2014-10-07|2014-10-07|NaT||||29||1|1|1|1|M|Black|Other African|18|No|Father|28212|9|One Parent: Male|Unknown|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2014|Match Support|M|White||38|28277|Juris Doctorate (JD)|Married|Law: Lawyer|28202|8|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504050606|504052630|31|31|1|503972019|1|0|1|500781247|10|1|500014504||2|1|500014505, 500014506|-1|500014506|-1|0|4|||7462|13|||1|500014505, 500014506|702163000107564368|0
M2070|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2412|Green||2010-07-07|2010-07-30|NaT||||79.2||1|1|1|1|M|Black|Other African|17|No|Mother|28269|11|One Parent: Female|Unknown|||Y|Yes||Relative|General Community||Match Support|M|White||35|28205|Masters Degree|Married|Tech: Engineer|28115|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501872144|501872517|31|31|1|502063676|1|0|1|500460156|10|2|-2||2|1||-2||-2|0|3|||46|2|||1||253338316288302752|8242487816501170810
M2071|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1995|Green|2010-2012 OJJDP JJI|2011-09-06|2011-09-20|NaT||||65.5||1|1|1|1|M|Black|Other African|15|No|Mother|29732|10|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|29720|Bachelors Degree|Married|Business: Sales|28134|4|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502455004|502074089|31|31|1|502680045|1|0|1|500553363|10|2|-2||2|1|500005291|-2||-2|0|4|||7464|9|||1|500005291|0|0
M2072|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|622|Red|VOL - Mentoring Hispanic Youth|2014-11-15|2014-12-16|2016-08-29|Child: Family structure changed|Child: Family structure changed||20.4||1|1|1|1|M|Hispanic|Other Central American|13|No|Mother|28214|6|One Parent: Female|Unknown|||Y|Yes||Therapist/Counselor|General Community|VOL - Mentoring Hispanic Youth|Match Support|M|Hispanic||37|28078|Associate Degree|Single|Finance|28217|0|3|Coworker|Workplace Partner|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|1|0|1|0|277|60|598|500000170|500017777|504059280|504061304|3|14|1|503998203|3|0|1|500796014|10|2|-2||4|3|500011312|-2|500011312|-2|0|5|||7447|3|||1|500011312|5604470640552265812|0
M2073|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|375|Yellow|VOL - Mentoring Hispanic Youth|2014-09-19|2014-09-29|2015-10-09|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||12.3||2|2|2|2|F|Hispanic|Other Central American|10|No|Mother|28217|1|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|RTBM|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500017777|503355390|503348836|3|14|2|503843020|3|0|2|500777040|7|2|-2||4|2|500011312, 500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|500011312|0|0
M2074|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1232|Green||2013-10-08|2013-10-22|NaT||||40.5||1|1|1|1|F|Hispanic|Other Central American|9|No|Mother|28262|3|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||30|28214|Bachelors Degree|Single|Law: Paralegal|28214|2|5|Self|Self|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|503467766|502751081|3|14|2|503543048|1|0|2|500717156|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1||4356567821563751981|0
M2075|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3253|Green||2007-07-10|2007-07-20|2016-06-15|Child: Graduated|Child: Graduated||106.9||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28273|12|Two Parent|Less than $10,000|||Y|No||Self|General Community||Match Support|F|White||36|28269|Masters Degree|Married|Education|28205|6|6|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|500896588|500896858|3|15|2|500924445|1|0|2|500183434|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1||8735132144641863371|0
M2076|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3044|Green||2008-10-08|2008-11-05|NaT||||100||1|1|1|1|M|Hispanic|Other South American|17|No|Mother|28273|8|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|501023408|501023677|3|15|1|501356600|1|0|1|500296545|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1||0|0
M2077|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|767|Green||2015-01-22|2015-01-30|NaT||||25.2||1|1|1|1|F|Hispanic|Other South American|16|No|Mother|28215|7|Two Parent|$10,000 to $14,999|||Y|Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||30|28211|Masters Degree|Married|Tech: Support, Writing|28202|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503860710|503862704|3|15|2|504115693|1|0|2|500809450|10|2|-2||2|1|500011312|-2||-2|0|10|||17159|12|||1||8202428416367135871|0
M2078|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|770|Yellow|PERL 2014-2016|2015-01-16|2015-01-27|NaT||||25.3||2|2|1|1|F|Hispanic|Other South American|14|No|Mother|28212|8|Two Parent|Unknown||||Yes|Big|Neighbor/Friend|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|Hispanic||26|28215|Bachelors Degree|Single|Student: College||0|0|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|502215233|502215660|3|15|2|504119825|3|0|2|500808734|10|2|-2||2|2|500011312, 500014681|-2|500000294, 500014681|-2|6854|8|||7464|9|||1|500014681|2811191761055817959|0
M2079|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|697|Green||2013-11-04|2013-11-15|2015-10-13|Volunteer: Time constraint|Volunteer: Time constraint||22.9||2|2|1|1|F|Hispanic|Other South American|13|No|Mother|28208|5|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Hispanic||39|28278|Associate Degree|Married|Finance||1|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502485856|502486303|3|15|2|503544124|3|0|2|500726848|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1||3935539763241716148|0
M2080|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|3856|Green||2005-03-30|2005-03-30|2015-10-20|Child/Family: Time constraints|Child/Family: Time constraints||126.7||1|2|1|2|F|Multi-Race (None of the above)||19|No|Father|28208|10|Two Parent|Unknown||||No||Self|General Community||Match Support|F|White||45|28226|Bachelors Degree||Business: Human Resources||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|500186798|500187961|7|0|2|500189825|1|0|2|500037945|10|1|-1||4|1||-2||-2|0|10|||7464|9|||1||702163000107564368|0
M2081|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|3123|Green||2007-11-14|2007-11-27|2016-06-15|Child: Graduated|Child: Graduated||102.6||3|4|1|2|F|Black||19||Mother|28208|3|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|White||37|28012|Some College|Married|Finance: Banking|28208|8|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|500771746|500772014|31|0|2|500996153|1|0|2|500218182|10|1|500000295|2128173567|4|1||-2||-2|0|4|||7464|9|||1||46835895261850668|0
M2082|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2266|Yellow||2008-11-05|2008-11-21|2015-02-04|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||74.4||1|2|2|3|F|White||18|No|Mother|28031|5|Other/Unknown|Unknown||||No||School|General Community||Match Support|F|White||68|28036||Divorced|Business: Sales||5|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500011349|501513669|501513961|1|0|2|500824400|1|0|2|500310460|10|1|-1||4|2||-2||-2|0|4|||7464|9|||1||927920773840777760|0
M2083|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2597|Green||2009-03-19|2009-03-20|2016-04-29|Child: Graduated|Child: Graduated||85.3||1|2|1|2|F|Black||18|No|Mother|28216|11|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|F|Black||38|28269|Masters Degree|Single|Medical: Nurse|28262|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018851|501609876|501610196|31|0|2|501425392|31|0|2|500350904|10|1|500000295|2128190544|4|1|500004640|-2||-2|0|4|||7464|9|||1||2374609189072499123|7044657180546140448
M2084|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|3599|Green||2007-04-30|2007-04-30|NaT||||118.2||1|2|1|2|M|Black||18||Mother|28213|9|Other/Unknown|Unknown||||No||School|General Community||Match Support|F|Black||38|28213||Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500881634|500881903|31|0|1|500816190|31|0|2|500174321|10|1|500000295|2128173562|2|1||-2||-2|0|4|||46|2|||1||253338316288302752|0
M2085|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|882|Green||2014-10-07|2014-10-07|NaT||||29||1|2|1|2|F|Hispanic||18|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|F|Some Other Race||34|28216|Masters Degree|Living w/ Significant Other|Finance|28202|0|0|Local Print|Media|Big|General Community|mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504043329|504045347|3|0|2|503918707|41|0|2|500781130|10|1|500014504||2|1|500014505, 500014506|-2|500014506|-2|0|4|||7439|1|||1||702163000107564368|0
M2086|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|3542|Green||2007-02-27|2007-03-01|2016-11-10|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||116.4||1|2|1|2|M|Black||17||Mother|28217|9|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|Multi-Race (None of the above)||38|29710|Bachelors Degree|Single|Architect||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|500835156|500835425|31|0|1|500466903|7|0|1|500163828|10|1|500000295|2128173557|4|1||-2||-2|0|4|||46|2|||1||7501346876523517480|0
M2087|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2549|Green||2008-10-15|2008-10-22|2015-10-15|Volunteer: Moved|Volunteer: Moved||83.7||2|3|1|2|F|Black||17||Mother|28213|9|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|White||35|85254|Bachelors Degree|Married|Medical: Admin|28217|2|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|501132052|501076355|31|0|2|501356464|1|0|2|500299659|10|1|500000295|2128173561|4|1||-2||-2|0|4|||7446|3|||1||7960300212314874874|0
M2088|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2591|Green||2007-12-12|2007-12-12|2015-01-15|Child: Family structure changed|Child: Family structure changed||85.1||1|2|4|6|F|Black||17||Mother|28217|8|Two Parent|Unknown||||No||School|General Community||Match Support|F|Black||48|28273|Bachelors Degree|Married|Business: Mgt, Admin|28273|4|0|Recruitment Event|Neighbor/Friend|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500018987|501129781|501130055|31|0|2|500189245|31|0|2|500230585|10|1|500000295|2128190544|4|1||-2||-2|0|4|||7459|10|||1||8981704271528751143|0
M2089|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2414|Yellow||2008-12-18|2009-01-14|2015-08-25|Child: Lost interest|Child: Lost interest||79.3||1|2|1|2|F|Black||17||Mother|28031|10|Other/Unknown|Unknown||||No||School|General Community||Match Support|F|Black||36|28205|Bachelors Degree|Single|Business: Mgt, Admin|28036|0|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|501488919|501489205|31|0|2|501392684|31|0|2|500328107|10|1|-1||4|2||-2||-2|0|4|||7464|9|||1||3455806768141331471|0
M2090|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|882|Green||2014-10-07|2014-10-07|NaT||||29||1|2|1|2|F|Black||17|No|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|Black||27|28202|Masters Degree|Single|Business|28202|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500017732|504042339|504044357|31|0|2|503984783|31|0|2|500781137|10|1|500014504||2|1||-2|500014506|-2|0|4|||7462|13|||1||702163000107564368|0
M2091|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|753|Green||2014-10-06|2014-10-06|2016-10-28|Child/Family: Moved|Child/Family: Moved||24.7||1|2|1|2|F|White||17|No|Mother|28217|9|One Parent: Female|Unknown|||Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|F|White||44|28226|Masters Degree|Single|Human Services: Social Worker|28226|0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017786|504043224|504045242|1|0|2|503985439|1|0|2|500780901|10|1|500014504||4|1|500014505, 500014506|-2||-2|0|4|||7462|13|||1||702163000107564368|0
M2092|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2183|Red||2010-10-28|2010-11-16|2016-11-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||71.7||3|4|1|2|F|White||17|No|GrandFather|28147|10|Grandparents|Unknown||||No||School|General Community|Cabarrus County|Match Support|F|White||29|28078||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500022817|501160242|501160516|1|0|2|502325100|1|0|2|500487111|10|1|-1||4|3|500016374|-2|500016374|-2|0|4|||7496|10|||1||0|0
M2093|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|753|Yellow||2014-10-06|2014-10-06|2016-10-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||24.7||1|2|1|2|F|Black||17|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|F|White||31|28278|Bachelors Degree|Married|Business: Mgt, Admin|28202|4|0|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017786|504043260|504045278|31|0|2|503969480|1|0|2|500780787|10|1|500014504||4|2|500014505, 500014506|-2|500014506|-2|0|4|||7462|13|||1||702163000107564368|0
M2094|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1952|Green|Amachi|2011-02-14|2011-02-15|2016-06-20|Child: Lost interest|Child: Lost interest||64.1||1|2|4|5|F|Black||16|Yes|Mother|28206|10|One Parent: Female|Unknown||||Yes||School|General Community|Amachi|Match Support|F|Black||52|28216|Some College|Divorced|Business: Clerical|28202|16|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|502445356|502445803|31|0|2|501026290|31|0|2|500517278|10|1|500000295|2128173561|4|1|500000294|-2||-2|0|4|||46|2|||1|500000294|2374609189072499123|0
M2095|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|882|Green||2014-10-07|2014-10-07|NaT||||29||1|2|1|2|M|Black||16|Yes|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|M|White||26|28210|Bachelors Degree||Business|28281|0|5|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504043128|504045146|31|0|1|503985272|1|0|1|500781233|10|1|500014504||2|1|500014505, 500014506|-2|500014506|-2|0|4|||7462|13|||1||702163000107564368|0
M2096|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|882|Green||2014-10-07|2014-10-07|NaT||||29||1|2|1|2|M|Black||16|No|Mother|28208|9|One Parent: Female|Unknown|||Y|Yes||School|General Community|mentor2.0, mentor2.0 2014|Match Support|M|White||60|28211|Masters Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|0|1|277|60|598|500000170|500022907|504043397|504045415|31|0|1|503922094|1|0|1|500781234|10|1|500014504||2|1|500014505, 500014506|-2|500014506|-2|0|4|||7671|13|||1||702163000107564368|0
M2097|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1593|Green||2012-10-26|2012-10-26|NaT||||52.3||1|2|1|2|F|Black||16|No|Mother|28217|11|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|White||48|28078|Some College|Married|Finance|28217|7|0|LPL Financial|Workplace Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503239475|503241272|31|0|2|503162880|1|0|2|500651859|10|1|500009132|2128207319|2|1||-2||-2|0|4|||11247|3|1204|3|1||253338316288302752|0
M2098|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|3736|Green||2006-12-14|2006-12-14|NaT||||122.7||2|3|4|5|M|Black||16||GrandMother|28208|6|Grandparents|Unknown||||No||School|General Site||Match Support|M|Black||49|28217|Associate Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site||Match Support|1|0|0|1|277|60|598|500000170|500017732|500337327|500251937|31|0|1|500189300|31|0|1|500148261|10|1|500000295|2128173561|2|1||-1||-1|0|4|||7464|9|||1||5424205421938369753|0
M2099|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|3964|Red||2006-04-19|2006-04-19|2017-02-24|Child: Graduated|Child: Graduated||130.2||1|2|1|2|F|Black||16||Mother|28208|0|One Parent: Female|Unknown||||No||School|General Site||Match Support|F|White||34|28210|Bachelors Degree|Single|Business: Mgt, Admin|29715|0|0|Radio|Media|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500008321|500399844|500400094|31|0|2|500188569|1|0|2|500089058|10|1|500000295|2128173567|4|3||-1||-1|0|4|||131|1|||1||46835895261850668|0
M2100|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|498|Green|mentor2.0, mentor2.0 2015|2015-09-23|2015-10-26|NaT||||16.4||1|2|2|3|M|White||16|No|Mother|28208|10|Two Parent|Unknown||||Yes||School|General Community|mentor2.0, mentor2.0 2015|Match Support|M|White||33|28202|Bachelors Degree|Married|Finance|28202|0|2|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0, mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500022907|504419889|504422142|1|0|1|503976384|1|0|1|500841736|10|1|500014504||2|1|500014505, 500015184|-2|500014505, 500014506|-2|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M2101|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1957|Green||2011-10-27|2011-10-28|NaT||||64.3||1|2|1|2|F|American Indian or Alaska Native||16|No|Aunt|28027|8|One Parent: Male|Unknown||||Yes||School|General Community|Cabarrus County|Match Support|F|White||49|28027|Bachelors Degree|Married|Business: Marketing|28025|14|0|ACN|Workplace Partner|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|502785308|504347632|6|0|2|502736971|1|0|2|500571594|10|1|500000295|2128212919|2|1|500016374|-2|500016374|-2|0|4|||13581|3|||1||5273065343662533495|1791051703918408849
M2102|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|479|Green|mentor2.0, mentor2.0 2014|2014-10-06|2014-10-06|2016-01-28|Child/Family: Moved|Child/Family: Moved||15.7||1|2|1|2|F|Black||16|No|Father|28216|9|One Parent: Male|Unknown|||Y|Yes||School|General Community||Match Support|F|Black||27|28269|Bachelors Degree|Single|Finance||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500017732|504043170|504045188|31|0|2|503974104|31|0|2|500780783|10|1|500014504||4|1||-2|500014506|-2|0|4|||7462|13|||1|500014505, 500014506|7301546317881317703|0
M2103|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|487|Green|mentor2.0, mentor2.0 2015|2015-10-12|2015-11-06|NaT||||16||1|2|1|2|F|Hispanic||16|No|Mother|28217||One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||33|28031||Married|Journalist/Media|28031|0|0|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|504445232|504447488|3|0|2|504431681|1|0|2|500846712|10|1|500014504||2|1||-2|500015184|-2|0|4|||7462|13|||1|500014505, 500015184|702163000107564368|0
M2104|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1732|Red|Amachi|2010-11-24|2010-12-03|2015-08-31|Volunteer: Time constraint|Volunteer: Time constraint||56.9||2|3|4|6|M|White||16|Yes|Mother|28146|8|One Parent: Female|Unknown||||Yes||School|General Community|Amachi|Match Support|M|White||41|28078|Bachelors Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|502034298|502034697|1|0|1|500188638|1|0|1|500499336|10|1|500004954||4|3|500000294|-2|500000294|-2|0|4|||7464|9|||1|500000294|0|0
M2105|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2029|Red|Project Big|2010-03-22|2010-03-31|2015-10-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||66.7||1|2|1|2|F|Black||16||Mother|28213|8|Other/Unknown|Unknown||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28262|||Business: Mgt, Admin|75234|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|502137546|502137975|31|0|2|501641708|31|0|2|500442568|10|1|500000295|2128173560|4|3|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640|5441374193599827162|0
M2106|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1888|Green|Project Big|2011-10-27|2011-12-29|2017-02-28|Volunteer: Moved|Volunteer: Moved||62||1|2|5|6|M|Black||16||Mother|28208|8|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Black|Other African|53|28277||Married|Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|502763586|502764498|31|0|1|500189754|31|31|1|500571093|10|1|500000295|2128173561|4|1||-2||-2|0|4|||7464|9|||1|500004640|4440360203097874486|0
M2107|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|3388|Yellow||2007-11-27|2007-11-27|NaT||||111.3||1|2|1|2|F|White||16||Mother|28270|1|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|White||55|28277|Masters Degree|Widowed|Consultant||5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501101149|501101423|1|0|2|500834694|1|0|2|500223542|10|1|500000295|2128183289|2|2||-2||-2|0|4|||7671|13|||1||7554307376683929204|0
M2108|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2520|Red|2010-2012 OJJDP JJI|2009-01-27|2009-02-13|2016-01-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||82.8||1|2|1|2|M|Hispanic||16||Mother|28031|5|Other/Unknown|Unknown||||No||School|General Community||Match Support|M|White||65|28031|Some College|Married|Tech: Sales, Mktg|4241|5|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017777|501618024|501618344|3|0|1|501500078|1|0|1|500336213|10|1|||4|3||-2||-2|0|4|||7462|13|||1|500005291|927920773840777760|0
M2109|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1191|Green||2013-10-22|2013-12-02|NaT||||39.1||1|2|1|2|F|Black||16|No|Mother|28205|9|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|Black||46|28214|Associate Degree|Married|Business|28202|2|10|Duke Energy|Workplace Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|503633704|503635645|31|0|2|503604638|31|0|2|500721771|10|1|500009132|2128173561|2|1||-2||-2|0|4|||16705|3|||1||2374609189072499123|0
M2110|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|493|Green||2015-10-16|2015-10-31|NaT||||16.2||1|2|2|3|F|Black||16|No|Mother|28217|9|Two Parent|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|Black||53|28226|Bachelors Degree|Single|Business: Mgt, Admin|28217|2|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500017732|504416193|504418445|31|0|2|504394474|31|0|2|500848798|10|1|500009132|2128207319|2|1||-2||-1|0|4|||11247|3|||1||702163000107564368|0
M2111|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|2345|Green||2010-09-13|2010-10-05|NaT||||77||1|2|1|2|M|Black||15|No|Mother|28031|8|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|Black||53|28078|PHD|Married|Medical|28078|2|0|AA Task Force|Special Event|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|502300563|502300995|31|0|1|502101059|31|0|1|500470033|10|1|-1||2|1||-2||-2|0|4|||11098|8|||1||4112464363801619560|0
M2112|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|2210|Green|Amachi|2011-02-14|2011-02-17|NaT||||72.6||1|2|1|2|M|Black||15|Yes|Mother|28206|9|One Parent: Female|Unknown||||Yes||School|General Community|Amachi|Match Support|M|White||34|28078|Bachelors Degree|Married|Business: Engineer|28202|12|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|502445373|502445803|31|0|1|502453180|1|0|1|500517348|10|1|500000295|2128173561|2|1|500000294|-2|500000294|-2|0|4|||7446|3|||1|500000294|702163000107564368|0
M2113|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|475|Green|mentor2.0, mentor2.0 2015|2015-11-06|2015-11-18|NaT||||15.6||1|2|1|2|F|Black||15|No|Mother|28217|9|One Parent: Female|Unknown||||Yes||School|General Community|mentor2.0 2015|Match Support|F|White||27|28031|Bachelors Degree|Married|Business: Sales|28277|4|0|Self|Self|Big|General Community|mentor2.0 2015|Match Support|0|1|0|1|277|60|598|500000170|500021786|502505660|502506109|31|0|2|504331356|1|0|2|500857003|10|1|500014504||2|1|500015184|-2|500015184|-2|0|4|||7464|9|||1|500014505, 500015184|702163000107564368|0
M2114|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|2660|Green||2009-11-06|2009-11-24|NaT||||87.4||4|5|1|2|F|Black||15||Aunt|28213|8|One Parent: Female|Unknown||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||40|29715|||Customer Service||2|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|500577150|500214349|31|0|2|501734288|1|0|2|500407385|10|1|500000295|2128173560|2|1|500004640, 500005291|-2||-2|0|4|||7464|9|||1||6381341368426079638|0
M2115|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|493|Green|PERL 2014-2016|2015-10-16|2015-10-31|NaT||||16.2||2|3|2|3|F|Black||15|No|Mother|28217|9|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2016, PERL 2014-2016|Match Support|F|Black||29|28209||Single|Customer Service|28217|0|6|Current/Previous Big|Other Big|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500017732|504416147|504418399|31|0|2|504212639|31|0|2|500848801|10|1|500009132|2128207319|2|1|500014505, 500014681, 500016394|-1|500014505, 500016394|-1|0|4|||17159|12|||1|500014681|702163000107564368|0
M2116|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1166|Red||2013-10-29|2013-11-18|2017-01-27|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38.3||1|2|1|2|M|Black||15|No|Mother|28206|7|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|White||31|28205|Masters Degree|Single|Business|28262|8|0|Duke Energy|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503635533|503580712|31|0|1|503604414|1|0|1|500724441|10|1|500009132|2128173561|4|3||-2||-2|0|4|||16705|3|||1||7960300212314874874|7044657180546140448
M2117|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|C|Completed|Match Support|374|Green|PERL 2014-2016|2015-07-15|2015-07-28|2016-08-05|Volunteer: Time constraint|Volunteer: Time constraint||12.3||1|3|1|3|F|Black||15|No|Mother|28208|8|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|Multi-race (Black & White)||41|28216||Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community|mentor2.0|Match Support|0|1|1|0|277|60|598|500000170|500008321|504308876|504311094|31|0|2|504215512|36|0|2|500833533|10|2|-2||4|1|500014681|-2|500014505|-2|34|2|||46|2|||1|500014681|3769714153336154386|2806833304218536184
M2118|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|393|Green||2016-02-04|2016-02-08|NaT||||12.9||1|2|2|3|F|Black||15|No|Mother|28216|8|One Parent: Female|$10,000 to $14,999||||Yes||School|General Community||Match Support|F|Black||30|28217|Bachelors Degree|Single|Business|28217|0|9|LPL Financial|Workplace Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|504579590|504581924|31|0|2|504397175|31|0|2|500877584|10|1|500009132|2128207319|2|1||-2||-2|0|4|||11247|3|||1||3935539763241716148|0
M2119|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2872|Green||2007-12-18|2007-12-18|2015-10-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||94.4||1|2|1|2|M|Black||14||Mother|28217|K|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||45|28273|Masters Degree|Single|Tech: Research/Design||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500017777|501129794|501130068|31|0|1|500922570|31|0|2|500232070|10|1|500000295|2128173557|4|1||-2||-2|0|4|||46|2|||1||8981704271528751143|0
M2120|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1870|Green||2012-01-11|2012-01-23|NaT||||61.4||1|2|1|2|F|White||14|No|Mother|28031|7|Two Parent|Unknown||||Yes||School|General Community||Match Support|F|White||61|28031|Bachelors Degree|Divorced|Business: Mgt, Admin||5|0|Newspaper|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502813454|502814731|1|0|2|502855397|1|0|2|500590919|10|1|500000295|2128173570|2|1||-2||-2|0|4|||129|1|||1||3974159976843499574|0
M2121|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1201|Green||2013-10-17|2013-11-15|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||39.5||1|2|2|3|F|Black||14|No|Father|28205|6|One Parent: Male|Unknown||||Yes||School|General Community||Match Support|F|White||49|28278|Masters Degree|Single|Business|28202|12|0|Duke Energy|Workplace Partner|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500017732|503624326|503626215|31|0|2|503605964|1|0|2|500720641|10|1|500009132|2128173561|4|1||-2||-1|0|4|||16705|3|||1||7960300212314874874|0
M2122|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|887|Yellow|PERL 2014-2016|2014-09-18|2014-09-25|2017-02-28|Volunteer: Time constraint|Volunteer: Time constraint||29.1||1|2|1|2|F|Black||14|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Community|PERL 2014-2016|Match Support|F|White||31|28211|Masters Degree|Single|Finance: Accountant|28202|1|0|Duke Energy|Workplace Partner|Big|General Community|PERL 2014-2016|Match Support|1|0|1|0|277|60|598|500000170|500008321|504012972|504014987|31|0|2|503975669|1|0|2|500776788|10|1|500009132|2128173561|4|2|500014681|-2|500014681|-2|0|4|||16705|3|||1|500014681|7960300212314874874|0
M2123|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1008|Green||2012-11-12|2012-11-20|2015-08-25|Child/Family: Moved|Child/Family: Moved||33.1||1|2|1|2|F|White||14|No|Mother|28083||Other/Unknown|Unknown||||No||School|General Community||Match Support|F|Some Other Race||44|28107|Bachelors Degree|Married|Finance|28025|0|0|ACN|Workplace Partner|Big|General Site|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|1|0|1|0|277|60|598|500000170|500012459|503292494|503294318|1|0|2|503216525|41|0|2|500658574|10|1|500000295|2128212919|4|1||-2|500007920, 500011315, 500011316|-1|0|4|||13581|3|||1||2437132833506538679|0
M2124|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1845|Green||2012-02-10|2012-02-17|NaT||||60.6||1|2|1|2|F|Black||14|No|Mother|28031|6|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||63|28031|Bachelors Degree|Married|Retired||0|0|Local Print|Media|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502813470|503507249|31|0|2|502889718|1|0|2|500597658|10|1|500000295|2128173570|2|1||-2||-2|0|4|||7439|1|||1||3974159976843499574|0
M2125|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1503|Green||2012-03-09|2012-03-23|2016-05-04|Child: Lost interest|Child: Lost interest||49.4||1|2|1|2|F|White||13|No|Non-Relative: Other|28164|4|Other/Unknown|Unknown||||Yes||School|General Community||Match Support|F|White||39|28031|Bachelors Degree|Single|Arts, Entertainment, Sports|28031|5|6|Local Print|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020752|502813513|502814790|1|0|2|502915648|1|0|2|500603223|10|1|500000295|2128173570|4|1||-2||-2|0|4|||7439|1|||1||0|1941858260967385324
M2126|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|523|Green||2015-09-22|2015-10-01|NaT||||17.2||2|3|1|2|F|Black||13|No|Mother|28217|8|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|Black||43|28075|Masters Degree|Divorced|Finance: Tax/Preparer|28202|6|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|504401898|504404140|31|0|2|504350243|31|0|2|500841372|10|1|500009132|2128212899|2|1||-2||-2|0|4|||7462|13|||1||7276767778509034039|0
M2127|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1969|Green||2011-10-10|2011-10-16|NaT||||64.7||1|2|1|2|F|Black||13|No|Mother|28206|8|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||31|28202|Bachelors Degree|Single|Retail: Mgt|28273|6|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|502776341|502777520|31|0|2|502631040|1|0|2|500563165|10|1|500000295|2128173557|2|1||-2||-2|0|4|||7464|9|||1||932861092942387634|0
M2128|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|385|Green||2014-09-04|2014-09-25|2015-10-15|Volunteer: Time constraint|Volunteer: Time constraint||12.6||1|2|1|2|F|Hispanic||13|No|Father|28216|5|Sibling Guardian|Unknown||||Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|Hispanic||28|28214|Bachelors Degree|Single|Business: Clerical|28214|2|9|Duke Energy|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500018987|503610353|503612230|3|0|2|503973144|3|0|2|500774532|10|1|500009132|2128173561|4|1|500011312|-2||-2|0|10|||16705|3|||1||7960300212314874874|0
M2129|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|896|Green||2014-09-12|2014-09-23|NaT||||29.4||1|2|2|3|F|Black||13|No|Mother|28206|5|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|Black||27|28213|Bachelors Degree|Single|Finance|28202|0|5|Ally Financial|Workplace Partner|Big|General Site||Match Support|1|0|0|1|277|60|598|500000170|500017732|503996726|503998741|31|0|2|503355514|31|0|2|500775721|10|1|500009132|2128173561|2|1||-2||-1|0|4|||12831|3|||1||7960300212314874874|0
M2130|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1073|Yellow||2012-04-17|2012-04-17|2015-03-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.3||2|3|1|2|F|American Indian or Alaska Native||13|No|Aunt|28027|3|Other Relative|Unknown||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||38|28027|Some College|Single|Arts, Entertainment, Sports|28025|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503012569|504347632|6|0|2|502966672|1|0|2|500610298|10|1|500000295|2128212919|4|2|500014681, 500016374|-2||-2|0|4|||7496|10|1360|3|1||2437132833506538679|1791051703918408849
M2131|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|519|Green||2015-09-21|2015-10-05|NaT||||17.1||1|2|2|3|M|Hispanic||13|No|Mother|28217|7|Two Parent|$15,000 to $19,999||||Yes||School|General Community|PERL 2014-2016|Match Support|M|Hispanic||34|28205|Masters Degree|Divorced|Tech: Engineer|28202|8|0|Duke Energy|Workplace Partner|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500018851|504396299|504398539|3|0|1|503973970|3|0|1|500841080|10|1|500009132|2128212899|2|1|500014681|-2|500014681|-2|0|4|||16705|3|||1||7276767778509034039|0
M2132|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1033|Green||2012-11-15|2012-11-16|2015-09-15|Child/Family: Moved|Child/Family: Moved||33.9||1|2|1|2|M|White||13|No|GrandMother|28083||Grandparents|Unknown||||No||School|General Community||Match Support|M|White||57|28027||Married|Business: Sales|28025|3|0|ACN|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503292427|503248831|1|0|1|503282196|1|0|1|500660366|10|1|500000295|2128212919|4|1||-2||-2|0|4|||13581|3|||1||2437132833506538679|0
M2133|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1206|Red||2012-10-30|2012-10-30|2016-02-18|Volunteer: Moved|Volunteer: Moved||39.6||2|3|2|3|M|Black||13|No|Mother|28031|6|Other/Unknown|Unknown||||Yes||School|General Community||Match Support|M|White||32|28078|Bachelors Degree||Business: Marketing|28031|2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|503250358|503252163|31|0|1|501721806|1|0|1|500653597|10|1|500000295|2128173570|4|3||-2||-2|0|4|||7464|9|||1||3974159976843499574|0
M2134|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1126|Red||2014-01-17|2014-01-27|2017-02-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||37||1|2|1|2|F|Hispanic||13|No|Mother|28217|3|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|White||45|28273|Some College|Single|Business|28217|2|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500020753|503779471|503781448|3|0|2|503040015|1|0|2|500743583|10|1|500000295|2128173557|4|3||-2||-2|0|4|||7464|9|||1||8981704271528751143|0
M2135|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|477|Green||2015-10-27|2015-11-16|NaT||||15.7||2|3|1|2|M|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Asian||26|28202|Bachelors Degree|Single|Finance: Banking|28202|2|9|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|503610226|503612103|31|0|1|504260675|4|0|1|500852497|10|1|500000295|2128173561|2|1||-2|500007920, 500011315, 500011316|-2|0|4|||7462|13|||1||7960300212314874874|0
M2136|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1943|Green||2011-11-02|2011-11-11|NaT||||63.8||1|2|1|2|F|Black||12|No|Mother|28031|5|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||62|28031|Masters Degree|Married|Real Estate: Realtor|28031|8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502813527|502814804|31|0|2|502691411|1|0|2|500573720|10|1|500000295|2128173570|2|1||-2||-2|0|4|||7496|10|||1||8034889377453131101|0
M2137|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1092|Green||2014-02-27|2014-03-11|NaT||||35.9||1|2|1|2|F|Black||12|Yes|Mother|28217|4|One Parent: Female|Unknown||||Yes||School|General Community|Amachi|Match Support|F|Black||78|28273|Masters Degree|Widowed|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|503807530|503809507|31|0|2|503381588|31|0|2|500751801|10|1|500000295|2128173557|2|1|500000294|-2||-2|0|4|||7464|9|||1||8981704271528751143|0
M2138|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|1035|Yellow||2012-11-29|2012-11-30|2015-10-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||34||1|2|1|2|F|Black||12|No|GrandMother|28027||Grandparents|Unknown||||Yes||School|General Community||Match Support|F|Black||46|28025||Divorced|Finance: Banking||0|0|ACN|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|503292675|503294499|31|0|2|503282391|31|0|2|500664592|10|1|500000295|2128212924|4|2||-2||-2|0|4|||13581|3|||1||3232906304025417619|0
M2139|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|519|Green||2015-09-22|2015-10-05|NaT||||17.1||1|2|2|3|F|White||12|No|Mother|28210|7|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|White||29|28209|Bachelors Degree|Single|Finance|28202|5|0|Duke Energy|Workplace Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|504396213|504398453|1|0|2|503615576|1|0|2|500841374|10|1|500009132|2128212899|2|1||-2||-2|0|4|||16705|3|||1||8568001799025358453|0
M2140|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|772|Yellow||2013-04-08|2013-04-10|2015-05-22|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||25.4||1|2|1|2|F|Black||12|No|Mother|28031|5|Other/Unknown|Unknown||||Yes||School|General Community||Match Support|F|White||56|28036|Bachelors Degree|Single|Arts, Entertainment, Sports||0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|503249895|503251700|31|0|2|503372833|1|0|2|500691940|10|1|500000295|2128173570|4|2||-2||-2|0|4|||7464|9|||1||8034889377453131101|0
M2141|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|2297|Green||2010-11-09|2010-11-22|NaT||||75.5||1|2|2|3|M|Black||12|No|Mother|28215|4|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||52|28207||Married|Medical: Doctor, Provider||0|0|Omega Psi Phi|Fraternity/Sorority|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502290745|502291177|31|0|1|501944716|31|0|1|500492413|10|1|500000295|2128173561|2|1||-2||-2|34|2|||8694|14|||1||2417657944362725638|0
M2142|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|711|Green||2015-03-02|2015-03-27|NaT||||23.4||1|2|1|2|M|Black||12|No|Mother|28216|5|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||36|28078|Masters Degree|Married|Finance: Banking|28205|1|4|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504183436|504185545|31|0|1|504053150|1|0|1|500816353|10|1|500000295|2128173561|2|1||-2||-2|0|4|||7439|1|||1||7960300212314874874|0
M2143|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|480|Red|PERL 2014-2016|2015-11-09|2015-11-13|NaT||||15.8||1|2|1|2|F|Black||12|No|Mother|28027|4|Other/Unknown|Unknown||||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||24|28216||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500022817|504198005|504200116|31|0|2|504222771|31|0|2|500857505|10|1|500000295|2128212924|2|3|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||46|2|||1|500014681|3232906304025417619|0
M2144|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|2195|Yellow|Amachi|2010-10-26|2010-10-28|2016-10-31|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||72.1||1|2|1|2|F|Black||11|Yes|Mother|28203|K|One Parent: Female|Unknown||||Yes||School|General Community|Amachi|Match Support|F|White||32|28226|||Consultant||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|502369374|501376144|31|0|2|501876592|1|0|2|500485591|10|1|-1||4|2|500000294|-2||-2|0|4|||7464|9|||1|500000294|8568001799025358453|0
M2145|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|684|Green||2015-04-20|2015-04-23|NaT||||22.5||1|2|1|2|F|Black||11|No|Mother|28208|5|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||53|28173|Some College|Divorced|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504257276|504259420|31|0|2|504250952|1|0|2|500824001|10|1|500000295|2128173557|2|1||-2||-2|0|4|||17159|12|||1||8981704271528751143|0
M2146|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Match Support|585|Green||2015-01-22|2015-02-23|2016-09-30|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||19.2||1|2|1|2|M|Black||10|No|Mother|28217|3|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||67|28104||Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|504184625|504186734|31|0|1|504016261|1|0|1|500809549|10|1|500000295|2128173557|4|1||-2||-2|0|4|||17159|12|||1||8981704271528751143|0
M2147|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Completed|Pending Match|1175|Red||2013-11-07|2013-11-19|2017-02-06|Volunteer: Time constraint|Volunteer: Time constraint||38.6||1|3|1|2|F|White||9|No|Mother|28025|3|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Cabarrus County|Pending Match|F|White||68|28025||Married|Retired||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500022817|503694497|503696462|1|0|2|503550540|1|0|2|500728658|9|1|500000295|2128212919|4|3|500016374|-2|500016374|-2|0|4|||7464|9|||1||4085045877112350207|0
M2148|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|96|Green|Cabarrus County|2016-11-17|2016-12-01|NaT||||3.2||1|2|2|3|F|White||9|No|Mother|28083|4|Two Parent|$30,000 to $34,999||||Yes||School|General Community|Cabarrus County|Match Support|F|Black||28|28083|Bachelors Degree|Single|Law|28147|0|2|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504936816|504939367|1|0|2|504528677|31|0|2|500928981|10|1|500000295|2128232374|2|1|500016374|-2|500016374|-2|0|4|||7496|10|||1|500016374|2043334928777030191|0
M2149|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|739|Green||2015-02-27|2015-02-27|NaT||||24.3||1|2|1|2|F|Hispanic||9||Mother|28031|4|Two Parent|Unknown||||Yes||School|General Community||Match Support|F|White||52|28036|Bachelors Degree|Divorced|Finance||1|3|TV|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500020910|504220499|504222613|3|0|2|504045698|1|0|2|500816057|10|1|500000295|2128173570|2|1||-2|500007920, 500011315, 500011316|-2|0|4|||130|1|||1||8034889377453131101|0
M2150|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|C|Active|Match Support|1256|Green||2013-09-12|2013-09-28|NaT||||41.3||1|3|1|3|F|Black||9|Yes|Mother|28205||One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community|Amachi|Match Support|F|White||33|28205|Masters Degree|Single|Education: Admin|28027|0|5|Recruitment Event|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|503457000|503458866|31|0|2|503552518|1|0|2|500710586|10|2|500014421||2|1|500000294|-2||-2|0|10|||7460|12|||1||0|4899444095790462270
M2151|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|335|Green||2016-04-01|2016-04-06|NaT||||11||1|2|1|2|F|Hispanic||7|No|Mother|28036|1|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||30|28031|Bachelors Degree|Single|Business: Sales|53158|3|9|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|504449667|504451923|3|0|2|504633714|1|0|2|500887478|10|1|500000295|2128173570|2|1||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||8034889377453131101|5081726734274569781
M2152|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|Y|S|Active|Match Support|1943|Green||2011-11-02|2011-11-11|NaT||||63.8||1|2|1|2|M|Hispanic|Mexican|15|No|Mother|28031|7|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28036|Some College|Married|Self-Employed, Entrepreneur|28036|20|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|502813442|502814719|3|10|1|502656402|1|0|1|500573668|10|1|500000295|2128173570|2|1|500005291|-2||-2|0|4|||7671|13|||1||3974159976843499574|0
