InterviewNum|AgencyName|AgencyGroup|OfficeName|TeamName|MatchType|MatchStatus|MatchOpenDate|MatchCloseDate|SurveyType|YOSScheduledDate|YOSCompletionDate|YOSCompletionType|YOSStatus|Q1|Q2Neg|Q3Neg|Q4Neg|Q5|Q6|SocAccept|Q1b|Q2b|Q3b|Q4b|Q5b|Q6b|SocAcceptB|SocAcceptPrcnt|Q7Neg|Q8|Q9|Q10Neg|Q11Neg|Q12|SchComp|Q7b|Q8b|Q9b|Q10b|Q11b|Q12b|SchCompB|SchCompPrcnt|Q13|Q14|Q15|EdExpect|Q13b|Q14b|Q15b|EdExpectb|EdExpectPrcnt|Q16|Q17|Q18|Q19|Grades|Q16b|Q17b|Q18b|Q19b|Gradesb|GradesPrcnt|Q20Neg|Q21Neg|Q22Neg|Q23Neg|Q24Neg|Q25Neg|Q26Neg|RiskAtt|Q20b|Q21b|Q22b|Q23b|Q24b|Q25b|Q26b|RiskAttb|RiskAttPrcnt|Q27|Q28|Q29|PTrust|Q27b|Q28b|Q29b|PTrustb|PTrustPrcnt|Q30Neg|Q31Neg|Truancy|Q30b|Q31b|Truancyb|TruancyPrcnt|Q32|SpAdult|Q32b|SpAdultb|SpAdultPrcnt|Q33Neg|JJustice|Q33b|JJusticeB|JJusticePrcnt|MatchSupportLevel|MatchReportSources|MatchClosureReasons|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildGrade|ChildLivingSituation|ChildIncomeLevel|ChildFamilyAssistance|ChildFreeReducedLunch|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|ChildPartKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolPartKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|MatchKey|MatchTypeKey|SiteTypeKey|MatchActivityKey|SiteKey|StatusKey|MatchSupportLevelKey|MatchReportSourceKey|ChildReportSourceKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|YOSSurveyKey|PriorBaselineYOSSurveyKey|YOSStatusKey|YOSCompletionTypeKey|SurveyTypeKey|CustodialAdultEmployerHash
21|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-26|NaT|Baseline|2015-02-24|2015-02-26|Complete|Done|3|3|4|3|3|3|3.17|||||||||4|4|3|4|4|3|3.67|||||||||4|4|3|3.67||||||4|4|5|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|||24.4||1|1|1|1|M|Black||14|No|Mother|28278|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|Black||29|28209|Bachelors Degree|Single|Finance|20877|0|8|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|504160892|504162947|31|0|1|504171934|31|0|1|500815454|2||-2||2|1|||-2||-2|0|4|||130|1|||1|854521|-1|4|3|44|2876415545463317777
21|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-02-26|NaT|Followup|2016-02-26|2016-05-12|Expired|Late||||||||3|3|4|3|3|3|3.17|||||||||4|4|3|4|4|3|3.67||||||4|4|3|3.67|||||||4|4|5|5|4.5||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|2|2.5||||1|1||||4|4||Green|||24.4||1|1|1|1|M|Black||14|No|Mother|28278|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|Black||29|28209|Bachelors Degree|Single|Finance|20877|0|8|TV|Media|Big|General Community||Match Support|277|60|598|500000170|500018851|504160892|504162947|31|0|1|504171934|31|0|1|500815454|2||-2||2|1|||-2||-2|0|4|||130|1|||1|855224|854521|4|0|45|2876415545463317777
27|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-16|NaT|Followup|2016-03-16|2016-05-16|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||23.8||1|1|1|1|M|Black||10|No|Mother|28211|2|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|M|White||31|28209|Bachelors Degree|Married|Medical|70112|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|503314773|503314167|31|0|1|504176084|1|0|1|500817494|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|979708||4|1|45|4253272603994307857
30|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-26|NaT|Baseline|2015-03-10|2015-03-26|Complete|Done|2|1|2|1|3|4|2.17|||||||||1|4|2|2|3|4|2.67|||||||||2|3|3|2.67||||||4|5|4|5|4.5|||||||3|2|4|4|4|2|2|3||||||||||4|4|3|3.67||||||1|2|1.5|||||1|1||||4|4||||Yellow|||23.5||1|1|1|1|F|Black||11|No|Mother|28227|3|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||29|28226|Bachelors Degree|Single|Finance: Accountant|28202|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|504194601|504184323|31|0|2|504032490|1|0|2|500817776|2||-2||2|2|||-2||-2|0|4|||7464|9|||1|859018|-1|4|3|44|5822555200185981373
30|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-26|NaT|Followup|2016-03-26|2016-04-22|Complete|Done|4|2|3|2|3|4|3|2|1|2|1|3|4|2.17|38.25|3|3|3|3|4|3|3.17|1|4|2|2|3|4|2.67|18.73|4|4|4|4|2|3|3|2.67|49.81|3|3|3|3|3|4|5|4|5|4.5|-33.33|4|4|4|4|4|4|4|4|3|2|4|4|4|2|2|3|33.33|4|4|4|4|4|4|3|3.67|8.99|3|3|3|1|2|1.5|100|2|2|1|1|100|4|4|4|4|0|Yellow|||23.5||1|1|1|1|F|Black||11|No|Mother|28227|3|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||29|28226|Bachelors Degree|Single|Finance: Accountant|28202|0|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500008321|504194601|504184323|31|0|2|504032490|1|0|2|500817776|2||-2||2|2|||-2||-2|0|4|||7464|9|||1|864248|859018|4|3|45|5822555200185981373
33|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-31|NaT|Baseline|2015-03-14|2015-03-31|Complete|Done|1|4|4|3|4|4|3.33|||||||||2|4|3|3|2|2|2.67|||||||||4|4|4|4||||||2|4|3|3|3|||||||4|4|4|4|3|4|3|3.71||||||||||3|3|2|2.67||||||3|2|2.5|||||2|2||||4|4||||Green|||23.3||1|1|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Business: Sales|28277|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|501843066|501843435|31|0|2|504152982|1|0|2|500818696|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|860440|-1|4|3|44|0
33|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-03-31|NaT|Followup|2016-03-31|2016-04-22|Complete|Done|2|3|4|3|4|4|3.33|1|4|4|3|4|4|3.33|0|3|4|3|3|3|3|3.17|2|4|3|3|2|2|2.67|18.73|4|4|4|4|4|4|4|4|0|3|3|3|3|3|2|4|3|3|3|0|4|4|4|4|3|4|4|3.86|4|4|4|4|3|4|3|3.71|4.04|2|3|3|2.67|3|3|2|2.67|0|3|2|2.5|3|2|2.5|0|2|2|2|2|0|4|4|4|4|0|Green|||23.3||1|1|1|1|F|Black||14|No|Mother|28208|6|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Business: Sales|28277|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|501843066|501843435|31|0|2|504152982|1|0|2|500818696|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|866058|860440|4|3|45|0
43|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Baseline|2015-04-24|2015-05-04|Complete|Done|4|2|3|3|3|4|3.17|||||||||2|3|3|3|2|3|2.67|||||||||4|3|3|3.33||||||4|3|2|2|2.75|||||||2|4|4|4|4|4|4|3.71||||||||||4|4|3|3.67||||||2|4|3|||||1|1||||4|4||||Green|||22.2||1|1|1|1|F|White||15|No|Mother|28227|8|One Parent: Female|$35,000 to $39,999||Yes||School|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Law: Paralegal|28211|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504235352|504237484|1|0|2|504200139|1|0|2|500825073|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|873520|-1|4|3|44|8961132295198487522
43|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Followup|2016-05-05|2016-05-09|Complete|Done|3|3|3|3|4|4|3.33|4|2|3|3|3|4|3.17|5.05|2|2|3|2|1|4|2.33|2|3|3|3|2|3|2.67|-12.73|3|3|2|2.67|4|3|3|3.33|-19.82|2|4|4|4|3.5|4|3|2|2|2.75|27.27|3|4|3|1|4|3|3|3|2|4|4|4|4|4|4|3.71|-19.14|3|3|2|2.67|4|4|3|3.67|-27.25|4|4|4|2|4|3|33.33|1|1|1|1|0|4|4|4|4|0|Green|||22.2||1|1|1|1|F|White||15|No|Mother|28227|8|One Parent: Female|$35,000 to $39,999||Yes||School|General Community||Match Support|F|White||26|28205|Bachelors Degree|Single|Law: Paralegal|28211|1|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504235352|504237484|1|0|2|504200139|1|0|2|500825073|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|877359|873520|4|3|45|8961132295198487522
44|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Baseline|2015-04-22|2015-05-04|Complete|Done|2|1|1|1|1|1|1.17|||||||||2|2|2|1|3|2|2|||||||||4|4|4|4||||||2|2|5|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||22.2||1|1|1|1|M|White||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999||Yes||School|General Community||Match Support|M|White||51|28173|Masters Degree|Married|Self-Employed, Entrepreneur|28173|19|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504235369|504237484|1|0|1|503937954|1|0|1|500824366|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|872406|-1|4|3|44|8961132295198487522
44|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-05|NaT|Followup|2016-05-05|2016-05-09|Complete|Done|3|2|1|1|2|3|2|2|1|1|1|1|1|1.17|70.94|2|3|4|2|1|3|2.5|2|2|2|1|3|2|2|25|4|4|4|4|4|4|4|4|0|3|3|3|3|3|2|2|5|5|3.5|-14.29|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|4|3.67|4|4|4|4|-8.25|3|4|3.5|4|4|4|-12.5|2|2|2|2|0|4|4|4|4|0|Green|||22.2||1|1|1|1|M|White||14|No|Mother|28227|6|One Parent: Female|$30,000 to $34,999||Yes||School|General Community||Match Support|M|White||51|28173|Masters Degree|Married|Self-Employed, Entrepreneur|28173|19|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504235369|504237484|1|0|1|503937954|1|0|1|500824366|2||-2||2|1|||-2||-2|0|4|||7464|9|||1|877351|872406|4|3|45|8961132295198487522
45|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-12|NaT|Followup|2016-05-12|2016-05-19|Complete|Done|3|1|2|2|1|4|2.17|||||||||2|1|4|4|4|4|3.17|||||||||2|4|4|3.33||||||4|3|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||21.9||1|1|1|1|F|White||10|No|Mother|28277|4|One Parent: Female|$45,000 to $49,999||Yes||Self|General Community||Match Support|F|White||29|29708|Bachelors Degree|Married|Medical|28105|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500013781|503889301|503891297|1|0|2|504021478|1|0|2|500823483|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|912396||4|3|45|6156547733130613405
46|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-13|NaT|Followup|2016-05-13|2016-05-25|Complete|Done|4|3|4|4|3|4|3.67|||||||||2|4|4|2|1|4|2.83|||||||||4|4|4|4||||||5|4|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||21.9||1|1|1|1|F|White||10|No|Mother|28214|4|One Parent: Female|$10,000 to $14,999|Y|Yes||Relative|General Community||Match Support|F|White||28|28206|Bachelors Degree|Single|Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500013781|504231269|504233379|1|0|2|503927707|1|0|2|500826291|2||-2||2|1|||-2||-2|0|3|||46|2|||1|954853||4|3|45|0
49|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-19|NaT|Followup|2016-05-19|2016-05-18|Complete|Done|4|4|2|4|4|4|3.67|||||||||1|1|4|2|2|4|2.33|||||||||4|3|3|3.33||||||4|5|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|3|2.5|||||1|1||||4|4||||Green|PERL 2014-2016||21.7||1|1|1|1|F|White||10|No|GrandMother|28210|3|Other Relative|Unknown||Yes||Self|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||28|28205|Some College|Single|Transport: Driver|28277|8|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504234369|503470938|1|0|2|504116244|35|0|2|500825294|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|10|||46|2|||1|910429||4|3|45|7044657180546140448
50|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-22|NaT|Baseline|2015-05-22|2015-05-22|Complete|Done|3|1|4|2|3|4|2.83|||||||||3|4|3|3|2|4|3.17|||||||||4|4|4|4||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||21.6||1|1|2|2|F|Black||13|No|Mother|28212|7|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500018851|502930499|502931919|31|0|2|502564910|31|0|2|500828045|2||-2||2|1|||-2||-2|0|10|||17161|11|||1|887615|-1|4|3|44|3402014428779854546
50|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-05-22|NaT|Followup|2016-05-22|2016-08-06|Expired|Late||||||||3|1|4|2|3|4|2.83|||||||||3|4|3|3|2|4|3.17||||||4|4|4|4|||||||4|5|5|4|4.5||||||||||4|4|4|4|4|4|2|3.71||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Green|||21.6||1|1|2|2|F|Black||13|No|Mother|28212|7|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|277|60|598|500000170|500018851|502930499|502931919|31|0|2|502564910|31|0|2|500828045|2||-2||2|1|||-2||-2|0|10|||17161|11|||1|887617|887615|4|0|45|3402014428779854546
54|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Baseline|2015-06-09|2015-06-16|Complete|Done|4|2|4|4|3|3|3.33|||||||||4|4|4|3|2|4|3.5|||||||||4|4|4|4||||||4|3|5|5|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|3|3.67||||||1|2|1.5|||||2|2||||4|4||||Green|PERL 2014-2016||20.8||1|1|1|1|M|Black||15|No|GrandMother|28208|7|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|3|10|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503944459|503946467|31|0|1|504260502|1|0|1|500829606|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7462|13|||1|901862|-1|4|3|44|7044657180546140448
54|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Followup|2016-06-16|2016-08-18|Declined|Late||||||||4|2|4|4|3|3|3.33|||||||||4|4|4|3|2|4|3.5||||||4|4|4|4|||||||4|3|5|5|4.25||||||||||4|4|4|4|3|4|3|3.71||||||4|4|3|3.67|||||1|2|1.5||||2|2||||4|4||Green|PERL 2014-2016||20.8||1|1|1|1|M|Black||15|No|GrandMother|28208|7|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|3|10|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020752|503944459|503946467|31|0|1|504260502|1|0|1|500829606|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7462|13|||1|905636|901862|4|1|45|7044657180546140448
55|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Baseline|2015-05-29|2015-06-16|Complete|Done|3|3|4|3|3|4|3.33|||||||||2|4|3|3|2|4|3|||||||||4|3|4|3.67||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||20.8||1|1|1|1|M|Black||13|No|Mother|28216|6|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Business|28217|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504247189|504249305|31|0|1|504228103|1|0|1|500828700|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|892042|-1|4|3|44|3402014428779854546
55|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-06-16|NaT|Followup|2016-06-16|2016-08-31|Expired|Late||||||||3|3|4|3|3|4|3.33|||||||||2|4|3|3|2|4|3||||||4|3|4|3.67|||||||4|4|3|4|3.75||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||3|3|3||||1|1||||4|4||Green|||20.8||1|1|1|1|M|Black||13|No|Mother|28216|6|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Business|28217|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504247189|504249305|31|0|1|504228103|1|0|1|500828700|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|905690|892042|4|0|45|3402014428779854546
66|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Baseline|2015-07-16|2015-07-27|Complete|Done|3|3|4|4|3|4|3.5|||||||||4|4|4|4|2|4|3.67|||||||||3|3|3|3||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||3|4|3|3.33||||||4|4|4|||||2|2||||4|4||||Green|||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||Relative|General Community||Match Support|F|White||29|28209|Bachelors Degree|Single|Retail: Mgt|28217|3|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504312629|504314787|31|0|2|504262612|1|0|2|500833665|2||-2||2|1|||-2||-2|0|3|||17159|12|||1|916650|-1|4|3|44|237874676114443178
66|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Followup|2016-07-27|2016-09-01|Complete|Done|3|4|4|4|3|4|3.67|3|3|4|4|3|4|3.5|4.86|4|3|4|4|4|4|3.83|4|4|4|4|2|4|3.67|4.36|4|4|4|4|3|3|3|3|33.33|3|4|3|4|3.5|4|5|5|4|4.5|-22.22|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|4|3|3.33|3|4|3|3.33|0|4|4|4|4|4|4|0|2|2|2|2|0|4|4|4|4|0|Green|||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||Relative|General Community||Match Support|F|White||29|28209|Bachelors Degree|Single|Retail: Mgt|28217|3|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504312629|504314787|31|0|2|504262612|1|0|2|500833665|2||-2||2|1|||-2||-2|0|3|||17159|12|||1|918944|916650|4|3|45|237874676114443178
67|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Baseline|2015-07-20|2015-07-27|Complete|Done|4|4|4|4|1|4|3.5|||||||||2|2|2|2|3|2|2.17|||||||||3|3|3|3||||||3|3|5|5|4|||||||4|4|4|4|4|4|4|4||||||||||3|4|4|3.67||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Asian||28|28203|Bachelors Degree|Single|Consultant|28202|1|1|Current/Previous Big|Other Big|Big|General Community|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500008321|504312569|504314787|31|0|2|504208036|4|0|2|500833808|2||-2||2|1|500014681|500014681|-2|500014505, 500015184|-2|0|4|||17159|12|||1|917230|-1|4|3|44|237874676114443178
67|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-07-27|NaT|Followup|2016-07-27|2016-09-01|Complete|Done|4|4|4|4|4|4|4|4|4|4|4|1|4|3.5|14.29|3|4|4|4|4|4|3.83|2|2|2|2|3|2|2.17|76.5|4|3|3|3.33|3|3|3|3|11|4|4|4|3|3.75|3|3|5|5|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|3|3|3|3|3|4|4|3.67|-18.26|3|3|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||19.4||1|1|1|1|F|Black||12|No|Mother|28202|4|One Parent: Female|$30,000 to $34,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Asian||28|28203|Bachelors Degree|Single|Consultant|28202|1|1|Current/Previous Big|Other Big|Big|General Community|mentor2.0, mentor2.0 2015|Match Support|277|60|598|500000170|500008321|504312569|504314787|31|0|2|504208036|4|0|2|500833808|2||-2||2|1|500014681|500014681|-2|500014505, 500015184|-2|0|4|||17159|12|||1|918957|917230|4|3|45|237874676114443178
70|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-13|NaT|Baseline|2015-08-13|2015-08-13|Complete|Done|4|2|3|2|4|4|3.17|||||||||3|3|4|2|3|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|2|2.5|||||2|2||||4|4||||Green|||18.9||1|1|1|1|F|Black||13|No|Mother|28214|6|One Parent: Female|$50,000 to $59,999||Yes||Self|General Community||Match Support|F|White||29|28273|Masters Degree|Married|Finance: Accountant|28210|3|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504328960|504331182|31|0|2|504215323|1|0|2|500836079|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|926159|-1|4|3|44|8503368421346667831
70|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-13|NaT|Followup|2016-08-13|2016-08-22|Complete|Done|4|3|3|2|4|4|3.33|4|2|3|2|4|4|3.17|5.05|3|4|4|4|4|4|3.83|3|3|4|2|3|4|3.17|20.82|4|4|4|4|4|4|4|4|0|5|5|5|5|5|5|5|5|5|5|0|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|3|3|3|3|2|2.5|20|2|2|2|2|0|4|4|4|4|0|Green|||18.9||1|1|1|1|F|Black||13|No|Mother|28214|6|One Parent: Female|$50,000 to $59,999||Yes||Self|General Community||Match Support|F|White||29|28273|Masters Degree|Married|Finance: Accountant|28210|3|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504328960|504331182|31|0|2|504215323|1|0|2|500836079|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|926293|926159|4|3|45|8503368421346667831
71|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-13|NaT|Followup|2016-08-13|2016-09-30|Declined|Late||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||18.9||1|1|1|1|F|Black||10|No|Mother|28216|2|One Parent: Female|$30,000 to $34,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||34|28031||Single|Self-Employed, Entrepreneur||9|8|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500017732|504186133|504188242|31|0|2|504122609|1|0|2|500834256|2||-2||2|1|||-2||-2|34|2|||17159|12|||1|937690||4|1|45|8136849793711030748
72|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-14|NaT|Baseline|2015-07-22|2015-08-14|Complete|Done|2|3|3|3|3|2|2.67|||||||||4|4|4|2|2|4|3.33|||||||||4|4|4|4||||||5|4|4|2|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||2|2||||3|3||||Green|||18.9||1|1|1|1|M|Black||13|No|Mother|28273|6|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|Black||56|28273|Some College|Married|Govt|28228|0|7|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|504284556|504286757|31|0|1|504260574|31|0|1|500834204|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|918085|-1|4|3|44|2392572474128905139
72|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-08-14|NaT|Followup|2016-08-14|2016-09-28|Complete|Done|4|4|4|2|3|3|3.33|2|3|3|3|3|2|2.67|24.72|2|4|3|3|4|3|3.17|4|4|4|2|2|4|3.33|-4.8|4|4|4|4|4|4|4|4|0|3|3|4|3|3.25|5|4|4|2|3.75|-13.33|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|4|3|3.33|4|4|3|3.67|-9.26|2|3|2.5|2|2|2|25|2|2|2|2|0|4|4|3|3|33.33|Green|||18.9||1|1|1|1|M|Black||13|No|Mother|28273|6|One Parent: Female|$35,000 to $39,999||No||Self|General Community||Match Support|M|Black||56|28273|Some College|Married|Govt|28228|0|7|Self|Self|Big|General Community|Amachi|Match Support|277|60|598|500000170|500008321|504284556|504286757|31|0|1|504260574|31|0|1|500834204|2||-2||2|1|||-2|500000294|-2|0|10|||7464|9|||1|926429|918085|4|3|45|2392572474128905139
80|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-16|NaT|Baseline|2015-09-10|2015-09-16|Complete|Done|4|4|4|4|3|4|3.83|||||||||3|4|4|2|4|4|3.5|||||||||3|3|4|3.33||||||4|3|4|2|3.25|||||||4|4|4|3|4|4|4|3.86||||||||||1|1|3|1.67||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016||17.8||1|1|1|1|M|Some Other Race||13|No|Mother|28217|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||38|28205|Masters Degree|Married|Human Services: Social Worker|28204|5|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504155180|501093096|41|0|1|502462446|1|0|1|500839295|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7464|9|||1|932973|-1|4|3|44|358434295995756137
80|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-16|NaT|Followup|2016-09-16|2016-09-19|Complete|Done|4|4|4|4|4|4|4|4|4|4|4|3|4|3.83|4.44|4|4|4|4|2|4|3.67|3|4|4|2|4|4|3.5|4.86|4|2|2|2.67|3|3|4|3.33|-19.82|5|4|5|4|4.5|4|3|4|2|3.25|38.46|4|4|4|4|4|4|3|3.86|4|4|4|3|4|4|4|3.86|0|4|4|1|3|1|1|3|1.67|79.64|3|3|3|4|4|4|-25|1|1|2|2|-50|4|4|4|4|0|Green|PERL 2014-2016||17.8||1|1|1|1|M|Some Other Race||13|No|Mother|28217|5|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||38|28205|Masters Degree|Married|Human Services: Social Worker|28204|5|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500013781|504155180|501093096|41|0|1|502462446|1|0|1|500839295|2||-2||2|1|500014681|500014681|-2|500014681|-2|0|4|||7464|9|||1|934749|932973|4|3|45|358434295995756137
81|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-22|NaT|Followup|2016-09-22|2016-10-31|Declined|Done||||||||3|1|3|1|4|4|2.67|||||||||2|4|3|1|2|2|2.33||||||4|4|4|4|||||||2|5|3|2|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|4|4|||||4|4|4||||1|1||||4|4||Green|PERL 2014-2016||17.6||2|2|1|1|F|Black||13|No|Mother|28205|6|One Parent: Female|Unknown||Yes||School|General Community|PERL 2014-2016|Match Support|F|White||26|28202|Bachelors Degree|Single|Finance: Banking|28262|1|7|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020752|504013056|504015071|31|0|2|504219921|1|0|2|500839610|2||-2||2|1|500014681|500014681|-2||-2|0|4|||17159|12|||1|936088|793476|4|1|45|0
82|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-23|NaT|Followup|2016-09-23|2016-10-31|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|PERL 2014-2016||17.5||2|2|1|1|M|Black||10|No|Mother|28214|2|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Black||25|28227|Bachelors Degree|Single|Insurance|28277|1|2|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|503779386|503781363|31|0|1|504333970|31|0|1|500839160|2||-2||2|1|500014681|500014681|-2||-2|0|4|||7464|9|||1|936510||4|1|45|1546374315672654438
83|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-28|NaT|Followup|2016-09-28|2016-10-26|Complete|Done|1|2|4|2|3|3|2.5|||||||||3|4|3|3|3|3|3.17|||||||||4|4|4|4||||||4||4|||||||||4|4|4|4|3|4|3|3.71||||||||||2|3|2|2.33||||||3|4|3.5|||||2|2||||4|4||||Green|||17.4||3|3|1|1|F|Black||14|No|Mother|28216|7|Two Parent|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|White||43|28269|Masters Degree|Single|Business: Mgt, Admin||0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|502186245|501610196|31|0|2|504248899|1|0|2|500836970|2||-2||2|1|||-2||-2|0|10|||17159|12|||1|938163||4|3|45|7044657180546140448
84|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-29|NaT|Baseline|2015-09-23|2015-09-29|Complete|Done|4|1|4|4|2|4|3.17|||||||||1|3|3|1|1|3|2|||||||||3|2|2|2.33||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||4|3|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||17.3||1|1|1|1|M|Black||11|No|Mother|28214|4|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28273|Bachelors Degree|Single|Insurance|28226|7|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|504153965|504156015|31|0|1|504372591|1|0|1|500841770|2||-2||2|1|500014681|500014681|-2||-2|0|4|||7464|9|||1|936574|-1|4|3|44|0
84|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-09-29|NaT|Followup|2016-09-29|2016-11-28|Declined|Late||||||||4|1|4|4|2|4|3.17|||||||||1|3|3|1|1|3|2||||||3|2|2|2.33|||||||3|3|3|3|3||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||4|3|3.5||||2|2||||4|4||Green|PERL 2014-2016||17.3||1|1|1|1|M|Black||11|No|Mother|28214|4|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28273|Bachelors Degree|Single|Insurance|28226|7|6|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500020752|504153965|504156015|31|0|1|504372591|1|0|1|500841770|2||-2||2|1|500014681|500014681|-2||-2|0|4|||7464|9|||1|938480|936574|4|1|45|0
85|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Baseline|2015-09-24|2015-10-05|Complete|Done|3|2|3|2|4|4|3|||||||||2|4|4|3|3|4|3.33|||||||||3|3|4|3.33||||||5|4|4|3|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|||||||2|2||||4|4||||Green|||17.1||1|1|1|1|F|Black||12|No|Mother|28215|6|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Multi-Race (None of the above)||27|28269|Bachelors Degree|Single|Transport: Flight Attendant|28208|1|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504358312|504320644|31|0|2|504048355|7|0|2|500842174|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|937130|-1|4|3|44|2141487034287122220
85|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Followup|2016-10-05|2016-11-18|Complete|Done|3|3|3|2|4|4|3.17|3|2|3|2|4|4|3|5.67|3|4|4|4|4|3|3.67|2|4|4|3|3|4|3.33|10.21|4|4|4|4|3|3|4|3.33|20.12|4|4|3|4|3.75|5|4|4|3|4|-6.25|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|3|3.67|4|4|4|4|-8.25|3|3|3|3||||2|2|2|2|0|3|3|4|4|-25|Green|||17.1||1|1|1|1|F|Black||12|No|Mother|28215|6|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|F|Multi-Race (None of the above)||27|28269|Bachelors Degree|Single|Transport: Flight Attendant|28208|1|5|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500008321|504358312|504320644|31|0|2|504048355|7|0|2|500842174|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|940717|937130|4|3|45|2141487034287122220
86|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Baseline|2015-09-28|2015-10-05|Complete|Done|4|2|4|1|2|4|2.83|||||||||4|4|3|1|2|2|2.67|||||||||4|4|4|4||||||3|5|5|4|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||1|1||||4|4||||Green|||17.1||1|1|1|1|M|Black||10|No|Mother|28213|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Consultant|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504179804|504181918|31|0|1|504337207|1|0|1|500842586|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|937970|-1|4|3|44|7044657180546140448
86|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-05|NaT|Followup|2016-10-05|2016-12-20|Expired|Late||||||||4|2|4|1|2|4|2.83|||||||||4|4|3|1|2|2|2.67||||||4|4|4|4|||||||3|5|5|4|4.25||||||||||4|4|4|4|4|4|4|4||||||4|4|4|4|||||2|1|1.5||||1|1||||4|4||Green|||17.1||1|1|1|1|M|Black||10|No|Mother|28213|3|One Parent: Female|Less than $10,000|Y|Yes||School|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Consultant|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504179804|504181918|31|0|1|504337207|1|0|1|500842586|2||-2||2|1|||-2||-2|0|4|||17159|12|||1|940706|937970|4|0|45|7044657180546140448
93|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Baseline|2015-09-21|2015-10-30|Complete|Done|4|1|4|2|3|4|3|||||||||1|3|3|2|2|3|2.33|||||||||4|4|4|4||||||1|1|2|2|1.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|1|2|||||2|2||||4|4||||Green|||16.3||1|1|1|1|F|Black||10|No|Mother|28216|4|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|F|Black||31|28216|Bachelors Degree|Single|Arts, Entertainment, Sports|28202|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504345626|504347850|31|0|2|504373316|31|0|2|500845709|2||-2||2|1|||-2||-2|0|10|||46|2|||1|935912|-1|4|3|44|1712849328738258411
93|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Followup|2016-10-30|2016-12-14|Complete|Done|3|2|4|2|3|3|2.83|4|1|4|2|3|4|3|-5.67|2|3|2|2|3|3|2.5|1|3|3|2|2|3|2.33|7.3|4|4|4|4|4|4|4|4|0|2|2|3|2|2.25|1|1|2|2|1.5|50|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|4|4|4|4|4|4|4|4|0|2|2|2|3|1|2|0|2|2|2|2|0|4|4|4|4|0|Green|||16.3||1|1|1|1|F|Black||10|No|Mother|28216|4|One Parent: Female|$35,000 to $39,999||Yes||Self|General Community||Match Support|F|Black||31|28216|Bachelors Degree|Single|Arts, Entertainment, Sports|28202|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|277|60|598|500000170|500008321|504345626|504347850|31|0|2|504373316|31|0|2|500845709|2||-2||2|1|||-2||-2|0|10|||46|2|||1|953778|935912|4|3|45|1712849328738258411
94|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Baseline|2015-10-08|2015-10-30|Complete|Done|2|4|3|2|4|3|3|||||||||2|3|4|4|3|3|3.17|||||||||3|4|3|3.33||||||4|5|2|3|3.5|||||||4|3|2|2|3|4|4|3.14||||||||||3|4|2|3||||||3|3|3|||||2|2||||4|4||||Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016||16.3|Y|1|1|1|1|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28204|Masters Degree|Married|Consultant||0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504254978|504257111|3|0|1|504379733|1|0|1|500845639|2||-2||2|1|500011312, 500014681|500014681|-2|500014681|-2|0|5|||46|2|||1|942403|-1|4|3|44|0
94|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-10-30|NaT|Followup|2016-10-30|2016-10-27|Complete|Done|2|2|2|2|3|4|2.5|2|4|3|2|4|3|3|-16.67|4|2|3|2|2|3|2.67|2|3|4|4|3|3|3.17|-15.77|4|4|4|4|3|4|3|3.33|20.12|3|2|3|3|2.75|4|5|2|3|3.5|-21.43|4|4|4|4|4|4|3|3.86|4|3|2|2|3|4|4|3.14|22.93|4|4|3|3.67|3|4|2|3|22.33|4|4|4|3|3|3|33.33|2|2|2|2|0|4|4|4|4|0|Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016||16.3|Y|1|1|1|1|M|Hispanic||10|No|Mother|28212|3|One Parent: Female|$10,000 to $14,999|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28204|Masters Degree|Married|Consultant||0|9|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020753|504254978|504257111|3|0|1|504379733|1|0|1|500845639|2||-2||2|1|500011312, 500014681|500014681|-2|500014681|-2|0|5|||46|2|||1|953996|942403|4|3|45|0
97|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-11|NaT|Baseline|2015-10-13|2015-11-11|Complete|Done|4|1|4|1|3|4|2.83|||||||||2|3|4|4|3|4|3.33|||||||||4|4|4|4||||||1|1|1|1|1|||||||4|4|4|3|1|4|3|3.29||||||||||4|3|1|2.67||||||4|1|2.5|||||1|1||||4|4||||Green|||15.9||1|1|1|1|M|Black||10|Yes|Mother|28216|5|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community|Amachi|Match Support|M|Black||41|28214|Some College|Married|Business|28287|0|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504207638|504209750|31|0|1|504357457|31|0|1|500850393|2||-2||2|1||500000294|-2||-2|0|4|||17159|12|||1|944553|-1|4|3|44|7674215580094440446
97|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-11|NaT|Followup|2016-11-11|2017-01-26|Expired|Late||||||||4|1|4|1|3|4|2.83|||||||||2|3|4|4|3|4|3.33||||||4|4|4|4|||||||1|1|1|1|1||||||||||4|4|4|3|1|4|3|3.29||||||4|3|1|2.67|||||4|1|2.5||||1|1||||4|4||Green|||15.9||1|1|1|1|M|Black||10|Yes|Mother|28216|5|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community|Amachi|Match Support|M|Black||41|28214|Some College|Married|Business|28287|0|3|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504207638|504209750|31|0|1|504357457|31|0|1|500850393|2||-2||2|1||500000294|-2||-2|0|4|||17159|12|||1|959794|944553|4|0|45|7674215580094440446
98|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-11|NaT|Followup|2016-11-11|2016-11-22|Complete|Done|4|2|3|2||4||||||||||2|3|3|2|2|3|2.5|||||||||4|4|4|4||||||4|2|2|4|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|PERL 2014-2016||15.9||1|1|1|1|F|Black||10|No|Mother|28216|3|One Parent: Female|$15,000 to $19,999|Y|Yes||Self|General Community||Match Support|F|Hispanic||26|28031|Bachelors Degree|Single|Tech: Research/Design|28117|0|8|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500018851|504390954|504393193|31|0|2|504231700|3|0|2|500853984|2||-2||2|1|500014681||-2||-2|0|10|||17159|12|||1|962340||4|3|45|3650724132819756420
102|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-16|NaT|Followup|2016-11-16|2016-11-30|Complete|Done|3|3|3|2|3|3|2.83|4|4|4|1|4|4|3.5|-19.14|3|4|4|4|4|4|3.83|4|4|3|1|2|4|3|27.67|4|4|4|4|4|4|4|4|0|4|4|4|4|4|3|4|5|5|4.25|-5.88|4|4|4|4|4|4|4|4|4|4|4|4|4|4|2|3.71|7.82|4|4|4|4|3|4|4|3.67|8.99|4|4|4|3|1|2|100|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||15.8||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||33|28216|Bachelors Degree|Married|Business|28202|0|10|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504378557|1|0|1|500856483|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|961771|905704|4|3|45|3402014428779854546
104|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Baseline|2015-11-10|2015-11-17|Complete|Done|3|1|1|1|3|1|1.67|||||||||1|1|2|1|1|4|1.67|||||||||4|4|4|4||||||2|5|1|1|2.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016, Cabarrus County||15.7||1|1|1|1|M|White||15|Yes|Mother|28025|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28025|High School Graduate|Single|Business: Sales|28025|5|0|Local TV|Media|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821678|503823656|1|0|1|504468148|1|0|1|500858177|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7438|1|||1|959176|-1|4|3|44|7044657180546140448
104|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Followup|2016-11-17|2016-11-14|Complete|Done|4|4|1|1|1|4|2.5|3|1|1|1|3|1|1.67|49.7|4|4|4|4|4|4|4|1|1|2|1|1|4|1.67|139.52|2|4|4|3.33|4|4|4|4|-16.75|5|4|4|5|4.5|2|5|1|1|2.25|100|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|2|3.33|4|4|3|3.67|-9.26|2|4|3|4|4|4|-25|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016, Cabarrus County||15.7||1|1|1|1|M|White||15|Yes|Mother|28025|8|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||26|28025|High School Graduate|Single|Business: Sales|28025|5|0|Local TV|Media|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821678|503823656|1|0|1|504468148|1|0|1|500858177|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7438|1|||1|962415|959176|4|3|45|7044657180546140448
105|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Baseline|2015-11-10|2015-11-17|Complete|Done|3|1|1|1|1|1|1.33|||||||||1|3|4|2|1|4|2.5|||||||||1|1|1|1||||||4|3|5|2|3.5|||||||4|4|4|4|4|4|4|4||||||||||3|2|4|3||||||4|4|4|||||1|1||||4|4||||Green|PERL 2014-2016, Cabarrus County||15.7||1|1|1|1|M|White||12|Yes|Mother|28025|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||32|28025|Bachelors Degree||Business: Sales||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821686|503823656|1|0|1|504460050|1|0|1|500858397|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7496|10|||1|959399|-1|4|3|44|7044657180546140448
105|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-17|NaT|Followup|2016-11-17|2016-11-14|Complete|Done|1|1|4|1|1|4|2|3|1|1|1|1|1|1.33|50.38|2|2|4|2|2|4|2.67|1|3|4|2|1|4|2.5|6.8|2|2|4|2.67|1|1|1|1|167|5|4|5|5|4.75|4|3|5|2|3.5|35.71|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|3|4|3.67|3|2|4|3|22.33|3|2|2.5|4|4|4|-37.5|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016, Cabarrus County||15.7||1|1|1|1|M|White||12|Yes|Mother|28025|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||32|28025|Bachelors Degree||Business: Sales||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|503821686|503823656|1|0|1|504460050|1|0|1|500858397|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7496|10|||1|962429|959399|4|3|45|7044657180546140448
108|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-23|NaT|Baseline|2015-11-06|2015-11-23|Complete|Done|3|4|1|4|4|4|3.33|||||||||2|4|3|1|2|3|2.5|||||||||3|4|4|3.67||||||3|4|2|2|2.75|||||||4|4|4|4|4|4|2|3.71||||||||||3|3|3|3||||||4|4|4|||||2|2||||4|4||||Green|PERL 2014-2016||15.5||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28208|3|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||30|28204|Some College|Single|Medical|28208|3|3|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504278828|504281028|38|0|2|504354967|35|0|2|500857068|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|957729|-1|4|3|44|2378213070582218846
108|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-23|NaT|Followup|2016-11-23|2016-11-25|Complete|Done|4|4|4|4|4|4|4|3|4|1|4|4|4|3.33|20.12|2|4|4|3|3|4|3.33|2|4|3|1|2|3|2.5|33.2|4|4|4|4|3|4|4|3.67|8.99|4|3|3|4|3.5|3|4|2|2|2.75|27.27|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|2|3.71|4.04|4|4|4|4|3|3|3|3|33.33|4|3|3.5|4|4|4|-12.5|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||15.5||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28208|3|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Multi-race (Hispanic & White)||30|28204|Some College|Single|Medical|28208|3|3|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504278828|504281028|38|0|2|504354967|35|0|2|500857068|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|965373|957729|4|3|45|2378213070582218846
109|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-24|NaT|Baseline|2015-09-22|2015-11-24|Complete|Done|4|3|4|4|3|4|3.67|||||||||2|4|4|2|3|4|3.17|||||||||4|4|4|4||||||3|3|3|4|3.25|||||||4|4|4|4|2|4|3|3.57||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||15.5||1|1|1|1|M|Black||12|No|Mother|28211|5|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||48|28105||Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504227502|504229617|31|0|1|504460839|31|0|1|500859784|2||-2||2|1||500000294|-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1|936163|-1|4|3|44|2077565980961547475
109|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-24|NaT|Followup|2016-11-24|2016-12-27|Declined|Done||||||||4|3|4|4|3|4|3.67|||||||||2|4|4|2|3|4|3.17||||||4|4|4|4|||||||3|3|3|4|3.25||||||||||4|4|4|4|2|4|3|3.57||||||4|4|4|4|||||4|4|4||||2|2||||4|4||Green|||15.5||1|1|1|1|M|Black||12|No|Mother|28211|5|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||48|28105||Married|Retired||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504227502|504229617|31|0|1|504460839|31|0|1|500859784|2||-2||2|1||500000294|-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1|966066|936163|4|1|45|2077565980961547475
110|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-30|NaT|Baseline|2015-11-17|2015-11-30|Complete|Done|2|2|1|2|2|3|2|||||||||2|3|3|2|3|4|2.83|||||||||2|3|2|2.33||||||4|4|5|3|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|VOL - Mentoring Hispanic Youth, PERL 2014-2016||15.3||1|1|2|2|F|Hispanic||13|No|Mother|28205|6|Two Parent|Unknown||Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504331538|504333760|3|0|2|503843020|3|0|2|500860738|2||-2||2|2|500011312, 500014681|500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|962816|-1|4|3|44|0
110|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-11-30|NaT|Followup|2016-11-30|2016-11-29|Complete|Done|2|4|4|4|1|1|2.67|2|2|1|2|2|3|2|33.5|2|4|3|2|4|3|3|2|3|3|2|3|4|2.83|6.01|4|4|4|4|2|3|2|2.33|71.67|5|3|3|4|3.75|4|4|5|3|4|-6.25|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|4|0|4|4|4|4|4|4|4|4|0|2|4|3|4|4|4|-25|2|2|2|2|0|4|4|4|4|0|Yellow|VOL - Mentoring Hispanic Youth, PERL 2014-2016||15.3||1|1|2|2|F|Hispanic||13|No|Mother|28205|6|Two Parent|Unknown||Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504331538|504333760|3|0|2|503843020|3|0|2|500860738|2||-2||2|2|500011312, 500014681|500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|967639|962816|4|3|45|0
114|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-14|NaT|Baseline|2015-11-20|2015-12-14|Complete|Done|3|3|2|1|2|3|2.33|||||||||2|3|3|3|2|4|2.83|||||||||4|4|3|3.67||||||4|4|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||2|3|1|2||||||4|3|3.5|||||2|2||||4|4||||Green|Amachi, PERL 2014-2016||14.9||1|1|1|1|F|Black||15|Yes|Mother|28215|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi, PERL 2014-2016|Match Support|F|White||30|28203|Bachelors Degree|Single|Business|60611|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|503611732|503613600|31|0|2|504421910|1|0|2|500862006|2||-2||2|1|500000294, 500014681|500000294, 500014681|-2|500014681|-2|0|10|||17159|12|||1|964751|-1|4|3|44|0
114|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-14|NaT|Followup|2016-12-14|2016-12-12|Complete|Done|4|4|3|3|3|3|3.33|3|3|2|1|2|3|2.33|42.92|2|4|3|1|2|4|2.67|2|3|3|3|2|4|2.83|-5.65|4|2|2|2.67|4|4|3|3.67|-27.25|4|4|5|2|3.75|4|4|4|5|4.25|-11.76|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|3|3|2|2.67|2|3|1|2|33.5|2|2|2|4|3|3.5|-42.86|2|2|2|2|0|4|4|4|4|0|Green|Amachi, PERL 2014-2016||14.9||1|1|1|1|F|Black||15|Yes|Mother|28215|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community|Amachi, PERL 2014-2016|Match Support|F|White||30|28203|Bachelors Degree|Single|Business|60611|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|277|60|598|500000170|500020910|503611732|503613600|31|0|2|504421910|1|0|2|500862006|2||-2||2|1|500000294, 500014681|500000294, 500014681|-2|500014681|-2|0|10|||17159|12|||1|973924|964751|4|3|45|0
115|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-15|NaT|Baseline|2015-11-30|2015-12-15|Complete|Done|2|2|2|3|3|2|2.33|||||||||4|2|4|4|4|4|3.67|||||||||4|4|4|4||||||4|3|3|3|3.25|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||2|2|2|||||1|1||||4|4||||Green|PERL 2014-2016||14.8||1|1|1|1|F|Black||15|No|Mother|28215|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||26|28213|Bachelors Degree|Single|Business: Mgt, Admin|28105|2|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500021785|504393421|504395660|31|0|2|504395484|31|0|2|500863556|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||46|2|||1|967546|-1|4|3|44|5081726734274569781
115|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2015-12-15|NaT|Followup|2016-12-15|2017-03-01|Expired|Late||||||||2|2|2|3|3|2|2.33|||||||||4|2|4|4|4|4|3.67||||||4|4|4|4|||||||4|3|3|3|3.25||||||||||4|4|4|4|4|4|3|3.86||||||4|4|3|3.67|||||2|2|2||||1|1||||4|4||Green|PERL 2014-2016||14.8||1|1|1|1|F|Black||15|No|Mother|28215|9|One Parent: Female|Less than $10,000|Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|Black||26|28213|Bachelors Degree|Single|Business: Mgt, Admin|28105|2|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500021785|504393421|504395660|31|0|2|504395484|31|0|2|500863556|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|5|||46|2|||1|974242|967546|4|0|45|5081726734274569781
120|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-01-14|NaT|Baseline|2015-11-24|2016-01-14|Complete|Done|1|1|3|3|2|1|1.83|||||||||1|1|4|4|4|4|3|||||||||4|4|4|4||||||2|5|2|5|3.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||13.8||1|1|1|1|F|Black||10|No|Mother|28203|3|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||25|28209|Bachelors Degree|Single|Business|28277|1|0|Bowl For Kids Sake|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504388295|504390534|31|0|2|504404378|1|0|2|500870013|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||132|8|||1|966128|-1|4|3|44|2141487034287122220
120|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-01-14|NaT|Followup|2017-01-14|2017-02-20|Complete|Done|3|3|3|2|3|3|2.83|1|1|3|3|2|1|1.83|54.64|2|4|3|2|2|3|2.67|1|1|4|4|4|4|3|-11|4|4|4|4|4|4|4|4|0|3|4|3|3|3.25|2|5|2|5|3.5|-7.14|4|4|4|4|4|4|3|3.86|4|4|4|4|4|4|3|3.86|0|3|4|3|3.33|4|4|4|4|-16.75|2|3|2.5|4|3|3.5|-28.57|2|2|2|2|0|4|4|4|4|0|Green|PERL 2014-2016||13.8||1|1|1|1|F|Black||10|No|Mother|28203|3|One Parent: Female|Less than $10,000|Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||25|28209|Bachelors Degree|Single|Business|28277|1|0|Bowl For Kids Sake|Special Event|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504388295|504390534|31|0|2|504404378|1|0|2|500870013|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|34|2|||132|8|||1|982719|966128|4|3|45|2141487034287122220
130|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-12|NaT|Baseline|2016-01-29|2016-02-11|Complete|Done|3|3|3|1|3|3|2.67|||||||||2|4|4|2|4|3|3.17|||||||||2|4|4|3.33||||||3|3|2|5|3.25|||||||4|4|4|4|3|4|3|3.71||||||||||3|4|4|3.67||||||1|4|2.5|||||1|1||||4|4||||Green|PERL 2014-2016||12.9||1|1|1|1|M|Black||11|Yes|Mother|28215|5|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||29|28262|Some College|Single|Business|28204|0|4|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT, VOL - Thrive - Intro|Match Support|277|60|598|500000170|500020753|504230975|504233090|31|0|1|504284612|31|0|1|500876290|2||-2||2|1|500014681|500000294, 500014681|-2|500008492, 500011315, 500011316, 500014681|-2|0|4|||7462|13|||1|988696|-1|4|3|44|7327400833679234452
130|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-12|NaT|Followup|2017-02-12|2017-02-02|Complete|Done|3|2|3|3|1|2|2.33|3|3|3|1|3|3|2.67|-12.73|4|3|3|3|1|3|2.83|2|4|4|2|4|3|3.17|-10.73|4|4|4|4|2|4|4|3.33|20.12|4|3|5|4|4|3|3|2|5|3.25|23.08|4|4|4|4|4|4|4|4|4|4|4|4|3|4|3|3.71|7.82|2|4|2|2.67|3|4|4|3.67|-27.25|4|4|4|1|4|2.5|60|2|2|1|1|100|4|4|4|4|0|Green|PERL 2014-2016||12.9||1|1|1|1|M|Black||11|Yes|Mother|28215|5|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||29|28262|Some College|Single|Business|28204|0|4|Recruitment Event|BBBS Board/Staff|Big|General Community|PERL 2014-2016, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT, VOL - Thrive - Intro|Match Support|277|60|598|500000170|500020753|504230975|504233090|31|0|1|504284612|31|0|1|500876290|2||-2||2|1|500014681|500000294, 500014681|-2|500008492, 500011315, 500011316, 500014681|-2|0|4|||7462|13|||1|993665|988696|4|3|45|7327400833679234452
131|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-13|NaT|Baseline|2016-02-01|2016-02-13|Complete|Done|4|1|1|3|4|2|2.5|||||||||2|2|3|1|1|4|2.17|||||||||3|4|3|3.33||||||3|5|2|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|Cabarrus County||12.8||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28025|3|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||28|28027|Masters Degree|Single|Govt|28273|3|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504468562|504470835|36|0|1|504556956|31|0|1|500876668|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|989695|-1|4|3|44|7044657180546140448
131|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-13|NaT|Followup|2017-02-13|2017-02-28|Complete|Done|3|1|3|2|1|3|2.17|4|1|1|3|4|2|2.5|-13.2|3|4|3|2|4|3|3.17|2|2|3|1|1|4|2.17|46.08|4|4|4|4|3|4|3|3.33|20.12|4|3|5|2|3.5|3|5|2|5|3.75|-6.67|4|4|4|4|4|4|4|4|4|4|4|4|4|4|3|3.86|3.63|4|4|4|4|4|4|4|4|0|3|4|3.5|3|3|3|16.67|2|2|2|2|0|4|4|4|4|0|Green|Cabarrus County||12.8||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28025|3|One Parent: Female|$20,000 to $24,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|Black||28|28027|Masters Degree|Single|Govt|28273|3|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504468562|504470835|36|0|1|504556956|31|0|1|500876668|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|994031|989695|4|3|45|7044657180546140448
135|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-22|NaT|Baseline|2016-01-14|2016-02-22|Complete|Done|3|2|3|4|3|3|3|||||||||3|2|4|3|3|4|3.17|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||12.6||1|1|1|1|F|Multi-race (Black & White)||10|Yes|Foster Parent|28216|4|One Parent: Female|$40,000 to $44,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||45|28208|Bachelors Degree|Single|Education: Teacher|28208|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504498650|504500981|36|0|2|504131389|31|0|2|500878445|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|34|2|||46|2|||1|982537|-1|4|3|44|0
136|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-02-23|NaT|Baseline|2016-02-10|2016-02-23|Complete|Done|4|2|4|1|4|4|3.17|||||||||4|4|4|3|4|4|3.83|||||||||4|4|4|4||||||4|5|4|4|4.25|||||||4|4|4|4|3|4|3|3.71||||||||||4|4|4|4||||||4|3|3.5|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||12.5||1|1|1|1|M|Black||11|No|Mother|28262|3|One Parent: Female|$30,000 to $34,999||No|BBBS National Site|Web Link|General Community||Match Support|M|White||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|277|60|598|500000170|500017732|504295805|504298006|31|0|1|504337975|1|0|1|500878715|2||-2||2|1|500007920, 500011315, 500011316||-2||-2|34|2|||7464|9|||1|992976|-1|4|3|44|5923747279518652886
144|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-03-10|NaT|Baseline|2015-06-24|2016-03-08|Complete|Done|4|4|4|4|4|4|4|||||||||3|4|4|3|2|4|3.33|||||||||4|4|4|4||||||4|4|3|4|3.75|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|2|2.5|||||1|1||||4|4||||Green|PERL 2014-2016||12||1|1|1|1|M|Black||13|No|Mother|28208|6|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|White||26|28202|Bachelors Degree|Single|Law|28202|0|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504237243|504239358|31|0|1|504456306|1|0|1|500881682|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||17159|12|||1|909217|-1|4|3|44|7044657180546140448
146|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-03-14|NaT|Baseline|2016-02-29|2016-03-14|Complete|Done|4|2|2|1|3|3|2.5|||||||||3|4|4|2|2|4|3.17|||||||||4|4|4|4||||||3|4|5|4|4|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|1|1.5|||||2|2||||4|4||||Green|||11.9||1|1|1|1|F|Black||13|No|Mother|28278|6|One Parent: Female|$15,000 to $19,999|Y|Yes||School|General Community||Match Support|F|White||39|28134|Bachelors Degree|Single|Business: Marketing|28204|2|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504161470|504162947|31|0|2|504396335|1|0|2|500882097|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|999485|-1|4|3|44|2876415545463317777
148|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-03-23|NaT|Baseline|2016-03-09|2016-03-23|Complete|Done|4|4|1|2|1|4|2.67|||||||||2|1|3|4|1|3|2.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Yellow|Cabarrus County||11.6||1|1|1|1|M|Black||10|No|Mother|28027|3|One Parent: Female|$10,000 to $14,999|Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||35|28083|High School Graduate|Married|Medical||8|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504563369|504565703|31|0|1|504600175|1|0|1|500883737|2||500016307||2|2|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||46|2|||1|1002382|-1|4|3|44|6200244613298520712
152|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-06|NaT|Baseline|2016-03-30|2016-04-06|Complete|Done|1|4|4|4|4|3|3.33|||||||||2|4|2|2|3|4|2.83|||||||||4|4|4|4||||||5|3|3|4|3.75|||||||4|4|4|4|3|4|4|3.86||||||||||3|4|3|3.33||||||4|4|4|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||11.1||1|1|1|1|M|Black||12|No|Mother|28208|5|One Parent: Female|$30,000 to $34,999||Yes||Relative|General Community||Match Support|M|White||32|28203|Juris Doctorate (JD)|Single|Law: Lawyer|28277|1|6|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|503952082|503954090|31|0|1|504546069|1|0|1|500887070|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|0|3|||46|2|||1|1008663|-1|4|3|44|0
153|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-19|NaT|Baseline|2016-04-08|2016-04-19|Complete|Done|3|2|3|4|3|3|3|||||||||4|1|4|4|3|4|3.33|||||||||4|4|4|4||||||5|4|5|5|4.75|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|||10.7||1|1|1|1|M|White||11|No|Mother|28277|4|One Parent: Female|$75,000 to $99,999||No||School|General Community||Match Support|M|White||53|28270|Masters Degree|Married|Self-Employed, Entrepreneur||15|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504581060|504583394|1|0|1|504503934|1|0|1|500888341|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1|1011466|-1|4|3|44|5081726734274569781
157|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-24|NaT|Baseline|2016-03-28|2016-04-24|Complete|Done|2|2|2|1|2|3|2|||||||||2|2|3|3|2|3|2.5|||||||||4|4|4|4||||||4|4|4|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||1|2|1.5|||||2|2||||4|4||||Green|Cabarrus County, mentor2.0 2016||10.5||1|1|1|1|F|Black||13|No|Mother|28027|7|Two Parent|$60,000 to $74,999||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||30|28269|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|2|Recruitment Event|BBBS Board/Staff|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504602680|504605091|31|0|2|504579649|1|0|2|500886605|2||500016307||2|1|500016374, 500016394|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|4|||7462|13|||1|1007638|-1|4|3|44|993637920138474088
158|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-25|NaT|Baseline|2016-04-08|2016-04-25|Complete|Done|4|2|3|2|3|4|3|||||||||3|3|3|3|2|3|2.83|||||||||4|3|4|3.67||||||4|5|5|4|4.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|||10.5||1|1|1|1|M|White||11|No|Mother|28277|5|One Parent: Female|$60,000 to $74,999||No||School|General Community||Match Support|M|White||40|28173|Bachelors Degree|Married|Business: Mgt, Admin|33637|9|4|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500008321|504240231|504242346|1|0|1|504523981|1|0|1|500888425|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1011564|-1|4|3|44|7406803744350640674
160|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-04-28|NaT|Baseline|2016-04-07|2016-04-27|Complete|Done|3|4|4|4|4|4|3.83|||||||||2|3|3|3|2|2|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|3|3.86||||||||||3|3|3|3||||||2|3|2.5|||||1|1||||4|4||||Green|PERL 2014-2016, Cabarrus County||10.4||1|1|1|1|M|White||10|No|GrandMother|28124|3|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||35|28027|Bachelors Degree|Single|Tech: Computer/Programmer|28202|2|6|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, mentor2.0, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504640447|504638197|1|0|1|504266263|1|0|1|500888255|2||500016307||2|1|500014681, 500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500014505, 500016374|-2|0|4|||17159|12|||1|1011251|-1|4|3|44|0
165|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-10|NaT|Baseline|2016-05-02|2016-05-09|Complete|Done|3|4|4|4|4|4|3.83|||||||||3|3|3|3|3|3|3|||||||||4|4|4|4||||||3|3|4|3|3.25|||||||4|4|4|4|4|4|4|4||||||||||4|4|3|3.67||||||3|2|2.5|||||2|2||||4|4||||Green|PERL 2014-2016||10||1|1|3|3|M|Multi-race (Black & White)||12|Yes|Mother|28215|6|One Parent: Female|$35,000 to $39,999||No||School|General Community|Amachi, PERL 2014-2016|Match Support|M|Black||57|28269|Bachelors Degree|Married|Finance: Accountant|28202|34|2|Omega Psi Phi|Fraternity/Sorority|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|502183411|502183840|36|0|1|500189229|31|0|1|500891295|2||-2||2|1|500014681|500000294, 500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||8694|14|||1|1019351|-1|4|3|44|4203557099934965158
169|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-24|NaT|Baseline|2016-03-15|2016-05-24|Complete|Done|4|3|3|4|3|3|3.33|||||||||4|3|3|4|4|3|3.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||2|2||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||9.5||1|1|1|1|F|Black||10|No|Mother|28208|4|One Parent: Female|$20,000 to $24,999|Y|Yes||School|General Community||Match Support|F|White||29|28210|Bachelors Degree|Single|Business: Sales|28269|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020910|504556546|504558880|31|0|2|504283498|1|0|2|500889681|2||-2||2|1|500007920, 500011315, 500011316||-2||-2|0|4|||17159|12|||1|1004119|-1|4|3|44|6084148439133243542
171|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-31|NaT|Baseline|2016-05-16|2016-05-31|Complete|Done|2|2|4|2|3|1|2.33|||||||||4|2|2|4|4|4|3.33|||||||||4|4|4|4||||||3|5|4|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||3|4|3.5|||||2|2||||4|4||||Green|||9.3||1|1|1|1|F|Black||15|No|Mother|28212|8|One Parent: Female|$40,000 to $44,999||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||48|28212|Associate Degree|Single|Finance||11|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504473782|504476056|31|0|2|504550297|1|0|2|500893115|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||7464|9|||1|1025743|-1|4|3|44|2806833304218536184
172|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-05-31|NaT|Baseline|2016-05-13|2016-05-31|Complete|Done|2|4|4|4|4|2|3.33|||||||||3|4|4|3|4|4|3.67|||||||||4|4|4|4||||||4|5|4|1|3.5|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||9.3||1|1|1|1|M|Black||13|No|Mother|28227|7|One Parent: Female|$10,000 to $14,999|Y|Yes||School|General Community||Match Support|M|Black||27|28205|Some College|Single|Retail: Sales|28210|2|6|Local Radio|Media|Big|General Community||Match Support|277|60|598|500000170|500017732|504425160|504427415|31|0|1|504509415|31|0|1|500893007|2||-2||2|1|||-2||-2|0|4|||7437|1|||1|1024882|-1|4|3|44|5544164653861671456
177|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-14|NaT|Baseline|2016-06-14|2016-06-14|Complete|Done|3|3|1|2|2|4|2.5|||||||||3|3|4|3|3|3|3.17|||||||||4|3|4|3.67||||||2|5|5|4|4|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|Cabarrus County||8.8||1|1|1|1|F|White||11|No|GrandMother|28124|5|Grandparents|$10,000 to $14,999|Y|Yes||School|General Community|Cabarrus County|Match Support|F|White||45|28025|Some College||Business|28262|1|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504635786|504638197|1|0|2|504662207|1|0|2|500896660|2||500016307||2|1|500016374|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|1048528|-1|4|3|44|0
178|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-16|NaT|Baseline|2016-05-27|2016-06-16|Complete|Done|3|3|4|3|3|4|3.33|||||||||1|4|3|3|4|4|3.17|||||||||4|4|4|4||||||2|3|3|4|3|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||3|4|3.5|||||2|2||||4|4||||Green|PERL 2014-2016||8.8||1|1|1|1|F|Multi-Race (None of the above)||14|No|Mother|28215|7|One Parent: Female|Less than $10,000|Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Black||26|28262|Bachelors Degree|Single|Journalist/Media|28206|2|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504507791|504510086|7|0|2|504650231|31|0|2|500895078|2||-2||2|1|500014681|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|1034810|-1|4|3|44|7044657180546140448
179|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-16|NaT|Baseline|2016-05-24|2016-06-16|Complete|Done|4|4|1|4|3|4|3.33|||||||||2|4|3|1|2|3|2.5|||||||||4|4|4|4||||||5|5|5|5|5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||3|3|3|||||2|2||||4|4||||Green|||8.8||1|1|1|1|F|Black||11|No|Mother|28216|4|One Parent: Female|$20,000 to $24,999||Yes||Self|General Community||Match Support|F|White||27|28209|Bachelors Degree|Single|Medical|28054|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500017732|504628520|504630931|31|0|2|504409458|1|0|2|500894207|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|1031243|-1|4|3|44|7044657180546140448
180|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-20|NaT|Baseline|2016-05-23|2016-06-20|Complete|Done|3|2|3|2|2|3|2.5|||||||||3|2|3|4|3|2|2.83|||||||||4|4|4|4||||||4|5|3|5|4.25|||||||4|4|4|4|4|4|3|3.86||||||||||3|4||||||||3|3|3|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||8.6||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28213|7|One Parent: Female|$30,000 to $34,999|Y|Yes||Self|General Community||Match Support|M|Asian||25|28204|Bachelors Degree|Single|Finance|28215|0|6|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020752|504691840|504694268|36|0|1|504535890|4|0|1|500894068|2||-2||2|1|500007920, 500011315, 500011316||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1|1030379|-1|4|3|44|8773162532572605235
183|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-06-30|NaT|Baseline|2016-06-16|2016-06-30|Complete|Done|3|1|1|1|2|2|1.67|||||||||1|1|2|1|1|1|1.17|||||||||4|4|4|4||||||1|1|5|1|2|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||4|4|4|||||1|1||||4|4||||Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment||8.3||1|1|1|1|F|Black||12|No|Mother|28211|6|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||27|28205|Some College||Medical|28269|0|4|Current/Previous Big|Other Big|Big|General Community||Match Support|277|60|598|500000170|500020910|504471617|504473895|31|0|2|504458762|31|0|2|500897003|2||-2||2|1|500007920, 500011315, 500011316||-2||-2|0|10|||17159|12|||1|1049879|-1|4|3|44|1545381051186164660
260|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-28|NaT|Baseline|2016-11-11|2016-11-22|Complete|Done|3|2|3|2|2|3|2.5|||||||||4|4|4|2|4|3|3.5|||||||||4|4|4|4||||||5|4|4|5|4.5|||||||4|4|4|4|4|4|3|3.86||||||||||4|4|4|4||||||2|2|2|||||1|1||||4|4||||Green|||3.4||1|1|1|1|M|White||13|No|Mother|28277|8|One Parent: Female|$60,000 to $74,999||No||Self|General Community|PERL 2014-2016|Match Support|M|White||26|28207|Masters Degree|Living w/ Significant Other|Tech: Engineer|28203|1|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504808434|504810913|1|0|1|504557160|1|0|1|500926948|2||-2||2|1||500014681|-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|1103507|-1|4|3|44|5571803589598086587
261|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-29|NaT|Baseline|2016-09-16|2016-11-29|Complete|Done|3|2|1|1|2|2|1.83|||||||||2|3|2|2|2|2|2.17|||||||||3|3|3|3||||||1|2|4|5|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||1|3|2|||||1|1||||4|4||||Green|||3.3||1|1|1|1|F|Black||15|No|Mother|28211|9|One Parent: Female|Less than $10,000|Y|Yes||Self|General Community||Match Support|F|Black||47|28215|Masters Degree|Married|Education|28202|5|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504471621|504473895|31|0|2|504580592|31|0|2|500925801|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|1078193|-1|4|3|44|1545381051186164660
262|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-29|NaT|Baseline|2016-10-24|2016-11-29|Complete|Done|3|2|3|2|1|4|2.5|||||||||3|3|3|2|2|3|2.67|||||||||4|4|4|4||||||3|4|1|4|3|||||||4|4|4|4|3|4|2|3.57||||||||||4|4|4|4||||||3|3|3|||||1|1||||4|4||||Green|||3.3||1|1|1|1|F|Black||11|No|Mother|28209|5|One Parent: Female|$25,000 to $29,999||Yes||Self|General Community||Match Support|F|White||23|28203|Bachelors Degree||Finance: Accountant|28031|0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500018851|504662612|504665039|31|0|2|504595097|1|0|2|500918825|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1093147|-1|4|3|44|2719955880210213907
263|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-11-30|NaT|Baseline|2016-10-20|2016-11-10|Complete|Done|3|1|1|1|1|1|1.33|||||||||1|3|1|||||||||||||4|4|4|4||||||2|1|5|4|3|||||||4|4|4|4|4|4|4|4||||||||||3|3|3|3||||||4|4|4||||||||||4|4||||Green|||3.3||1|1|1|1|F|White||12|Yes|Non-Relative: Other|28205|5|One Parent: Female|$25,000 to $29,999|Y|Yes||Self|General Community||Match Support|F|White||28|28202|Bachelors Degree|Single|Finance|28202|5|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020753|504539986|504538455|1|0|2|504793129|1|0|2|500926111|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|1092039|-1|4|3|44|2082620892288628337
264|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-04|NaT|Baseline|2016-11-22|2016-12-04|Complete|Done|3|3|3|3|3|2|2.83|||||||||2|3|2|2|3|2|2.33|||||||||4|3|3|3.33||||||3|3|4|5|3.75|||||||4|4|4|4|4|4|3|3.86||||||||||3|4|3|3.33||||||1|4|2.5|||||2|2||||4|4||||Green|Cabarrus County||3.2||1|1|1|1|F|Black||12|No|Mother|28027|7|One Parent: Female|$15,000 to $19,999||Yes||School|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||24|28262|Masters Degree|Single|Human Services: Social Worker|28027|0|1|BBBS National Site|Web Link|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500022817|504937152|504939686|31|0|2|504797758|31|0|2|500930335|2||500016307||2|1|500016374|500014681, 500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||46|2|||1|1108671|-1|4|3|44|0
267|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-06|NaT|Baseline|2016-11-11|2016-12-06|Complete|Done|4|4|4|2|4|4|3.67|||||||||2|4|3|3|4|4|3.33|||||||||4|3|3|3.33||||||5|3|3|3|3.5|||||||4|4|4|4|4|4|2|3.71||||||||||4|4|4|4||||||2|4|3|||||2|2||||4|4||||Green|||3.1||1|1|1|1|M|Black||12|No|Mother|28213|5|One Parent: Female|$20,000 to $24,999|Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||33|28203|Bachelors Degree|Married|Business|32207|9|0|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|502383218|502383656|31|0|1|504867282|1|0|1|500926962|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|6854|8|||46|2|||1|1103521|-1|4|3|44|20998188998147742
271|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-21|NaT|Baseline|2016-09-16|2016-12-19|Declined|Done||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||Green|||2.6||1|1|1|1|M|Black||15|No|Mother|28227|8|One Parent: Female|$25,000 to $29,999|Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||25|28277|Bachelors Degree|Single|Business|28208|1|8|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504662357|504664784|31|0|1|504791469|31|0|1|500933117|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|34|2|||17159|12|||1|1078180|-1|4|1|44|3557919386369667257
272|BBBS of Greater Charlotte|Default|BBBS of Greater Charlotte|Main Office|C|Active|2016-12-21|NaT|Baseline|2016-10-21|2016-12-21|Complete|Done|4|1|1|1|4|4|2.5|||||||||1|4|4|1|1|4|2.5|||||||||4|4|4|4||||||3|3|3|3|3|||||||4|4|4|4|4|4|4|4||||||||||4|4|4|4||||||3|3|3||||||||||4|4||||Green|||2.6||1|1|1|1|M|Black||12|No|Mother|28210|5|One Parent: Female|$25,000 to $29,999|Y|Yes||School|General Community||Match Support|M|Black||30|28210|Bachelors Degree|Married|Military||1|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|277|60|598|500000170|500020910|504565095|504567429|31|0|1|504860995|31|0|1|500932205|2||-2||2|1|||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|1092382|-1|4|3|44|6156547733130613405
