ChildPartKey|VolPartKey|MatchKey|OfficeName|TeamName|Hybrid|MatchType|MatchStatus|QueueDescription|TimeInQueue|MatchSupportLevel|MatchReportSources|PendingMatchDate|MatchOpenDate|MatchCloseDate|MatchClosureReasons|MatchClosurePrimaryReason|MatchClosureSecondaryReason|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildLivingSituation|ChildIncomeLevel|MilitaryParent|ParentDeployed|ChildFamilyAssistance|ChildFreeReducedlunch|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|Beg|Open|Close|End|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|QueueKey|MatchTypeKey|MatchActivityKey|MatchSiteKey|StatusKey|MatchSupportLevelKey|ChildReportSourcesKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|MatchReportSourcesKey
500186464|500189376|500037414|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4088|Green||1997-11-04|1997-11-04|2009-01-13|Strong Relationship: Support No Longer Needed|Strong Relationship: Support No Longer Needed||134.3||1|1|2|2|F|Black||26||Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||60|28269|Bachelors Degree|Married|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500188181|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186029|500188979|500036979|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3564|Green||1999-04-22|1999-04-22|2009-01-23|Strong Relationship: Support No Longer Needed|Strong Relationship: Support No Longer Needed||117.1||1|1|1|1|M|Black||26||Mother|28208|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|Black||54|28105|Bachelors Degree|Married|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187816|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500186349|500189349|500037384|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1925|Green||2004-07-07|2004-07-07|2009-10-14|Child: Graduated|Child: Graduated||63.2||1|1|2|2|M|Black||26||Mother|28208|One Parent: Female|Unknown|||Y|No||Neighbor/Friend|General Community||Match Support|M|White||45|28211|Bachelors Degree|Single|Finance: Economist||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500187958|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
500186030|500188980|500036980|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3186|Green||2000-05-04|2000-05-04|2009-01-23|Strong Relationship: Support No Longer Needed|Strong Relationship: Support No Longer Needed||104.7||1|1|1|1|M|Black||26||Mother|28216|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|White||42|29601||Single|Business: Engineer||0|0||Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187883|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||0|10|||1|
500376900|500376909|500083705|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1104|Green||2006-03-03|2006-03-03|2009-03-11|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||36.3||1|1|3|3|M|White||26|No|Mother|28217|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||53|28226||Married|Business: Marketing||0|0|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187797|1|0|1|1|0|1|10|2|-2||4|1||-2||-1|0|10|||7464|9|||1|
500186729|500750594|500159730|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|752|Green|Amachi|2007-02-12|2007-02-12|2009-03-05|Vol: Other Reason|Vol: Other Reason||24.7||1|1|1|1|F|Black||25|Yes|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||39|28269||Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188072|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500185930|500188909|500036909|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1492|Green||2005-08-15|2005-08-15|2009-09-15|Child: Graduated|Child: Graduated||49||1|1|1|1|F|Black||25||Mother|28212|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|Black||36|28027|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187520|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500185666|500188616|500036616|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3165|Red||2001-01-02|2001-01-02|2009-09-02|Child: Graduated|Child: Graduated||104||1|1|1|1|M|Black||25||Mother|28203|One Parent: Female|Unknown|||Y|No|Brochure|Media|General Community||Match Support|M|Black||41|28216|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500187312|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|51|1|||7464|9|||1|
500186575|500189451|500037508|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3043|Green||2001-06-27|2001-06-27|2009-10-26|Child: Graduated|Child: Graduated||100||1|1|1|1|F|Black||25||Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||45|28214|Bachelors Degree|Single|Finance: Banking||0|0|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500188004|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7458|9|||1|
500186688|500189748|500037863|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1940|Green|Amachi|2004-06-16|2004-06-16|2009-10-08|Child: Graduated|Child: Graduated||63.7||1|1|1|1|F|Black||25|Yes|Mother|28215|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||45|28269|||Finance: Banking|28202|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188155|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500186318|500189327|500037347|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2337|Red||2002-10-11|2002-10-11|2009-03-05|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||76.8||1|1|1|1|F|Black||25||Mother|28208|Other/Unknown|Unknown||||No||School|General Community||Match Support|F|Asian||39|28205|Some College||Medical: Healthcare Worker||0|0||Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500187946|31|0|2|4|0|2|10|2|-2||4|3||-2||-2|0|4|||0|9|||1|
500185688|500188604|500036604|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2841|Green||2002-10-22|2002-10-22|2010-08-02|Child: Graduated|Child: Graduated||93.3||1|1|1|1|M|White||25||Mother|28217|Two Parent|Unknown||||No||School|General Community||Match Support|M|White||78|28277||Divorced|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500187321|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
500185702|500188653|500036653|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3543|Green||2000-03-02|2000-03-02|2009-11-13|Child: Graduated|Child: Graduated||116.4||1|1|1|1|M|White||25||Mother|28120|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||43|28146|Some College|Married|Insurance|28202|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187490|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500186678|500188441|500050852|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1741|Green|Amachi|2005-11-01|2005-10-27|2010-08-03|Child: Graduated|Child: Graduated||57.2||2|2|1|1|F|Black||25|Yes|Mother|28269|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||32|28273||Single|Student: College||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188055|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|6854|8|||2238|7|||1|500000294
500185700|500188695|500036695|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2199|Green||2003-09-29|2003-09-29|2009-10-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||72.2||1|1|1|1|F|Black||25||Mother|28208|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||36|28277|Some College|Single|Unknown||0|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008629|500187327|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500636686|500569051|500142359|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1192|Green||2006-11-21|2006-11-21|2010-02-25|Volunteer: Time constraint|Volunteer: Time constraint||39.2||1|1|2|2|M|Black||25||Mother|28205|One Parent: Female|$25,000 to $29,999|||Y|No||School|General Community||Match Support|M|Black||34|28205|Bachelors Degree|Single|Tech: Research/Design||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500636946|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|4|||46|2|||1|
500186040|500188989|500036989|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3102|Green||2002-12-19|2002-12-19|2011-06-17|Child: Graduated|Child: Graduated||101.9||1|1|1|1|F|Black||24|No|GrandMother|28208|Grandparents|Unknown||||No||Self|General Community||Match Support|F|Black||48|28217|Bachelors Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500187836|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500764771|500189381|500170997|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1099|Green||2007-04-05|2007-04-05|2010-04-08|Child: Graduated|Child: Graduated||36.1||1|1|3|3|F|Black||24||Mother|28212|Two Parent|Unknown||||No||Self|General Community||Match Support|F|Black||56|28269|Bachelors Degree|Divorced|Arts, Entertainment, Sports||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500765039|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500815555|500842415|500176537|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1051|Red||2007-05-11|2007-05-21|2010-04-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.5||1|1|1|1|F|Black||24|No|Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||35|28216||Single|Finance: Accountant||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500815824|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|34|2|||46|2|||1|
500754629|500789803|500162386|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|736|Green||2007-02-22|2007-03-21|2009-03-26|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||24.2||1|1|1|1|M|White||24|No|Mother|28124||Unknown||||No||Self|General Community||Match Support|M|White||30|28025|Some College|Single|Transport: Mechanic|28075|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|500754897|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500185675|500188632|500036632|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2617|Green||2003-06-04|2003-06-04|2010-08-03|Child: Graduated|Child: Graduated||86||1|1|1|1|F|Black||24||Mother|28262|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||43|28278|Juris Doctorate (JD)|Single|Law: Lawyer|28205|0|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187557|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7459|10|||1|
500186507|500189413|500037454|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3364|Green||2003-11-12|2001-05-18|2010-08-03|Child: Graduated|Child: Graduated||110.5||1|1|1|1|M|Black||24||Mother|28205|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||46|28269|Masters Degree|Married|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500188167|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||7496|10|||1|
500806676|500878893|500181682|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1219|Yellow||2007-06-20|2007-06-25|2010-10-26|Child: Graduated|Child: Graduated||40||1|1|1|1|M|Black||24||Mother|28269|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Match Support|M|Black||39|28213|Some College|Single|Military|28213|13|0|Radio|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500806944|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||131|1|||1|
500186436|500189444|500037500|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2654|Green||2003-08-07|2003-08-07|2010-11-12|Child: Graduated|Child: Graduated||87.2||1|1|1|1|M|Black||24||Mother|28216|One Parent: Female|Unknown||||No|Brochure|Media|General Community||Match Support|M|Black||42|28213|Bachelors Degree|Married|Finance: Banking||0|0|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187988|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|51|1|||7458|9|||1|
500185758|500188703|500036703|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3882|Green||2000-10-30|2000-10-30|2011-06-17|Child: Graduated|Child: Graduated||127.5||1|1|1|1|F|Black||24||Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||46|28078|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500187350|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500867574|500775714|500184661|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|730|Green|Amachi|2007-07-17|2007-07-30|2009-07-29|Volunteer: Moved|Volunteer: Moved||24||1|1|1|1|M|Black||24|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|No||Faith Organization|General Community|Amachi|Match Support|M|White||34|28209|Bachelors Degree|Single|Business: Sales|28216|1|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500867843|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
500186222|500189174|500037174|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1422|Red||2005-03-14|2005-03-14|2009-02-03|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||46.7||1|1|1|1|M|Some Other Race||24||Mother|28208|Other/Unknown|Unknown||||No||Self|General Community||Match Support|M|Black||41|28078||Single|Business: Marketing||0|0||Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187886|41|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||0|9|||1|
500344284|500336791|500129982|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|867|Green|Amachi|2006-10-12|2006-10-20|2009-03-05||||28.5||1|1|2|2|M|Black||24|Yes|Mother|28205|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||52|28216|Bachelors Degree|Married|Clergy|28216|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500344425|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500186788|500189605|500037707|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2460|Green||2004-09-21|2004-09-21|2011-06-17|Child: Graduated|Child: Graduated||80.8||1|1|2|2|M|Black||24||Mother|28208|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||47|28204||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500188098|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|6854|8|||7496|10|||1|
500186331|500189281|500037291|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3905|Green||2000-04-12|2000-04-12|2010-12-21|Child: Graduated|Child: Graduated||128.3||1|1|2|2|M|Black||24||Mother|28216|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187969|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
500186332|500189281|500037292|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2871|Green||2003-02-14|2003-02-10|2010-12-21|Child: Graduated|Child: Graduated||94.3||1|1|2|2|M|Black||24||Mother|28216|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187969|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
500186775|500189599|500037701|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2038|Yellow|Amachi|2004-08-30|2004-08-30|2010-03-30|Volunteer: Time constraint|Volunteer: Time constraint||67||1|1|1|1|M|Black||24|Yes|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||59|28216|Bachelors Degree|Widowed|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001281|500188088|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500767205|500868727|500179032|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|590|Yellow||2007-06-04|2007-06-12|2009-01-22|Child/Family: Moved|Child/Family: Moved||19.4||1|1|4|4|F|Black||24||Mother|28216|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|Black||38|28214|Bachelors Degree|Single|Business: Clerical|28273|2|3|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500001281|500767473|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500185939|500188874|500036874|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1452|Green||2005-02-11|2005-02-11|2009-02-02|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||47.7||1|1|2|2|M|Black||24||Mother|28025|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|Black||41|28027|Some College|Married|Law: Police Officer||5|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|500187530|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500185819|500188758|500036758|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1733|Green||2004-05-06|2004-05-06|2009-02-02|Child (or Parent): Other Reason|Child (or Parent): Other Reason||56.9||1|1|2|2|M|Black||24||Mother|28205|Other/Unknown|Unknown||||No||Self|General Community||Match Support|M|White||40|28205||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500187407|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500402676|500339569|500102368|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2073|Yellow|Amachi|2006-06-27|2006-06-27|2012-02-29|Child: Graduated|Child: Graduated||68.1||1|1|1|1|M|White||24|||28211|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community|Amachi|Match Support|M|White||36|28208|Bachelors Degree|Single|Business: Mgt, Admin|28203|2|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500402926|1|0|1|1|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|5|||2238|7|||1|500000294
500993537|500940949|500200304|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|442|Red||2007-10-02|2007-11-14|2009-01-29|Child/Family: Feels incompatible with volunteer Volunteer: Feels incompatible with child/family|Child/Family: Feels incompatible with volunteer|Volunteer: Feels incompatible with child/family|14.5||1|1|1|1|F|Black||24|No|Father|28104|One Parent: Male|$50,000 to $59,999||||No|BBBS National Site|Web Link|General Community||Match Support|F|Black||38|28269||Single|Customer Service||1|0|BBBS National Site|Web Link|Big|General Community||RTBM|1|0|1|0|277|60|598|500000170|500001267|500993810|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|34|2|||46|2|||1|
500186336|500189301|500037314|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3233|Green||2002-09-20|2002-09-20|2011-07-28|Child: Graduated|Child: Graduated||106.2||1|1|1|1|M|Black||24||Mother|28208|One Parent: Female|Unknown|||Y|No||School|General Community||Match Support|M|White||57|28277|Bachelors Degree|Married|Business: Sales||0|0|Billboard|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011184|500187974|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||125|1|||1|
500761777|500776552|500185821|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|560|Green||2007-07-24|2007-08-27|2009-03-09|Volunteer: Moved|Volunteer: Moved||18.4||1|1|2|2|M|Black||24||Mother|28215|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|Black||32|28202|Bachelors Degree|Single|Finance: Banking||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500762045|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500378573|500923396|500184849|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1135|Green|Amachi|2007-07-18|2007-08-14|2010-09-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||37.3||2|2|1|1|M|Black||24|Yes|Mother|28217|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||47|28213|Associate Degree|Single|Education: Teacher||4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500378823|31|0|1|31|0|1|10|2|-2||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500540838|501077532|500250641|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1028|Green|Amachi|2008-03-06|2008-03-07|2010-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||33.8||2|2|1|1|M|Black||23|Yes|Mother|28208|One Parent: Female|Unknown||||No||Service Organization|General Community|Amachi|Match Support|M|Black||39|28210|Bachelors Degree|Single|Business: Clerical||4|0|AA Task Force|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500541089|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|11|||6247|12|||1|500000294
500186291|500189241|500037241|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2432|Green||2004-11-30|2004-11-30|2011-07-29|Child: Graduated|Child: Graduated||79.9||1|1|2|2|F|Black||23||Foster Parent|28269|Other Relative|Unknown|||Y|No||Self|General Community||Match Support|F|Black||49|28269|Bachelors Degree|Divorced|Finance|28282|0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008629|500219859|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500342076|500188562|500080816|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2205|Green||2006-02-14|2006-02-14|2012-02-28|Child: Graduated|Child: Graduated||72.4||1|1|1|1|M|Black||23||Mother|28216|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|White||35|28207|Bachelors Degree|Single|Business: Marketing||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500342211|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1|
500870996|500869085|500176243|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1589|Green||2007-05-09|2007-05-16|2011-09-21|Child: Graduated|Child: Graduated||52.2||1|1|1|1|M|Black||23|No|Mother|28208|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|M|White||41|28209|Bachelors Degree|Divorced|Business: Sales|28202|0|7|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500871265|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500825243|500872550|500179954|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1143|Yellow||2007-06-12|2007-07-09|2010-08-25|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||37.6||1|1|1|1|M|Black||23|No|Relative: Other|28262|Two Parent|$10,000 to $14,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||31|28262|Some College|Single|Student: College|28203|0|6|TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500010765|500825512|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|34|2|||130|1|||1|
501234601|501223094|500271822|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1527|Yellow||2008-06-10|2008-06-24|2012-08-29|Child: Graduated|Child: Graduated||50.2||1|1|2|2|F|Black||23|No|Mother|28215|Grandparents|Unknown||||No|TV|Media|General Community||Match Support|F|Black||48|28211|Bachelors Degree|Single|Consultant|28278|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|1|0|1|0|277|60|598|500000170|500008629|501234877|31|0|2|31|0|2|10|2|-2||4|2||-2|500014505, 500015184|-1|56|1|||7462|13|||1|
501299223|501158791|500273953|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|852|Red||2008-06-18|2008-06-26|2010-10-26|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||28||1|1|1|1|F|White||23|No|Father|28214|One Parent: Male|Unknown||||No||Therapist/Counselor|General Community||Match Support|F|White||35|28207|Associate Degree|Single|Business: Mgt, Admin|28217|2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501299501|1|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|5|||7464|9|||1|
500185706|500188657|500036657|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4011|Green||2000-07-28|2000-07-28|2011-07-22|Child: Graduated|Child: Graduated||131.8||1|1|1|1|M|White||23||Mother|28226|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||46|28078|Bachelors Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187480|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501000034|501184263|500277856|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|160|Red||2008-07-15|2008-07-29|2009-01-05|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||5.3||1|1|1|1|M|Black||23|No|Mother|28262|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community||Match Support|M|Black||50|28213|Bachelors Degree|Married|Finance: Banking||3|0|AA Task Force|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|501000307|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|5|||6247|12|||1|
500948379|500952605|500192958|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1330|Yellow||2007-08-28|2007-08-30|2011-04-21|Child: Lost interest|Child: Lost interest||43.7||1|1|1|1|M|Black||23|No|Mother|28214|One Parent: Female|$30,000 to $34,999||||Yes||Neighbor/Friend|General Community||Match Support|M|Black||48|28273||Married|Tech: Research/Design||0|0|General|Other Big|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500011639|500948655|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|8|||6450|12|||1|
500463808|500498479|500117634|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1540|Yellow||2006-08-09|2006-08-15|2010-11-02|Volunteer: Time constraint|Volunteer: Time constraint||50.6||1|1|1|1|M|Black||23||Mother|28269|One Parent: Female|$50,000 to $59,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28269|Juris Doctorate (JD)|Single|Law: Lawyer||0|8|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500464059|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|34|2|||6450|12|||1|
501098842|500967139|500247572|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1496|Green||2008-02-25|2008-02-25|2012-03-31|Child: Graduated|Child: Graduated||49.1||1|1|2|2|M|Black||23|No|Mother|28216|One Parent: Female|$25,000 to $29,999||||No||Neighbor/Friend|General Community||Match Support|M|Black||60|28269|Bachelors Degree|Married|Business: Sales|28079|9|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501099116|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||4748|14|||1|
500186088|500188966|500036966|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2945|Green||2003-10-03|2003-10-03|2011-10-26|Child: Graduated|Child: Graduated||96.8||1|1|1|1|M|Black||23|No|Mother|28203|Other/Unknown|Unknown||||No||School|General Community||Match Support|M|White||44|28210|Bachelors Degree|Single|Finance: Banking|28211|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500002335|500187606|31|0|1|1|0|1|10|2|-2||4|1||-2||-1|0|4|||7496|10|||1|
500795704|500723270|500154833|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1583|Green|Amachi|2007-01-25|2007-01-30|2011-06-01|Child: Lost interest|Child: Lost interest||52||1|1|1|1|F|Multi-Race (None of the above)||23|Yes|Mother|28081|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||42|28075||Single|Medical: Pharmacist|28025|7|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500002335|500766037|7|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500474840|500708340|500172756|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1084|Yellow||2007-04-18|2007-04-18|2010-04-06|Child: Lost interest|Child: Lost interest||35.6||2|2|1|1|F|Black||23|No|Mother|28214|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||59|28205||Single|Law: Security Officer||11|0|Recruitment Event|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500009007|500474735|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|34|2|||7458|9|||1|
500575861|501202981|500274108|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1060|Green||2008-06-19|2008-07-22|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||34.8||2|2|1|1|F|Black||23||Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|No||Neighbor/Friend|General Community||Match Support|F|White||37|28209|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500576113|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
501202342|501213387|500262140|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|522|Green|Amachi|2008-04-22|2008-05-05|2009-10-09|Volunteer: Moved|Volunteer: Moved||17.1||1|1|1|1|F|Multi-race (Black & White)||23|Yes|Mother|28226|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|Asian||38|28205|Bachelors Degree|Single|Tech: Computer/Programmer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501202616|36|0|2|4|0|2|10|2|500003586||4|1|500000294|-2||-2|0|5|||2238|7|||1|500000294
500465521|500542558|500118432|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2110|Green|Amachi|2006-08-18|2006-08-21|2012-05-31|Child: Graduated|Child: Graduated||69.3||1|1|1|1|F|Black||23|Yes|Mother|28262|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|F|White||42|28209|Masters Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500465757|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294
500548831|500189256|500140290|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1249|Green||2006-11-14|2006-11-14|2010-04-16|Child/Family: Time constraints|Child/Family: Time constraints||41||1|1|6|6|F|Black||23||Mother|28262|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|F|Black||38|28269|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Site|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500001281|500549079|31|0|2|31|0|2|10|2|-2||4|1||-2|500007920, 500011315, 500011316, 500016374|-1|0|10|||7464|9|1360|3|1|
500398859|500954503|500274760|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|303|Yellow||2008-06-24|2008-07-07|2009-05-06|Child (or Parent): Other Reason Volunteer: Lost contact with child/agency|Child (or Parent): Other Reason|Volunteer: Lost contact with child/agency|10||3|3|1|1|F|Black||23||Mother|28227|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community||Match Support|F|White||38|28211|||Business: Clerical||1|0|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008062|500399109|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|5|||46|2|||1|
500809082|500878459|500178590|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1747|Yellow||2007-05-30|2007-06-01|2012-03-13|Child: Graduated|Child: Graduated||57.4||1|1|1|1|M|Black||23||Mother|28210|One Parent: Female|$35,000 to $39,999||||No||Self|General Community||Match Support|M|White||34|28203|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||RTBM|1|0|1|0|277|60|598|500000170|500011746|500809351|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500871235|500932548|500186929|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|590|Green|Amachi|2007-08-02|2007-08-14|2009-03-26|Volunteer: Lost contact with child/agency Child/Family: Lost contact with volunteer/agency|Volunteer: Lost contact with child/agency|Child/Family: Lost contact with volunteer/agency|19.4||1|1|1|1|M|Black||23|Yes|Mother|28083|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||57|28025||Married|Landscaper/Groundskeeper||13|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500001262|500871502|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500705925|500908500|500182939|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1338|Yellow||2007-07-03|2007-07-23|2011-03-22|Child/Family: Moved|Child/Family: Moved||44||1|1|2|2|M|Black||23||Relative: Other|28269|Other Relative|$60,000 to $74,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|Black||48|28269||Divorced|Tech: Engineer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500706192|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|34|2|||7496|10|||1|
500357337|501211519|500317956|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|698|Green||2008-11-19|2008-11-21|2010-10-20|Child/Family: Moved|Child/Family: Moved||22.9||2|2|1|1|F|White||23||Mother|28215|One Parent: Female|Unknown||||No||Relative|General Community||Match Support|F|White||47|28105|||Medical: Admin|28204|0|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500002335|500187556|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
500185781|500188751|500244796|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1538|Red||2008-02-13|2008-02-13|2012-04-30|Child: Graduated|Child: Graduated||50.5||2|2|2|2|M|Black||23||Mother|28262|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||34|28105||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013709|500187370|31|0|1|1|0|1|10|2|||4|3||-2||-2|6854|8|||7464|9|||1|
501086305|500189590|500251964|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|460|Green|Amachi|2008-03-12|2008-03-20|2009-06-23|Child/Family: Moved|Child/Family: Moved||15.1||1|1|5|5|M|Black||23|Yes|Mother|28277|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Some Other Race||46|28134|Bachelors Degree|Separated|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501086579|31|0|1|41|0|1|10|2|500003586||4|1|500000294|-2||-2|34|2|||2238|7|||1|500000294
500867579|500577903|500195387|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2019|Green|Amachi|2007-09-13|2007-09-22|2013-04-02|Child: Graduated|Child: Graduated||66.3||1|1|1|1|M|Black||23|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|No||Faith Organization|General Community|Amachi|Match Support|M|Black||42|28269||Single|Finance: Banking||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500867843|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
500185644|500188593|500036593|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3384|Red||2002-03-12|2002-03-12|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||111.2||1|1|1|1|M|Black||23||Mother|28269|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||46|28213|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500187279|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|8|||7496|10|||1|
500186926|500189699|500037812|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2669|Green|Amachi|2004-08-30|2004-08-30|2011-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||87.7||1|1|1|1|M|Some Other Race||23|Yes|Mother|28213|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||60|28277|Bachelors Degree|Married|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188133|41|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
501200793|500965108|500270284|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|300|Green||2008-06-06|2008-07-11|2009-05-07|Child/Family: Time constraints|Child/Family: Time constraints||9.9||1|1|2|2|M|Multi-race (Black & White)||22|No|Mother|28277|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||41|28211|||Finance: Banking||0|1|BBBS National Site|Web Link|Big|General Community||RTBM|1|0|1|0|277|60|598|500000170|500001281|501201067|36|0|1|31|0|1|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
500185745|500188692|500036692|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2223|Yellow||2004-01-05|2004-01-05|2010-02-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||73||1|1|1|1|M|Black||22||Mother|28278|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|White||42|28209|Masters Degree|Married|Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187340|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|8|||7464|9|||1|
500393176|500415570|500101074|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2206|Green|Amachi|2006-06-08|2006-06-07|2012-06-21|Child: Graduated|Child: Graduated||72.5||1|1|1|1|F|Black||22||Relative: Other|28216|Other Relative|Unknown||||No||Relative|General Community|Amachi|Match Support|F|Black||35|28213||Single|Tech: Engineer||2|0|Bellafonte Presbyter|Faith Organization|Big|General Site|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500013781|500187361|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-1|0|3|||2238|7|||1|500000294
500185712|500188663|500036663|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3079|Green||2000-09-28|2000-09-28|2009-03-04|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||101.2||1|1|1|1|M|White||22|No|Mother|28212|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||53|28227||Married|Business: Clerical||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500187555|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500186925|500189697|500037810|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2491|Green|Amachi|2005-02-24|2005-02-24|2011-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||81.8||1|1|1|1|M|Black||22|Yes|Mother|28205|One Parent: Female|Unknown|||Y|No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||59|28269|Masters Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188151|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500414113|500846653|500179366|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|925|Green||2007-06-07|2007-06-07|2009-12-18|Volunteer: Moved|Volunteer: Moved||30.4||1|1|1|1|F|Black||22||Mother|28208|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Enrollment|F|White||33|28226|||Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500414363|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|8|||46|2|||1|
500732462|500878773|500184327|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1686|Green||2007-07-13|2007-07-18|2012-02-28|Child: Graduated|Child: Graduated||55.4||1|1|1|1|F|Black||22||Mother|28205|One Parent: Female|$30,000 to $34,999|||Y|No||School|General Community||Match Support|F|Black||40|28269|Masters Degree|Single|Education: Admin|28223|1|9|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500732729|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||7458|9|||1|
500186615|500403330|500093132|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1969|Green|Amachi|2006-05-09|2006-05-09|2011-09-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||64.7||2|2|1|1|F|Black||22||Mother|28278|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||39|28269|PHD|Single|Medical: Doctor, Provider||0|8|Other|BBBS Board/Staff|Big|General Site|Amachi, mentor2.0 2014|Enrollment|1|0|1|0|277|60|598|500000170|500008629|500188023|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2|500000294, 500014506|-1|0|10|||7671|13|||1|500000294
500432759|500415680|500099996|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1587|Yellow||2006-05-26|2006-05-26|2010-09-29|Volunteer: Time constraint|Volunteer: Time constraint||52.1||1|1|1|1|F|Black||22||Mother|28205|One Parent: Female|Unknown||||No||Faith Organization|General Community||Match Support|F|Black||37|28216|Bachelors Degree|Single|Human Services: Non-Profit|28205|2|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500433090|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|9|||7464|9|||1|
501078559|501262050|500279449|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1417|Green|Amachi|2008-07-25|2008-08-04|2012-06-21|Child: Graduated|Child: Graduated||46.6||1|1|1|1|M|Black||22|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||37|28269|Bachelors Degree|Single|Medical: Admin|19380|0|9||Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501078832|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||0|11|||1|500000294
501185625|501170831|500274914|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|512|Green||2008-06-25|2008-07-28|2009-12-22|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||16.8||1|1|1|1|F|Black||22|No|Mother|28208|One Parent: Female|$20,000 to $24,999||||Yes||Neighbor/Friend|General Community||Match Support|F|Black||39|28208|Masters Degree|Single|Human Services: Social Worker|28025|0|1|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500009242|501185899|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|8|||46|2|||1|
500185628|500190654|500117464|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2213|Red||2006-08-07|2006-08-09|2012-08-30|Child: Graduated|Child: Graduated||72.7||2|2|2|2|M|American Indian or Alaska Native||22||Mother|28031|Other/Unknown|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|White||51|28078|Bachelors Degree|Married|Business: Sales|28269|0|6|Igniting Breakfast|Special Event|Big|General Community|mentor2.0, mentor2.0 2015|RTBM|1|0|1|0|277|60|598|500000170|500008321|500187262|6|0|1|1|0|1|10|2|||4|3||-2|500014505, 500015184|-2|0|8|||17266|8|||1|
500892907|500188541|500268211|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1566|Red|Amachi|2008-05-22|2008-05-29|2012-09-11|Child: Graduated|Child: Graduated||51.4||1|1|3|3|F|Black||22|No|Mother|28216|One Parent: Female|Unknown||||No||Faith Organization|General Community|Amachi|Match Support|F|Hispanic||37|28203|Some College|Single|Education: Teacher|28217|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|500893173|31|0|2|3|0|2|10|2|-2||4|3|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
500892903|501189856|500268753|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1669|Yellow|Amachi|2008-05-28|2008-05-29|2012-12-23|Child: Graduated|Child: Graduated||54.8||1|1|1|1|F|Black||22|Yes|Mother|28216|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||36|28273|Juris Doctorate (JD)|Single|Law: Lawyer|28052|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|500893173|31|0|2|31|0|2|10|2|-2||4|2|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500186136|500188550|500043731|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1684|Red||2005-09-23|2005-09-23|2010-05-04|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||55.3||2|2|1|1|F|Black||22||GrandMother|28205|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||38|28016|Some College|Single|Finance: Banking||7|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500187727|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
500186004|500188958|500036958|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2594|Green||2003-02-22|2003-02-22|2010-03-31|Volunteer: Moved|Volunteer: Moved||85.2||1|1|1|1|M|Black||22||Mother|28217|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|White||39|28134|Bachelors Degree|Single|Arts, Entertainment, Sports||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500187639|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
500186949|501212924|500262563|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1114|Green|Amachi|2008-04-23|2008-05-05|2011-05-24|Child: Lost interest|Child: Lost interest||36.6||2|2|1|1|M|Black||22|Yes|Mother|28215|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||37|28213|Bachelors Degree|Single|Consultant||2|6|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500188131|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||2238|7|||1|500000294
501285486|501161038|500274153|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|512|Green||2008-06-19|2008-06-19|2009-11-13|Child/Family: Moved|Child/Family: Moved||16.8||1|1|1|1|M|Black||22|No|Mother|28227|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|M|White||41|28203|Bachelors Degree|Single|Business: Mgt, Admin|28202|4|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501285764|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
500186830|500189605|500037708|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2164|Green||2005-07-14|2005-07-14|2011-06-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||71.1||1|1|2|2|M|Black||22||Mother|28208|Other/Unknown|Unknown||||No||Self|General Community||Match Support|M|White||47|28204||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500188106|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501074353|501116955|500247181|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|971|Green|Amachi|2008-02-21|2008-02-22|2010-10-20|Volunteer: Moved|Volunteer: Moved||31.9||1|1|1|1|M|Black||22|Yes|GrandMother|28025|Grandparents|Unknown||||No||Faith Organization|General Community|Amachi|Match Support|M|White||40|28269|Some College|Married|Business: Mgt, Admin|28273|10|3|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500002335|501074618|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||7464|9|||1|500000294
500378578|501537034|500341556|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|794|Green|Amachi|2009-02-17|2009-02-23|2011-04-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||26.1||2|2|1|1|F|Black||22|Yes|Mother|28217|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||64|28212|Masters Degree|Divorced|Education: Admin|28216|0|0|Recruitment Event|College Partner|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|500378823|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2|500000294|-2|0|8|||7448|5|||1|500000294
500876742|500865849|500178866|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|612|Green|Amachi|2007-06-01|2007-06-01|2009-02-02|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||20.1||1|1|2|2|M|Black||22|Yes|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||55|28083||Single|Govt: Mgmt/Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001262|500876680|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500186962|500367387|500086009|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1491|Green|Amachi|2006-03-24|2006-03-24|2010-04-23|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||49||2|2|1|1|F|Black||22||Mother|28269|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Enrollment|F|Black||55|28269||Married|Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500010355|500188165|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500186054|500189004|500037004|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2494|Green||2003-11-24|2003-11-24|2010-09-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||81.9||1|1|1|1|F|Black||22||Non-Relative: Other|28277|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||58|28078|Bachelors Degree|Married|Unknown||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500187666|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500958312|501249632|500271938|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|368|Green|Amachi|2008-06-10|2008-07-17|2009-07-20|Volunteer: Moved|Volunteer: Moved||12.1||2|2|1|1|M|Black||22|Yes|Mother|28212|One Parent: Female|$40,000 to $44,999|||Y|No||Service Organization|General Community|Amachi|Enrollment|M|White||35|28205|Bachelors Degree|Single|Journalist/Media|28205|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|500958582|31|0|1|1|0|1|5|2|500003586||4|1|500000294|-2||-2|0|11|||7464|9|||1|500000294
501249455|501488627|500317964|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1366|Red||2008-11-19|2008-12-03|2012-08-30|Child: Graduated|Child: Graduated||44.9||1|1|1|1|M|Black||22|No|Mother|28269|One Parent: Female|Unknown||||Yes|Brochure|Media|General Community||Match Support|M|Black||36|28262|Masters Degree|Single|Finance: Banking||6|6|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008321|501249731|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|51|1|||7464|9|||1|
501409300|501287416|500346626|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|501|Yellow||2009-03-03|2009-03-09|2010-07-23|Volunteer: Moved|Volunteer: Moved||16.5||1|1|1|1|F|Black||22|No|Mother|28278|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||37|76054|PHD|Single|Medical: Doctor, Provider|28203|1|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|501409585|31|0|2|31|0|2|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1|
500186683|501240668|500266144|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|275|Green|Amachi|2008-05-14|2008-06-03|2009-03-05|Child/Family: Lost contact with volunteer/agency Volunteer: Lost contact with child/agency|Child/Family: Lost contact with volunteer/agency|Volunteer: Lost contact with child/agency|9||3|3|1|1|M|Black||22|Yes|Mother|28262|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|M|Black||50|28213|Some College|Married|Tech: Engineer|28025|4|7|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500188164|31|0|1|31|0|1|5|2|500003586||4|1|500000294|-2||-2|0|10|||2238|7|||1|500000294
500780323|500992707|500203090|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|630|Green||2007-10-11|2007-10-30|2009-07-21|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.7||1|1|1|1|M|Black||22||Mother|28105|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||37|28270|Bachelors Degree|Single|Business: Mgt, Admin||3|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500780591|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500185729|500188672|500223221|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1745|Green||2007-11-26|2007-11-26|2012-09-05|Child: Graduated|Child: Graduated||57.3||2|2|2|2|M|Black||22||Relative: Other|28208|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||35|2109||Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500187496|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501373971|501359582|500290822|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|221|Green|Amachi|2008-09-24|2008-10-02|2009-05-11|Child: Lost interest|Child: Lost interest||7.3||1|1|2|2|F|Black||22|Yes|Mother|28273|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|F|Black||34|28273|Masters Degree|Living w/ Significant Other|Consultant|28273|1|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501374245|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|3|||7464|9|||1|500000294
500186800|500189320|500037337|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2849|Green||2004-10-06|2004-10-06|2012-07-25|Child: Graduated|Child: Graduated||93.6||1|1|3|3|F|Black||22||Mother|28216|Other/Unknown|Unknown||||No||School|General Community||Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500012459|500188103|31|0|2|31|0|2|10|2|-2||4|1||-2|500016374|-2|0|4|||7464|9|||1|
500764773|501091276|500235607|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1258|Red||2008-01-04|2008-01-06|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||41.3||2|2|1|1|F|Black||22||Mother|28212|Two Parent|Unknown||||No||Self|General Community||Match Support|F|White||36|28205|Bachelors Degree|Single|Medical: Nurse||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500765039|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
500526569|500497534|500118230|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1012|Green|Amachi|2006-08-16|2006-09-14|2009-06-22|Child: Lost interest Child/Family: Lost contact with volunteer/agency|Child: Lost interest|Child/Family: Lost contact with volunteer/agency|33.2||1|1|1|1|F|Black||22||Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community|Amachi|Match Support|F|Black||52|28212|Bachelors Degree|Married|Finance: Banking|28202|8|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500003657|500526820|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|5|||2238|7|||1|500000294
500414909|500188447|500510533|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|565|Green|2010-2012 OJJDP JJI|2011-01-12|2011-01-12|2012-07-30|Child: Graduated|Child: Graduated||18.6||3|3|3|3|M|White||22|No|Mother|28027|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||56|28078|Bachelors Degree|Single|Business: Sales|28027|14|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500002335|500415159|1|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|0|10|||7446|3|||1|500005291
500414909|500188447|500173974|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1280|Green||2007-04-26|2007-04-26|2010-10-27|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||42.1||3|3|3|3|M|White||22|No|Mother|28027|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||56|28078|Bachelors Degree|Single|Business: Sales|28027|14|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500002335|500415159|1|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|0|10|||7446|3|||1|
500186047|501176920|500276662|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|298|Green||2008-07-07|2008-07-10|2009-05-04|Vol: Lost Interest|Vol: Lost Interest||9.8||3|3|1|1|F|Black||22||Mother|28206|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|White||31|28206|Bachelors Degree|Single|Finance: Banking||0|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500187662|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|8|||46|2|||1|
500234359|500251451|500068942|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2008|Red||2005-12-17|2005-12-17|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||66||1|1|1|1|M|Black||22||Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||33|28269|Bachelors Degree|Single|Finance: Banking|28262|2|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500234368|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500185678|500188619|500036619|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3446|Green||2003-02-23|2003-02-23|2012-07-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||113.2||1|1|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||42|28277|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500187309|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500916715|500871928|500183554|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|555|Green||2007-07-11|2007-07-11|2009-01-16|Child: Lost interest|Child: Lost interest||18.2||1|1|1|1|F|Black||22|No|Mother|28227|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|Black||47|28270|Masters Degree||Education||2|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008062|500916985|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186453|500189369|500037407|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2828|Green||2002-09-14|2001-09-18|2009-06-16|Volunteer: Moved Child (or Parent): Other Reason|Volunteer: Moved|Child (or Parent): Other Reason|92.9||1|1|1|1|M|Black||22||Non-Relative: Other|28205|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||50|28216|Bachelors Degree|Married|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500188176|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186813|500189600|500037702|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2389|Red||2004-10-05|2004-10-05|2011-04-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||78.5||1|1|2|2|M|Black||22||Mother|28273|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||46|28214|Bachelors Degree|Single|Finance: Economist|28217|14|0|Brochure|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500188094|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|8|||127|1|||1|
501459095|501508823|500335575|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|692|Yellow||2009-01-26|2009-01-28|2010-12-21|Volunteer: Moved|Volunteer: Moved||22.7||1|1|1|1|F|Black||22|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||31|28202|Bachelors Degree|Single|Retail: Sales|28226|0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501459380|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500186970|500189743|500037857|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1661|Green||2005-04-04|2005-04-04|2009-10-21|Child/Family: Moved|Child/Family: Moved||54.6||1|1|1|1|F|Hispanic||22||Mother|28215|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||36|28209|||Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500548897|3|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500824047|500923510|500193080|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|726|Green||2007-08-29|2007-09-05|2009-08-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||23.9||1|1|1|1|M|Black||22|No|Mother|28269|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||Enrollment|M|Some Other Race||40|28277|Masters Degree|Married|Human Services: Youth Worker|29730|7|9|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|500824306|31|0|1|41|0|1|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500186374|500419439|500102160|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2022|Yellow||2006-06-23|2006-06-28|2012-01-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||66.4||2|2|1|1|F|Black||22||Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||55|28269|High School Graduate|Single|Business: Human Resources|28202|5|0|AA Task Force|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500187968|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||6247|12|||1|
500186107|500392161|500102003|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2309|Green||2006-06-22|2006-06-22|2012-10-17|Child: Graduated|Child: Graduated||75.9||2|2|1|1|M|Black||22||Mother|28206|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|Black||52|28210|Masters Degree|Married|Business: Mgt, Admin||0|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500187654|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||2230|7|||1|
500186325|500189265|500047102|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3298|Green||2005-10-19|2003-11-19|2012-11-29|Child: Graduated|Child: Graduated||108.4||2|2|2|3|M|Black||22||Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||39|28202|Bachelors Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|500187951|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186924|500483618|500108918|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1057|Green|Amachi|2006-07-25|2006-07-31|2009-06-22|Child: Cust. Adult Unsupportive/Interfered|Child: Cust. Adult Unsupportive/Interfered||34.7||2|2|1|1|M|Black||22|Yes|Mother|28217|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|M|White||69|28203|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188132|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
501171388|501126269|500247001|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|456|Green||2008-02-21|2008-02-27|2009-05-28|Vol: Lost Interest Vol: Family Change|Vol: Lost Interest|Vol: Family Change|15||1|1|1|1|F|Black||22|No|Mother|28025|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||45|28075||Married|Business: Clerical||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|501171662|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|34|2|||7671|13|||1|
501030388|501169473|500290065|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|164|Red||2008-09-22|2008-12-15|2009-05-28|Volunteer: Moved|Volunteer: Moved||5.4||1|1|2|2|M|Black||22|No|Mother|28210|One Parent: Female|$40,000 to $44,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||42|28277|Bachelors Degree|Single|Business: Sales|28208|5|7|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|501030661|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
501099294|500897787|500244827|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1205|Yellow||2008-02-13|2008-02-28|2011-06-17|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||39.6||1|1|1|1|F|Black||22|No|Mother|28206|One Parent: Female|$15,000 to $19,999||||Yes||Neighbor/Friend|General Community||Match Support|F|White||40|28205|Bachelors Degree|Single|Business: Sales|28277|0|3|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501099568|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|8|||46|2|||1|
501457664|501728924|500368257|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|469|Green||2009-06-10|2009-06-17|2010-09-29|Volunteer: Moved|Volunteer: Moved||15.4||1|1|1|1|M|Black||22|No|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||36|28203||Single|Business: Marketing||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501457949|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
500185676|500192243|500046426|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1209|Yellow||2005-10-13|2005-10-13|2009-02-03|Child (or Parent): Other Reason Vol: Other Reason|Child (or Parent): Other Reason|Vol: Other Reason|39.7||2|2|1|1|M|Black||22||Mother|28215|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||35|28215||Single|Retail: Sales|28027|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187307|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|8|||46|2|||1|
500185535|500921223|500182913|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|714|Green||2007-07-03|2007-07-11|2009-06-24|Vol: Family Change|Vol: Family Change||23.5||1|1|1|1|F|Black||22||GrandMother|28208|Grandparents|Unknown|||Y|No||Neighbor/Friend|General Community||Match Support|F|Some Other Race||48|28216|||Medical: Nurse||0|0|Essence Magazine|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187160|31|0|2|41|0|2|10|2|-2||4|1||-2||-2|0|8|||3892|1|||1|
501184653|501216727|500256896|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|382|Green||2008-04-04|2008-04-04|2009-04-21|Vol: Other Reason|Vol: Other Reason||12.6||1|1|1|1|M|White||22|No|Mother|28081|One Parent: Female|Unknown||||No||Self|General Community||RTBM|M|White||39|28081||Married|Transport: Driver||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|501184919|1|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186327|500189289|500037301|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3611|Red||2003-01-11|2003-01-11|2012-11-30|Child: Graduated|Child: Graduated||118.6||1|1|1|1|M|Black||22||Mother|28208|One Parent: Female|Unknown|||Y|No||School|General Community||Match Support|M|White||63|28211|Some College|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008321|500187974|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
500187030|500189679|500037792|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2149|Green||2005-02-23|2005-02-23|2011-01-12|Child: Lost interest|Child: Lost interest||70.6||1|1|1|1|F|Hispanic||22|No|Mother|28027|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|White||50|28078|Bachelors Degree|Married|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500188205|3|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500726828|500863980|500173102|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1582|Green||2007-04-23|2007-05-14|2011-09-12|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||52||1|1|3|3|M|Black||22||Mother|28027|One Parent: Female|$40,000 to $44,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||49|28027|Bachelors Degree|Married|Transport: Driver|28208|6|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500002335|500187529|31|0|1|31|0|1|10|2|-2||4|1||-2|500014505, 500014506|-1|34|2|||7671|13|||1|
500185972|500492482|500120588|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2303|Green|Amachi|2006-09-01|2006-09-01|2012-12-21|Child: Graduated|Child: Graduated||75.7||2|3|1|1|F|Black||22|Yes|Mother|28206|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Match Support|F|Black||38|28213|Bachelors Degree|Single|Education: Teacher|28202|2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500187610|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501315399|500957632|500328684|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|298|Green||2008-12-22|2009-01-08|2009-11-02|Child/Family: Moved|Child/Family: Moved||9.8||1|1|2|2|F|Black||22|No|Mother|28269|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|F|Black||32|28209|Bachelors Degree||Finance: Banking||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501315677|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|8|||46|2|||1|
500872449|500846955|500178294|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2101|Red||2007-05-25|2007-05-30|2013-02-28|Volunteer: Time constraint|Volunteer: Time constraint||69||1|1|2|2|M|Black||22|No|Mother|28211|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Match Support|M|White||37|28209|Masters Degree|Single|Business: Marketing|28208|1|9|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500872718|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500697380|500752342|500168910|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1466|Yellow||2007-03-27|2007-04-16|2011-04-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||48.2||1|1|2|2|M|White||22||Mother|28105|One Parent: Female|$25,000 to $29,999||||Yes||Therapist/Counselor|General Community||Match Support|M|White||53|28227|||Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500697647|1|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|5|||46|2|||1|
500186473|500344294|500092470|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1638|Green|Amachi|2006-05-03|2006-05-02|2010-10-26|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||53.8||3|3|1|1|F|Black||22|Yes|Mother|28205|One Parent: Female|Unknown|||Y|No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||43|28215|Masters Degree|Single|Business: Engineer|28269|1|3|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500187991|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500186146|500191447|500049095|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1237|Green||2005-10-27|2005-10-27|2009-03-17|Child/Family: Lost contact with volunteer/agency Volunteer: Moved|Child/Family: Lost contact with volunteer/agency|Volunteer: Moved|40.6||2|2|1|1|M|Black||22||Mother|28213|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||42|28205|Masters Degree|Divorced|Business: Marketing||3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500187734|31|0|1|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500187077|500189823|500037943|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2863|Green||2005-05-31|2005-05-31|2013-04-02|Child: Graduated|Child: Graduated||94.1||2|2|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||43|28210|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500188224|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500187077|500189824|500037944|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2863|Green||2005-05-31|2005-05-31|2013-04-02|Child: Graduated|Child: Graduated||94.1||2|2|1|1|M|Black||22||Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||41|28210|Bachelors Degree|Married|Medical: Pharmacist||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500188224|31|0|1|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500736888|501355773|500309757|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|779|Green||2008-11-03|2008-11-11|2010-12-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||25.6||2|2|1|1|M|Black||22||Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|No||School|General Community||Match Support|M|White||31|28226|Bachelors Degree|Married|Finance: Banking|28255|6|0|Neighbor/Friend|Neighbor/Friend|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500008629|500737155|31|0|1|1|0|1|10|2|-2||4|1||-2|500014505, 500014506|-1|0|4|||7496|10|||1|
500488488|500226756|500108788|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1217|Yellow||2006-07-24|2006-07-27|2009-11-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||40||1|1|2|2|M|Black||22||Aunt|28217|Other Relative|Unknown|||Y|No||Neighbor/Friend|General Community||Match Support|M|Black||33|28207|Bachelors Degree|Single|Business: Sales||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500488739|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|8|||46|2|||1|
500186385|500189269|500037278|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3620|Green||2003-02-11|2003-02-11|2013-01-09|Child: Graduated|Child: Graduated||118.9||1|1|1|1|M|Black||22||Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||43|28269|Bachelors Degree|Single|Finance: Accountant|28262|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500004169|500187967|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500965126|501572572|500341377|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|568|Yellow||2009-02-16|2009-02-17|2010-09-08|Child/Family: Moved|Child/Family: Moved||18.7||2|2|1|1|M|White||22|No|Mother|28134|One Parent: Female|$45,000 to $49,999||||No||Therapist/Counselor|General Community||Match Support|M|White||31|28105|High School Graduate|Single|Retail: Mgt|28105|4|0||Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|500965396|1|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|5|||0|11|||1|
501097465|501012178|500236354|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1034|Green||2008-01-09|2008-01-25|2010-11-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34||1|1|1|1|F|White||22|No|Father|28027|One Parent: Male|Unknown||||Yes||School|General Community||Match Support|F|White||51|28075||Single|Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501097739|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||46|2|||1|
501234992|501009895|500265126|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|733|Red||2008-05-07|2008-05-21|2010-05-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.1||1|1|1|1|F|Black||22|No|Mother|28273|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||32|28273|Bachelors Degree|Single|Business: Sales|20190|0|4|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|501235268|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||6450|12|||1|
501002521|501363548|500294584|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|643|Yellow||2008-10-03|2008-12-04|2010-09-08|Volunteer: Time constraint|Volunteer: Time constraint||21.1||2|2|1|1|F|Black||22|No|Mother|28214|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|F|White||32|28209|Bachelors Degree|Single|Human Services: Non-Profit||1|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501002794|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501333719|501172171|500289665|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|567|Yellow|Amachi|2008-09-19|2008-09-26|2010-04-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.6||1|1|1|1|F|Black||22|Yes|Mother|28212|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||35|28262|Associate Degree|Single|Education: Teacher|28205|3|3|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501333998|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2||-2|0|8|||6450|12|||1|500000294
500577965|500458869|500127631|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1074|Green||2006-10-06|2006-10-10|2009-09-18|Child/Family: Moved|Child/Family: Moved||35.3||1|1|1|1|M|Black||22||Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|No||Neighbor/Friend|General Community||Match Support|M|White||40|28209|Bachelors Degree|Single|Business: Engineer|28217|1|0|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500001281|500578217|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|8|||46|2|||1|
500574639|500724574|500140736|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1399|Green||2006-11-15|2006-11-15|2010-09-14|Volunteer: Moved|Volunteer: Moved||46||1|1|1|1|M|Black||22||Aunt|28269|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|Black||32|28277||Single|Arts, Entertainment, Sports||1|6|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500574891|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7447|3|||1|
501114443|501180846|500290376|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1751|Green|Amachi|2008-09-23|2008-10-08|2013-07-25|Child: Graduated|Child: Graduated||57.5||1|1|2|2|M|Black||22|No|Uncle|28206|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||34|28205|Juris Doctorate (JD)|Married|Law: Lawyer||0|4|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501114708|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||46|2|||1|500000294
500402978|500414710|500103314|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2140|Yellow|Amachi|2006-06-29|2006-06-29|2012-05-08|Child/Family: Time constraints|Child/Family: Time constraints||70.3||1|1|1|1|M|White||22||Mother|28211|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||33|28203|Bachelors Degree|Single|Business: Sales|27609|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500402926|1|0|1|1|0|1|10|2|-2||4|2|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
501820715|501049119|500387870|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|403|Green||2009-09-24|2009-10-23|2010-11-30|Volunteer: Health|Volunteer: Health||13.2||1|1|2|2|M|Black||22|No|Mother|28227|One Parent: Female|Unknown|||Y|Yes||Relative|General Community||Match Support|M|Black||68|28212|Associate Degree|Married|Craftsman||25|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|501821070|31|0|1|31|0|1|10|2|-2||4|1||-2|500000294|-2|0|3|||2238|7|||1|
500764136|501915488|500428501|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|925|Green|Amachi|2010-01-20|2010-02-10|2012-08-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||30.4||3|3|1|1|M|Black||22|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community|Amachi|Match Support|M|White||32|28210|Some College|Single|Business: Mgt, Admin|28206|8|2|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|500764404|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
500764136|501377225|500320856|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|328|Green|Amachi|2008-11-26|2008-12-03|2009-10-27|Volunteer: Time constraint|Volunteer: Time constraint||10.8||3|3|1|1|M|Black||22|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Finance: Accountant|28202|0|1|other|College Partner|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500764404|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7670|5|||1|500000294
501630156|500188758|500344438|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|665|Green||2009-02-24|2009-02-24|2010-12-21|Child: Lost interest|Child: Lost interest||21.8||1|1|2|2|M|Black||22|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||40|28205||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|500187407|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500906209|500871224|500272050|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|348|Green||2008-06-11|2008-06-25|2009-06-08|Volunteer: Moved|Volunteer: Moved||11.4||1|1|1|1|F|Black||22|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Enrollment|F|White||39|28205|Bachelors Degree|Single|Service: Tourism|28255|3|10|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500008628|500906479|31|0|2|1|0|2|5|2|-2||4|1||-2||-1|0|10|||7464|9|||1|
501431901|501780241|500384909|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|654|Green||2009-09-15|2009-09-22|2011-07-08|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.5||1|1|1|1|M|Black||22|No|Mother|28083|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||48|28081||Single|Medical: Healthcare Worker||0|0|AA Task Force|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501432186|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||9226|6|||1|
500185596|500310736|500068627|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1963|Green||2005-12-15|2005-12-19|2011-05-05|Child: Lost interest|Child: Lost interest||64.5||1|1|1|1|M|Black||22||Mother|28205|Other/Unknown|Unknown||||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500187230|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500840811|501391123|500308254|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|251|Green|Amachi|2008-10-30|2008-11-07|2009-07-16|Child: Lost interest|Child: Lost interest||8.2||2|2|3|3|F|Black||22|Yes|Mother|28083|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|Black||41|28027|PHD|Single|Medical: Doctor, Provider|28075|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500001262|500408385|31|0|2|31|0|2|10|2|500003586||4|1||-2|500016374|-2|0|8|||7464|9|||1|500000294
500185721|500188678|500036678|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3096|Green||2003-12-03|2003-12-03|2012-05-25|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||101.7||1|1|1|1|M|Black||22||Mother|28054|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||43|28207||Single|Unknown||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187333|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500843860|501340550|500320896|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|837|Green|Amachi|2008-11-26|2008-12-14|2011-03-31|Volunteer: Moved|Volunteer: Moved||27.5||2|2|1|1|M|Black||22|Yes|Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|No|TV|Media|General Community||Match Support|M|White||33|28202|Bachelors Degree|Single|Finance: Banking|28255|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500844129|31|0|1|1|0|1|10|2|500003586||4|1||-2||-2|56|1|||46|2|||1|500000294
501310912|501348323|500286597|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|436|Green||2008-09-08|2008-09-29|2009-12-09|Volunteer: Moved|Volunteer: Moved||14.3||1|1|1|1|F|Black||21|No|Mother|28262|One Parent: Female|Unknown||||No||Relative|General Community||Match Support|F|White||34|28269|Masters Degree|Single|Medical: Healthcare Worker|27103|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501311190|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
500911245|500852314|500278884|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|719|Green|Amachi|2008-07-22|2008-08-07|2010-07-27|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||23.6||2|2|2|2|F|Black||21|Yes|Mother|28075|One Parent: Female|$15,000 to $19,999|||Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||53|28262|Bachelors Degree|Married|Medical: Nurse|28207|6|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500911515|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|9|||7464|9|||1|500000294
501457406|501720969|500375964|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1426|Green||2009-07-28|2009-08-20|2013-07-16|Child: Graduated|Child: Graduated||46.9||1|1|1|1|M|Black||21|No|Mother|28269|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28205|||Finance: Banking|28217|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|501457691|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|6854|8|||7464|9|||1|
501314431|501564923|500338142|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|386|Yellow||2009-02-03|2009-02-09|2010-03-02|Volunteer: Time constraint|Volunteer: Time constraint||12.7||1|1|1|1|M|Black||21||GrandMother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||54|28215|Some College|Divorced|Business: Human Resources|28269|23|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|500947529|31|0|1|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500186662|500189813|500037930|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1635|Yellow|Amachi|2005-08-11|2005-08-11|2010-02-01|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||53.7||2|2|2|2|F|Black||21||Mother|28278|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Enrollment|F|Black||39|28278|Bachelors Degree|Single|Finance: Accountant|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500188023|31|0|2|31|0|2|5|2|500003586||4|2|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500186247|500189197|500037197|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2645|Red||2005-06-30|2005-06-30|2012-09-26|Child: Graduated|Child: Graduated||86.9||1|1|2|2|M|Black||21||Mother|28213|Other/Unknown|Unknown||||No||Self|General Community||Match Support|M|Black||39|28269|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Site|mentor2.0 2014|RTBM|1|0|1|0|277|60|598|500000170|500008321|500187842|31|0|1|31|0|1|10|2|-2||4|3||-2|500014506|-1|0|10|||7464|9|||1|
500185815|501356152|500419960|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|615|Green||2009-12-09|2009-12-17|2011-08-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.2||5|5|2|2|F|Black||21|No|Mother|28213|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||44|28211|Bachelors Degree|Single|Transport: Flight Attendant||10|0|Other|Service Organization|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500001281|500187403|31|0|2|1|0|2|10|2|-2||4|1||-2||-1|0|10|||7452|6|||1|
500185815|500556707|500254150|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|587|Green||2008-03-25|2008-04-02|2009-11-10|Volunteer: Moved|Volunteer: Moved||19.3||5|5|2|2|F|Black||21|No|Mother|28213|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||35|28269||Single|Child/Day Care Worker|28012|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500187403|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500544934|501213248|500269480|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1009|Yellow||2008-06-02|2008-06-17|2011-03-23|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||33.1||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|No||Neighbor/Friend|General Community||Match Support|F|Black||67|28215||Married|Education: Teacher||0|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500010765|500545186|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|8|||2230|7|||1|
500186138|500189040|500037040|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1726|Yellow||2004-05-04|2004-05-14|2009-02-03|Volunteer: Moved|Volunteer: Moved||56.7||1|1|1|1|M|Black||21||Mother|28208|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|White||45|28270|Masters Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187729|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501363890|500189279|500315105|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1377|Yellow||2008-11-14|2008-11-21|2012-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||45.2||1|1|2|2|M|Black||21|No|Mother|28216|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||37|28213|Masters Degree|Single|Medical: Healthcare Worker||2|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|501356607|31|0|1|31|0|1|10|2|-2||4|2||-2|500000294|-2|0|8|||7464|9|||1|
501045211|501132288|500239114|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1328|Green||2008-01-23|2008-01-23|2011-09-12|Child/Family: Moved|Child/Family: Moved||43.6||1|1|1|1|M|Black||21|No|GrandMother|28269|Grandparents|$20,000 to $24,999||||Yes||BBBS Board/Staff|General Community||Match Support|M|Black||47|28226|Bachelors Degree|Married|Business: Marketing||1|2|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501045484|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|13|||7671|13|||1|
500874202|501251394|500274520|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|299|Green||2008-06-23|2008-06-30|2009-04-25|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||9.8||1|1|1|1|M|Black||21|No|Mother|28205|One Parent: Female|$35,000 to $39,999||||No||Self|General Community||Enrollment|M|White||35|28203|Bachelors Degree|Single|Customer Service|28255|2|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500874471|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500261314|501842294|500426381|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|216|Yellow||2010-01-12|2010-01-20|2010-08-24|Child/Family: Time constraints|Child/Family: Time constraints||7.1||2|2|1|1|M|Hispanic||21||Mother|28213|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||36|28262|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|500261329|3|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501340105|501514453|500322778|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1658|Red|Amachi|2008-12-04|2008-12-12|2013-06-27|Child: Graduated|Child: Graduated||54.5||1|1|1|1|F|Multi-race (Black & Hispanic)||21|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||53|28269||Married|Medical: Admin||4|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501340376|38|0|2|1|0|2|10|2|-2||4|3|500000294|-2||-2|0|10|||7464|9|||1|500000294
502108064|502146885|500460150|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1295|Yellow||2010-07-07|2010-07-22|2014-02-06|Child: Graduated|Child: Graduated||42.5||1|1|1|1|F|White||21|No|Father|28277|One Parent: Male|Unknown||||No||Relative|General Community||Match Support|F|White||48|28277|High School Graduate|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502108491|1|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|3|||7464|9|||1|
500848341|500851040|500175773|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1035|Red||2007-05-04|2007-05-08|2010-03-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||34||1|1|1|1|M|Black||21|No|Mother|28277|One Parent: Female|$40,000 to $44,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||38|29732|||Business: Clerical||4|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500848610|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||46|2|||1|
500186765|500189359|500037396|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3266|Green||2004-09-15|2004-09-05|2013-08-15|Child: Graduated|Child: Graduated||107.3||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||46|28078|Masters Degree|Widowed|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500004169|500188083|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501811375|501391123|500374230|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1493|Yellow||2009-07-16|2009-07-27|2013-08-28|Child: Graduated|Child: Graduated||49.1||1|1|3|3|F|Black||21|No|Mother|28027|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|Black||41|28027|PHD|Single|Medical: Doctor, Provider|28075|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|501811730|31|0|2|31|0|2|10|2|-2||4|2||-2|500016374|-2|0|8|||7464|9|||1|
502221899|502188288|500461229|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|707|Green|Amachi|2010-07-15|2010-07-22|2012-06-28|Child: Severity of challenges|Child: Severity of challenges||23.2||1|1|1|1|F|Black||21|Yes|Mother|28216|One Parent: Female|Unknown||||Yes|Arby's|Workplace Partner/Business|General Community||Match Support|F|White||33|28262|Masters Degree|Single|Govt: Mgmt/Admin||5|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|502222330|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|3394|14|||7464|9|||1|500000294
500185734|500188688|500036688|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3592|Red||2003-10-15|2003-10-15|2013-08-15|Child: Graduated|Child: Graduated||118||1|1|1|1|F|Black||21||Mother|28203|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|White||45|28202|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500004169|500187476|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|8|||7464|9|||1|
500903146|501299088|500287883|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|665|Green|Amachi|2008-09-12|2008-09-30|2010-07-27|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||21.8||2|2|1|1|M|Black||21|No|Mother|28211|One Parent: Female|Less than $10,000|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Enrollment|M|Black||48|28105|Some College|Single|Finance: Accountant|28217|7|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500903416|31|0|1|31|0|1|5|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||7453|7|||1|500000294
500791133|500459674|500164598|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1157|Yellow|Amachi|2007-03-02|2007-03-06|2010-05-06|Child/Family: Moved|Child/Family: Moved||38||1|1|4|4|F|Black||21|Yes|Mother|28269|One Parent: Female|$35,000 to $39,999||||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||38|28219||Single|Finance: Banking|28273|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001281|500791401|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|6854|8|||2238|7|||1|500000294
500763132|500956022|500257067|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|630|Green|Amachi|2008-04-07|2008-04-09|2009-12-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.7||2|2|2|2|F|Black||21|Yes|Mother|28208|Other/Unknown|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||41|28277|Bachelors Degree|Single|Business: Mgt, Admin||9|0|General|Other Big|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500003657|500763400|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|5635|9|||6450|12|||1|500000294
501672971|500868727|500365034|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|302|Yellow||2009-05-22|2009-06-15|2010-04-13|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||9.9||1|1|4|4|F|Black||21|No|Mother|28205|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|Black||38|28214|Bachelors Degree|Single|Business: Clerical|28273|2|3|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|501673309|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|8|||7464|9|||1|
501021329|501035673|500235713|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|396|Green||2008-01-07|2008-01-08|2009-02-07|Volunteer: Moved|Volunteer: Moved||13||1|1|1|1|F|Black||21|No|Mother|28215|One Parent: Female|Less than $10,000||||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|Black||31|28215|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501021602|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|34|2|||46|2|||1|
500186938|500189708|500037821|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2675|Yellow|Amachi|2004-08-24|2004-08-24|2011-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||87.9||1|1|1|1|F|Black||21||Mother|28215|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||40|28217|Bachelors Degree|Single|Finance: Accountant|28277|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188131|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500539983|500540103|500143721|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1457|Yellow||2006-11-28|2006-12-05|2010-12-01|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||47.9||1|1|1|1|M|Black||21|No|Mother|28078|One Parent: Female|$25,000 to $29,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||47|28078|Some College|Married|Business: Mgt, Admin|3801|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500010765|500540234|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|34|2|||46|2|||1|
500186646|500189263|500047741|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2895|Yellow||2005-10-20|2005-10-20|2013-09-23|Child: Graduated|Child: Graduated||95.1||3|3|3|3|F|Some Other Race||21||Mother|28217|Other/Unknown|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|Black||39|28216|Some College||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|500188044|41|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|8|||7464|9|||1|
500392419|500746900|500162012|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2368|Yellow||2007-02-21|2007-03-06|2013-08-29|Child/Family: Moved|Child/Family: Moved||77.8||2|2|1|1|F|Black||21||Father|28105|One Parent: Male|Unknown||||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||32|28277||Single|Business: Sales||0|5|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011746|500392669|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|6855|8|||7464|9|||1|
501253984|500914930|500256894|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|482|Green|Amachi|2008-04-04|2008-04-09|2009-08-04|Child/Family: Moved|Child/Family: Moved||15.8||1|1|2|2|F|Black||21|No|Mother|28213|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||42|28027|Bachelors Degree|Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001262|501254241|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500478936|501284751|500275964|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1946|Green||2008-06-30|2008-07-14|2013-11-11|Child: Graduated|Child: Graduated||63.9||1|1|3|3|M|Black||21|No|Mother|28078|One Parent: Female|$25,000 to $29,999||||No||Neighbor/Friend|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|1|0|277|60|598|500000170|500017777|500479187|31|0|1|31|0|1|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|8|||132|8|||1|
501791114|501343064|500375189|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|419|Green||2009-07-23|2009-07-30|2010-09-22|Volunteer: Time constraint|Volunteer: Time constraint||13.8||1|1|1|1|F|Black||21|No|Mother|28262|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community||Match Support|F|Black||39|28215|Bachelors Degree|Single|Tech: Management|28202|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501791469|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|5|||7496|10|||1|
500850236|500189198|500169235|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2357|Green||2007-03-28|2007-04-04|2013-09-16|Child: Graduated|Child: Graduated||77.4||1|1|2|2|M|Black||21|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|M|Black||37|28262|Bachelors Degree|Single|Real Estate: Realtor||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011746|500850505|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500781988|500773716|500160560|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2392|Green||2007-02-14|2007-02-16|2013-09-04|Child/Family: Moved|Child/Family: Moved||78.6||1|1|1|1|M|White||21||Mother|28027||Unknown||||No||Self|General Community||Match Support|M|White||71|28083|Some College|Married|Business: Mgt, Admin|28027|13|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500782256|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500398853|500795095|500155431|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1603|Green|2010-2012 OJJDP JJI|2007-01-29|2007-02-16|2011-07-08|Child: Lost interest|Child: Lost interest||52.7||1|1|1|1|M|Black||21|No|Mother|28083|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||40|28269|Masters Degree|Married|Govt: Mgmt/Admin|28202|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500399103|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||2238|7|||1|500005291
500465511|500527675|500118120|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2628|Yellow|Amachi|2006-08-15|2006-08-21|2013-10-31|Child: Graduated|Child: Graduated||86.3||1|1|1|1|M|Black||21|Yes|Mother|28262|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|M|White||54|28210|Masters Degree|Married|Finance: Accountant||0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500465757|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2|500000294|-2|0|4|||2230|7|||1|500000294
501535013|501609664|500351430|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|848|Yellow||2009-03-23|2009-03-26|2011-07-22|Volunteer: Moved|Volunteer: Moved||27.9||1|1|1|1|M|Black||21|No|Mother|28273|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||36|28277|Bachelors Degree|Single|Retail: Mgt|28105|3|3|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|501535305|31|0|1|31|0|1|10|2|-2||4|2||-2|500000294|-2|0|10|||7496|10|||1|
500903951|501167853|500252953|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1789|Yellow|Amachi|2008-03-18|2008-04-04|2013-02-26|Child: Lost interest|Child: Lost interest||58.8||1|1|1|1|M|Black||21|Yes|Mother|28203|One Parent: Female|Less than $10,000|||Y|No||Faith Organization|General Community|Amachi|Match Support|M|White||34|28202|Bachelors Degree|Single|Finance: Banking||3|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500012459|500904221|31|0|1|1|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
502222992|502085103|500461244|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1245|Green||2010-07-16|2010-07-16|2013-12-12|Child: Graduated|Child: Graduated||40.9||1|1|1|1|F|Black||21|No|Aunt|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||32|28213|Bachelors Degree|Single|Education|28223|7|0|BBBS National Site|Web Link|Big|General Site||Enrollment|0|1|1|0|277|60|598|500000170|500017732|502223423|31|0|2|31|0|2|10|2|-2||4|1||-2||-1|6854|8|||46|2|||1|
501560189|501388335|500337198|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|180|Green||2009-01-30|2009-02-05|2009-08-04|Volunteer: Moved|Volunteer: Moved||5.9||2|2|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||40|28202|Bachelors Degree|Living w/ Significant Other|Business: Marketing|28202|1|1|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500001281|501560485|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501560189|501621478|500439156|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|806|Green||2010-03-04|2010-03-11|2012-05-25|Volunteer: Moved|Volunteer: Moved||26.5||2|2|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||39|28273||Single|Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501560485|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500713145|500932892|500187379|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1218|Green|Amachi|2007-08-08|2007-08-30|2010-12-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||40||1|1|1|1|M|Black||21|Yes|GrandMother|28227|One Parent: Female|Less than $10,000|||Y|No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||48|28227||Married|Military||21|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500713412|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500380928|500836517|500186930|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|605|Green||2007-08-02|2007-09-07|2009-05-04|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||19.9||2|2|1|1|F|Black||21||GrandMother|28216|One Parent: Female|Unknown||||No||Service Organization|General Community||Enrollment|F|Black||47|28216||Single|Finance: Banking|28216|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500381178|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|11|||46|2|||1|
500867581|500708515|500195388|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2323|Green|Amachi|2007-09-13|2007-09-28|2014-02-06|Child: Graduated|Child: Graduated||76.3||1|1|2|2|M|Black||21|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999||||No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||40|28269|Masters Degree|Single|Finance: Accountant|28255|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500015820|500867843|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|5635|9|||2238|7|||1|500000294
500480596|500491267|500120915|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2682|Green|Amachi|2006-09-05|2006-09-13|2014-01-16|Child: Graduated|Child: Graduated||88.1||1|1|1|1|M|Black||21|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Married|Business: Sales|28203|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500480847|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
500185627|500191338|500056611|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1354|Red||2005-11-14|2005-11-14|2009-07-30|Child: Severity of challenges|Child: Severity of challenges||44.5||1|1|1|1|M|American Indian or Alaska Native||21||Mother|28031|Other/Unknown|Unknown||||No||Faith Organization|General Community||Match Support|M|White||66|28031||Married|Business: Human Resources||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500001267|500187261|6|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|9|||7496|10|||1|
500382619|500385268|500085979|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1081|Green|Amachi|2006-03-23|2006-04-10|2009-03-26|Volunteer: Lost contact with child/agency Child/Family: Lost contact with volunteer/agency|Volunteer: Lost contact with child/agency|Child/Family: Lost contact with volunteer/agency|35.5||1|1|1|1|M|Black||21|Yes|Mother|28083|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|M|White||40|28081|Bachelors Degree|Single|Finance: Banking|28117|0|1|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001262|500382869|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294
500186352|500189280|500037290|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4175|Green||2002-07-29|2002-07-29|2014-01-02|Child: Graduated|Child: Graduated||137.2||4|4|2|2|M|Black||21||Mother|28212|One Parent: Female|Unknown|||Y|No|Big|Neighbor/Friend|General Community||Match Support|M|White||45|28226|Masters Degree|Married|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|500187945|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|6854|8|||7496|10|||1|
500186352|500189260|500037267|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4175|Green||2002-07-29|2002-07-29|2014-01-02|Child: Graduated|Child: Graduated||137.2||4|4|2|2|M|Black||21||Mother|28212|One Parent: Female|Unknown|||Y|No|Big|Neighbor/Friend|General Community||Match Support|F|White||40|28226|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|500187945|31|0|1|1|0|2|10|2|-2||4|1||-2||-2|6854|8|||7464|9|||1|
501227519|501216868|500255834|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|346|Green|Amachi|2008-03-31|2008-03-31|2009-03-12|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||11.4||1|1|3|3|M|Black||21|Yes|Mother|28025|Sibling Guardian|Unknown||||No||School|General Community|Amachi|Match Support|M|White||32|28078||Single|Education: Teacher||0|0|other|College Partner|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500001262|501227795|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||7670|5|||1|500000294
500187075|500189550|500037643|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3404|Green||2004-09-21|2004-09-21|2014-01-16|Child: Graduated|Child: Graduated||111.8||1|1|6|6|F|Black||21||Mother|28205|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||38|28209|Bachelors Degree|Single|Human Services: Non-Profit||0|0|Recruitment Event|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500012459|500188223|31|0|2|1|0|2|10|2|-2||4|1||-2||-1|0|10|||7458|9|||1|
501190094|500721829|500314463|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Red||2008-11-13|2008-11-20|2011-04-21|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29||1|1|1|1|F|Black||21||Aunt|28215|Two Mothers|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|F|Black||42|28215||Single|Business: Clerical||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501190365|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|34|2|||46|2|||1|
501343402|501371488|500287282|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|201|Green||2008-09-10|2008-09-18|2009-04-07|Vol: Lost Interest|Vol: Lost Interest||6.6||2|2|1|1|M|Some Other Race||21|No|Mother|28027|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||79|28025|Bachelors Degree|Divorced|Self-Employed, Entrepreneur|28025|0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|501343681|41|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
501343402|501567853|500355892|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|279|Green||2009-04-07|2009-04-07|2010-01-11|Volunteer: Time constraint|Volunteer: Time constraint||9.2||2|2|1|1|M|Some Other Race||21|No|Mother|28027|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||53|28027||Married|Business: Mgt, Admin|28027|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501343681|41|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501255133|501306527|500278242|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|681|Green||2008-07-17|2008-07-30|2010-06-11|Child: Lost interest|Child: Lost interest||22.4||2|2|4|5|F|White||21|No|Father|28025|One Parent: Male|Unknown||||Yes||Self|General Community||Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|1|0|1|0|277|60|598|500000170|500002335|501255409|1|0|2|1|0|2|10|2|-2||4|1||-2|500014681, 500016374|-2|0|10|||7464|9|||1|
500185890|500188833|500036833|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2020|Green||2005-04-09|2005-04-09|2010-10-20|Child/Family: Moved|Child/Family: Moved||66.4||1|1|1|1|M|White||21||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||54|28202||Married|Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500187556|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500916976|501262371|500273621|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|843|Green|Amachi|2008-06-17|2008-09-08|2010-12-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||27.7||1|1|1|1|M|Black||21|Yes|Mother|28216|One Parent: Female|$20,000 to $24,999||||Yes||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||35|28269|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500917246|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|8|||7496|10|||1|500000294
501622497|501446203|500350734|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1032|Green||2009-03-19|2009-03-31|2012-01-27|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||33.9||1|1|1|1|M|Black||21|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||43|28227||Married|Business: Engineer|28227|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501622817|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501626199|501293622|500351814|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1649|Green||2009-03-24|2009-03-26|2013-09-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||54.2||1|1|1|1|F|Black||21|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||33|28203|Masters Degree|Single|Finance: Accountant|28211|1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|501622822|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501508070|501447548|500334682|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|239|Green||2009-01-21|2009-01-27|2009-09-23|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||7.9||1|1|1|1|M|Black||21|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||33|28078|Bachelors Degree|Single|Tech: Engineer|28078|1|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501508362|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500767208|501341042|500276669|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2083|Green|Project Big|2008-07-07|2008-07-10|2014-03-24|Child: Graduated|Child: Graduated||68.4||1|1|1|1|F|Black||21||Mother|28216|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|Black||32|28216|Masters Degree|Single|Human Services|28215|0|7|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Enrollment|1|0|1|0|277|60|598|500000170|500017732|500767473|31|0|2|31|0|2|10|2|500004641||4|1||-2|500014506|-1|0|10|||7671|13|||1|500004640
500186943|500224697|500048942|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2120|Green|Amachi|2005-10-26|2005-10-26|2011-08-16|Volunteer: Time constraint|Volunteer: Time constraint||69.7||2|2|1|1|F|Black||21||Mother|28269|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||40|28297|||Human Services: Social Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188139|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
501130354|501124346|500245525|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1749|Red|Amachi|2008-02-15|2008-02-15|2012-11-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||57.5||1|1|1|1|M|Black||21|Yes|Mother|28213|One Parent: Female|Less than $10,000|||Y|Yes||BBBS Board/Staff|General Community|Amachi|Match Support|M|White||43|28205|Bachelors Degree|Married|Finance: Banking||7|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501130628|31|0|1|1|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|13|||46|2|||1|500000294
500483980|500423426|500120592|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2761|Green||2006-09-01|2006-09-01|2014-03-24|Child: Graduated|Child: Graduated||90.7||1|1|2|2|M|Black||21||Mother|28227|One Parent: Female|$10,000 to $14,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||71|28270||Single|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|500484231|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|6854|8|||7464|9|||1|
500185691|500188680|500036680|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2100|Green||2004-02-04|2004-02-04|2009-11-04|Volunteer: Moved|Volunteer: Moved||69||1|1|1|1|M|Black||21||GrandMother|28206|Other/Unknown|Unknown||||No|Brochure|Media|General Community||Match Support|M|White||44|28206||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500187323|31|0|1|1|0|1|10|2|||4|1||-2||-2|51|1|||7496|10|||1|
501201068|501771844|500396764|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1034|Green||2009-10-19|2009-10-30|2012-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||34||1|1|1|1|M|Black||21|No|Mother|28215|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||60|28262|Masters Degree|Single|Tech: Engineer||5|0|AA Task Force|Service Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|501201342|31|0|1|31|0|1|10|2|-2||4|1||-2|500000294|-2|6854|8|||9226|6|||1|
501618778|501610596|500353343|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|217|Green||2009-03-30|2009-04-08|2009-11-11|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||7.1||1|1|2|2|M|Black||21|No|Mother|28083|One Parent: Female|Unknown||||No||Workplace Partner/Business|General Community||Enrollment|M|Black||42|28027|Bachelors Degree|Single|Finance|28262|0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500001262|501618544|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|14|||7464|9|||1|
500186169|500189147|500037147|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1975|Red||2004-11-09|2004-11-09|2010-04-07|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||64.9||1|1|1|1|F|Black||21||Mother|28204|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||36|28278|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500187754|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501994934|501930790|500457779|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|395|Green||2010-06-22|2010-06-29|2011-07-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13||1|1|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||||No||BBBS Board/Staff|General Community||Match Support|F|Black||29|28202|||Tech: Production Line||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501843047|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|13|||7464|9|||1|
502294587|502389185|500499438|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|87|Green||2010-11-24|2010-12-07|2011-03-04|Volunteer: Moved|Volunteer: Moved||2.9||1|1|1|1|M|Black||21|No|Mother|28215|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||31|28204|Juris Doctorate (JD)|Single|Law: Lawyer|28280|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|501712404|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|6854|8|||7496|10|||1|
500185593|500234684|500062071|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1969|Yellow||2005-12-05|2005-12-05|2011-04-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||64.7||1|1|2|2|M|Black||21||Mother|28262|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||34|28213|Bachelors Degree|Single|Finance: Banking|28202|0|2|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187227|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|8|||7458|9|||1|
500877524|501077565|500229736|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|928|Yellow||2007-12-11|2007-12-15|2010-06-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||30.5||1|1|1|1|M|Black||21|No|Mother|28273|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||RTBM|M|Black||35|28213|Bachelors Degree|Single|Human Services: Youth Worker|28025|1|6|AA Task Force|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500877793|31|0|1|31|0|1|7|2|-2||4|2||-2||-2|0|10|||6247|12|||1|
501296349|501471640|500318555|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1914|Yellow||2008-11-20|2008-12-01|2014-02-27|Child: Graduated|Child: Graduated||62.9||1|1|1|1|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||42|28214|Bachelors Degree|Single|Business: Mgt, Admin|28205|3|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500012459|501296627|31|0|2|31|0|2|10|2|||4|2||-2|500000294|-2|0|4|||7464|9|||1|
501086649|501833794|500399391|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1146|Red||2009-10-23|2009-11-20|2013-01-09|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||37.7||1|1|1|1|M|Black||21|No|Mother|28216|One Parent: Female|$20,000 to $24,999||||Yes||Relative|General Community||Match Support|M|White||39|28205|Bachelors Degree|Single|Transport: Pilot|30320|2|0|Other Church Partner|Faith Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|501086923|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|3|||7453|7|||1|
500897083|501862348|500407273|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1102|Red|Amachi|2009-11-06|2009-11-13|2012-11-19|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||36.2||1|1|1|1|M|Black||21|Yes|Mother|28269|One Parent: Female|Unknown|||Y|No||Service Organization|General Community|Amachi|Match Support|M|White||54|28210||Married|Self-Employed, Entrepreneur||0|0|Holy Comforter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500015820|500897335|31|0|1|1|0|1|10|2|-2||4|3|500000294|-2|500000294|-2|0|11|||9216|7|||1|500000294
500981435|501623866|500374604|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|524|Red||2009-07-20|2009-07-24|2010-12-30|Volunteer: Time constraint|Volunteer: Time constraint||17.2||2|2|1|1|F|Multi-Race (None of the above)||21|No|Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||42|28203|||Business: Mgt, Admin|28210|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|500981706|7|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500981435|501130006|500241571|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|487|Red||2008-02-01|2008-02-07|2009-06-08|Volunteer: Moved|Volunteer: Moved||16||2|2|1|1|F|Multi-Race (None of the above)||21|No|Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||38|28205|Bachelors Degree|Single|Human Services: Non-Profit||1|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500981706|7|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7446|3|||1|
500185463|501470938|500330778|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|142|Green|Amachi|2009-01-06|2009-01-31|2009-06-22|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||4.7||2|2|1|1|M|Black||21|Yes|Non-Relative: Other|28205|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||35|28204||Single|Finance: Banking|28207|1|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|500187095|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
500186170|500648150|500147412|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1038|Red||2006-12-12|2006-12-13|2009-10-16|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||34.1||2|2|1|1|M|Black||21||Mother|28216|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|White||37|28209|Bachelors Degree|Single|Education: Teacher||0|0|General|Other Big|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500009007|500187755|31|0|1|1|0|2|10|2|-2||4|3||-2||-2|0|10|||6450|12|||1|
501614157|501596246|500374258|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1345|Green||2009-07-16|2009-07-29|2013-04-04|Volunteer: Moved|Volunteer: Moved||44.2||1|1|1|1|F|Black||21|No|Mother|28202|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||33|28273|||Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|501614477|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186071|500189012|500037012|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3768|Green||2004-01-05|2004-01-05|2014-04-30|Child: Graduated|Child: Graduated||123.8||1|1|1|1|M|White||21|No|Mother|28277|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||40|28277|Masters Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500187670|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500185897|500549520|500155451|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2552|Red|Project Big|2007-01-29|2007-02-05|2014-01-31|Child: Graduated|Child: Graduated||83.8||2|2|1|1|M|Black||21|No|Relative: Other|28208|Other Relative|Unknown||||No||Self|General Community||Match Support|M|White||39|28277|Bachelors Degree|Single|Tech: Computer/Programmer||4|0|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008321|500187458|31|0|1|1|0|1|10|2|500004641||4|3||-2||-2|0|10|||46|2|||1|500004640
500922736|501248121|500278235|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|171|Green||2008-07-17|2008-08-04|2009-01-22|Vol: Lost Interest|Vol: Lost Interest||5.6||1|1|1|1|F|Black||21|No|Mother|28083|One Parent: Female|Unknown||||No||School|General Community||Enrollment|F|Black||33|28025||Single|Finance: Banking|28262|0|0|TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500923006|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|4|||130|1|||1|
500552971|500565140|500147762|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1105|Green||2006-12-12|2006-12-13|2009-12-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||36.3||1|1|1|1|M|Black||21||Mother|28269|One Parent: Female|$30,000 to $34,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|Black||56|28078|Bachelors Degree|Married|Finance: Banking||9|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500553223|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
500186665|500189566|500037664|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3145|Red||2004-07-20|2004-07-20|2013-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||103.3||1|1|1|1|M|Black||21||Mother|28202|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|Black||40|28207||Single|Medical: Nurse||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500188050|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
501791424|501310838|500373905|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|350|Yellow||2009-07-14|2009-07-27|2010-07-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.5||1|1|1|1|F|Black||21|No|Mother|28202|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||32|28212|Some College|Single|Tech: Production Line|28212|2|9|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501791779|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7438|1|||1|
500344292|501166827|500341565|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|174|Yellow|Amachi|2009-02-17|2009-02-27|2009-08-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.7||2|2|1|1|F|Black||21|Yes|Mother|28205|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||30|28213|||Student: College||0|0|other|College Partner|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|500344425|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7670|5|||1|500000294
500186853|500189632|500037741|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2640|Yellow||2004-11-04|2004-11-04|2012-01-27|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||86.7||1|1|1|1|M|Black||21||Mother|28210|Other/Unknown|Unknown||||No||Self|General Community||Match Support|M|Black||36|28203|Bachelors Degree||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500264223|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500998929|502332678|500497432|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|284|Green|Amachi|2010-11-18|2010-11-19|2011-08-30|Volunteer: Moved|Volunteer: Moved||9.3||1|1|1|1|F|Black||21|Yes|Mother|28212|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|Amachi|Match Support|F|White||29|28204|Bachelors Degree|Single|Medical: Nurse|28202|0|0|Big Champions|Other Big|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008629|500999202|31|0|2|1|0|2|10|2|-2||4|1|500000294|-2|500000294, 500004640|-2|0|10|||7461|12|||1|500000294
500924153|500954048|500209749|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|741|Green||2007-10-25|2007-10-31|2009-11-10|Child: Severity of challenges|Child: Severity of challenges||24.3||1|1|1|1|M|Multi-Race (None of the above)||21|No|Mother|28277|One Parent: Female|$40,000 to $44,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||46|28277||Divorced|Business: Sales||11|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500924423|7|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
500910040|501600417|500363806|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1805|Red||2009-05-14|2009-05-29|2014-05-08|Child: Graduated|Child: Graduated||59.3||1|1|1|1|M|White||21|No|Mother|28270|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||31|28209|||Human Services: Non-Profit|28273|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|500910310|1|0|1|1|0|1|10|2|||4|3||-2||-2|0|10|||7464|9|||1|
500186427|501362883|500297556|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|293|Green||2008-10-10|2008-10-15|2009-08-04|Volunteer: Moved|Volunteer: Moved||9.6||3|3|1|1|M|Black||21||GrandMother|28202|One Parent: Female|Unknown||||No|Brochure|Media|General Community||Match Support|M|Black||41|28262|Some College|Single|Self-Employed, Entrepreneur|28216|1|6|Radio|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187983|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|51|1|||131|1|||1|
500186427|501811850|500380093|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|96|Green||2009-08-20|2009-08-27|2009-12-01|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.2||3|3|3|3|M|Black||21||GrandMother|28202|One Parent: Female|Unknown||||No|Brochure|Media|General Community||Match Support|M|White||36|28202|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009242|500187983|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|51|1|||7464|9|||1|
501164174|501241280|500276864|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|704|Green|Amachi|2008-07-08|2008-08-22|2010-07-27|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||23.1||1|1|1|1|F|Black||21|Yes|Mother|28212|One Parent: Female|$50,000 to $59,999||||No||Self|General Community|Amachi|Match Support|F|Black||36|28273|Some College|Single|Business: Clerical|28255|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501164448|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||2238|7|||1|500000294
501389722|500787778|500337267|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1903|Green||2009-01-30|2009-02-06|2014-04-24|Child: Graduated|Child: Graduated||62.5||1|1|1|1|F|White||21|No|Mother|28027|Two Parent|Unknown||||No||Self|General Community||Match Support|F|White||56|28027||Divorced|Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500012459|501390003|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500954724|500922418|500187226|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1396|Yellow||2007-08-07|2007-08-21|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||45.9||1|1|1|1|F|Black||21|No|GrandMother|28273|One Parent: Female|Less than $10,000|||Y|No||Service Organization|General Community||Match Support|F|Black||38|28273|||Finance: Accountant||0|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500954994|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|11|||46|2|||1|
500946666|500982086|500198334|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1113|Red||2007-09-26|2007-10-09|2010-10-26|Volunteer: Moved|Volunteer: Moved||36.6||1|1|1|1|M|Black||21|No|Mother|28227|One Parent: Female|$30,000 to $34,999||||Yes||Neighbor/Friend|General Community||Match Support|M|Black||35|28212|Bachelors Degree|Single|Finance: Banking||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500946936|31|0|1|31|0|1|10|2|||4|3||-2||-2|0|8|||46|2|||1|
500190624|501129024|500344200|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|365|Red||2009-02-24|2009-03-10|2010-03-10|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||12||2|2|2|2|M|Black||21||Mother|28227|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|Black||44|28212|Bachelors Degree|Single|Law: Security Officer|28208|2|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|500190627|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501448470|501194872|500298923|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|654|Red||2008-10-14|2008-11-04|2010-08-20|Volunteer: Time constraint|Volunteer: Time constraint||21.5||1|1|1|1|F|White||21|No|Mother|28031|Two Parent|Unknown||||No||School|General Community||Match Support|F|White||38|28115|Some College|Single|Business: Clerical||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500010765|501448755|1|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||46|2|||1|
500185630|500542491|500688663|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|548|Green||2013-03-19|2013-03-19|2014-09-18|Child: Graduated|Child: Graduated||18||3|3|2|2|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||39|28211|High School Graduate|Single|Finance: Banking|28208|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|500187264|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
500185630|500542491|500122710|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2172|Green||2006-09-19|2006-09-26|2012-09-06|Child/Family: Time constraints|Child/Family: Time constraints||71.4||3|3|2|2|F|Black||21|No|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||39|28211|High School Graduate|Single|Finance: Banking|28208|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500187264|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
500185863|500188915|500036915|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3351|Green||2005-03-12|2005-03-12|2014-05-15|Child: Graduated|Child: Graduated||110.1||1|1|1|1|F|Black||20||Mother|28213|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||43|28202|Bachelors Degree|Married|Student: College||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|500187435|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501784421|501615736|500374160|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|418|Yellow||2009-07-15|2009-07-31|2010-09-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||13.7||1|1|1|1|F|Black||20|No|Mother|28206|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||33|28269|||Medical: Pharmacist|28203|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501784776|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501674375|501687861|500369936|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|269|Red||2009-06-18|2009-06-26|2010-03-22|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||8.8||1|1|1|1|F|Black||20|No|Mother|28203|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||45|28273|Associate Degree|Single|Business||15|0|Coca Cola|Workplace Partner|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|501674713|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||9610|3|||1|
500729762|501213239|500278874|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|358|Red||2008-07-22|2008-08-06|2009-07-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||11.8||2|2|1|1|F|Black||20|No|Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|No||School|General Community||Match Support|F|Black||45|28209|Bachelors Degree|Single|Human Services: Social Worker|28203|1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500730029|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||46|2|||1|
502245018|501811850|500469733|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|148|Green||2010-09-10|2010-09-21|2011-02-16|Volunteer: Moved|Volunteer: Moved||4.9||1|1|3|3|M|Hispanic||20|No|Mother|28217|One Parent: Female|Unknown||||No|Radio|Media|General Community||Match Support|M|White||36|28202|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|502245449|3|0|1|1|0|1|10|2|-2||4|1||-2||-2|55|1|||7464|9|||1|
502418103|502430938|500528075|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|152|Yellow|2010-2012 OJJDP JJI|2011-03-29|2011-04-08|2011-09-07|Child/Family: Moved|Child/Family: Moved||5||1|1|1|1|M|Black||20|No|Mother|28027|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28027|Bachelors Degree|Married|Business: Mgt, Admin|28273|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|502418541|31|0|1|31|0|1|10|2|-2||4|2|500005291|-2||-2|34|2|||7496|10|||1|500005291
500186141|501046739|500254296|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2219|Green||2008-03-25|2008-04-02|2014-04-30|Child: Graduated|Child: Graduated||72.9||3|3|1|1|F|Black||20|No|Mother|28213|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|Black||45|28269|Bachelors Degree|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500008321|500187731|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||46|2|||1|
501619710|501380737|500344198|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|815|Green||2009-02-24|2009-03-16|2011-06-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||26.8||1|1|1|1|M|Black||20|No|Mother|28208|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|M|Black||38|28211|Masters Degree|Single|Finance: Banking|28202|0|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501620030|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
500187090|500189320|500125754|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2521|Green||2006-10-04|2006-10-04|2013-08-29|Child: Graduated|Child: Graduated||82.8||2|2|3|3|F|Black||20||Mother|28216|Two Parent|Unknown||||No||School|General Community||Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|1|0|277|60|598|500000170|500012459|500188103|31|0|2|31|0|2|10|2|-2||4|1||-2|500016374|-2|0|4|||7464|9|||1|
500741571|500938541|500187546|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1609|Green||2007-08-09|2007-08-15|2012-01-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||52.9||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Some Other Race||31|28262|||Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500724899|31|0|1|41|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501987736|502109789|500456045|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1450|Green||2010-06-08|2010-06-29|2014-06-18|Child: Graduated|Child: Graduated||47.6||1|1|1|1|F|White||20|No|Father|28217|One Parent: Male|Unknown||||No|AARTF|Neighbor/Friend|General Community||Match Support|F|White||40|28203|Masters Degree|Single|Finance||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|501988135|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|6855|8|||7464|9|||1|
501868918|501921115|500454496|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1456|Green||2010-05-26|2010-05-27|2014-05-22|Child: Graduated|Child: Graduated||47.8||1|1|1|1|M|Black||20|No|Mother|28211|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||35|27612|Juris Doctorate (JD)|Living w/ Significant Other|Law|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|501869291|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500398862|500866741|500181635|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|689|Green||2007-06-20|2007-06-26|2009-05-15|Vol: Other Reason|Vol: Other Reason||22.6||1|1|1|1|F|Black||20||Mother|28227|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community||Enrollment|F|White||34|28205||Married|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500399109|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|5|||46|2|||1|
500383915|500540512|500274279|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1532|Green||2008-06-20|2008-06-20|2012-08-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||50.3||2|2|2|2|F|Black||20||GrandMother|28205|One Parent: Female|Unknown||||No|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||64|28269||Married|Finance: Economist||0|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008321|500384165|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|6855|8|||7464|9|||1|
501686310|501818631|500392214|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1230|Red||2009-10-07|2009-10-30|2013-03-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||40.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28211|One Parent: Female|Unknown||||No|Radio|Media|General Community||Match Support|M|Black||34|28202|Juris Doctorate (JD)|Single|Law: Lawyer||1|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501686648|36|0|1|31|0|1|10|2|-2||4|3||-2||-2|55|1|||7446|3|||1|
501249335|501482897|500328407|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|690|Green|Amachi|2008-12-19|2009-01-23|2010-12-14|Volunteer: Moved|Volunteer: Moved||22.7||1|1|1|1|M|White||20|Yes|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|RTBM|M|Some Other Race||28|28227|Some College|Single|Student: College|28205|6|2|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|501249611|1|0|1|41|0|1|7|2|500003586||4|1|500000294|-2||-2|0|10|||46|2|||1|500000294
500897406|500843337|500181575|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1218|Green|Amachi|2007-06-19|2007-06-26|2010-10-26|Volunteer: Moved|Volunteer: Moved||40||1|1|1|1|F|Black||20|Yes|Mother|28270|Two Parent|$20,000 to $24,999|||Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||37|28262|Masters Degree||Human Services: Social Worker||2|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501224558|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||7464|9|||1|500000294
501045216|500991938|500225279|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|850|Green||2007-11-30|2007-11-30|2010-03-29|Volunteer: Time constraint|Volunteer: Time constraint||27.9||1|1|1|1|F|Black||20|No|GrandMother|28269|Grandparents|$20,000 to $24,999||||Yes||BBBS Board/Staff|General Community||Enrollment|F|Black||49|28226|Associate Degree|Married|Self-Employed, Entrepreneur||20|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501045484|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|13|||7671|13|||1|
501045214|500953330|500217682|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2938|Green||2007-11-13|2007-11-30|2015-12-16|Child: Graduated|Child: Graduated||96.5||1|1|2|2|F|Black||20|No|Relative: Other|28269|Grandparents|$20,000 to $24,999||||Yes||BBBS Board/Staff|General Community||Match Support|F|Black||35|28213|Masters Degree|Single|Business||4|0|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|1|0|0|1|277|60|598|500000170|500002335|501045484|31|0|2|31|0|2|10|2|-2||4|1||-2|500014505, 500016394|-1|0|13|||46|2|||1|
501409296|501632500|500357952|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|919|Yellow||2009-04-17|2009-05-06|2011-11-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||30.2||1|1|1|1|M|Black||20|No|Mother|28278|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||54|28278|High School Graduate|Married|Tech: Management||0|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500001281|501409581|31|0|1|31|0|1|10|2|-2||4|2||-2|500007920, 500011315, 500011316|-2|0|10|||17159|12|||1|
500186206|500189157|500037157|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3140|Red||2005-02-24|2005-02-24|2013-09-30|Child/Family: Moved|Child/Family: Moved||103.2||1|1|1|1|M|Black||20||GrandMother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||44|28214|PHD|Married|Medical: Doctor, Provider||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500004169|500187812|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500185776|500188720|500036720|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1830|Green||2004-02-23|2004-02-23|2009-02-26|Volunteer: Moved|Volunteer: Moved||60.1||1|1|1|1|F|Black||20|No|Aunt|28216|One Parent: Female|Unknown||||No||Self|General Community||RTBM|F|Black||37|28227||Single|Human Services: Non-Profit|28205|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187366|31|0|2|31|0|2|7|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500357354|500824176|500169087|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|963|Green||2007-03-28|2007-04-27|2009-12-15|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.6||3|3|1|1|F|Hispanic||20|No|Mother|28208|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|Multi-Race (None of the above)||34|28277|Bachelors Degree|Single|Child/Day Care Worker||0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500357603|3|0|2|7|0|2|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
501967613|502311344|500498762|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|788|Yellow||2010-11-23|2010-12-31|2013-02-26|Volunteer: Time constraint|Volunteer: Time constraint||25.9||1|1|1|1|F|Black||20|No|Mother|28273|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Finance: Accountant|28277|3|5|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500012459|501968011|31|0|2|1|0|2|10|2|-2||4|2||-2|500000294, 500004640|-2|34|2|||7496|10|||1|
500896018|501225232|500269506|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2233|Green|Amachi|2008-06-02|2008-07-03|2014-08-14|Child: Graduated|Child: Graduated||73.4||1|1|1|1|F|Black||20|Yes|Mother|28027|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||40|28027|Bachelors Degree|Separated|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500896288|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
500858259|500773625|500174656|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|658|Green||2007-05-01|2007-05-01|2009-02-17|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||21.6||1|1|2|2|F|Black||20|No|Aunt|28025|Other Relative|Unknown||||No||Self|General Community||Match Support|F|Black||39|28083|Bachelors Degree|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|500858528|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500190264|500829745|500165110|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|953|Green|Amachi|2007-03-05|2007-03-20|2009-10-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||31.3||4|4|1|1|F|White||20|Yes|Mother|28083|One Parent: Female|Unknown||||No||Neighbor/Friend|General Site||Enrollment|F|White||50|28083|Bachelors Degree|Married|Real Estate: Realtor|28025|0|0||Other Big|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001262|500190267|1|0|2|1|0|2|5|2|500003586||4|1||-1|500000294|-2|0|8|||0|12|||1|500000294
501201092|501285276|500280817|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1343|Red||2008-08-06|2008-08-26|2012-04-30|Volunteer: Moved|Volunteer: Moved||44.1||1|1|1|1|M|White||20|No|Mother|28105|One Parent: Female|Unknown||||No||Relative|General Community||Match Support|M|White||35|28270|Bachelors Degree|Single|Tech: Engineer|48121|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011746|501201366|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|3|||7464|9|||1|
500186675|500865601|500185332|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2198|Red|Amachi|2007-07-19|2007-08-23|2013-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||72.2||4|4|1|1|F|Black||20|Yes|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||38|28221||Single|Human Services: Youth Worker||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500188055|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500227043|500205341|500149633|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1204|Yellow||2006-12-20|2006-12-21|2010-04-08|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||39.6||2|2|3|4|F|Black||20||Mother|28206|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||48|28213|Masters Degree|Divorced|Finance: Economist|28202|13|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500009007|500227051|31|0|2|31|0|2|10|2|-2||4|2||-2|500000294|-2|0|4|||46|2|||1|
500577339|501634485|500353354|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|813|Green||2009-03-30|2009-04-16|2011-07-08|Child/Family: Moved|Child/Family: Moved||26.7||1|1|1|1|M|Black||20|No|Mother|28083|Two Parent|Unknown||||No||Self|General Community||Match Support|M|White||37|28075|Some College|Married|Military||11|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|500577557|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7446|3|||1|
500892914|500826359|500267382|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|593|Green|Amachi|2008-05-16|2008-05-16|2009-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.5||2|2|2|2|M|Black||20|Yes|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28277|||Education: Teacher||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500893173|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|5|||2238|7|||1|500000294
500892914|501964388|500429157|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1668|Red|Amachi|2010-01-22|2010-02-16|2014-09-11|Child: Graduated|Child: Graduated||54.8||2|2|1|1|M|Black||20|Yes|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|White||30|28203|Bachelors Degree|Single|Business: Sales|28269|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|500893173|31|0|1|1|0|1|10|2|500003586||4|3|500000294|-2||-2|0|5|||7464|9|||1|500000294
501938310|501306527|500456460|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|60|Green||2010-06-11|2010-06-25|2010-08-24|Child: Lost interest|Child: Lost interest||2||1|1|4|5|F|White||20|Yes|Father|28081|Two Parent|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|0|1|1|0|277|60|598|500000170|500002335|501938708|1|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500014681, 500016374|-2|0|10|||7464|9|||1|
500186217|500541585|500139849|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1481|Yellow|Amachi|2006-11-13|2006-11-17|2010-12-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||48.7||3|4|1|1|M|Black||20|Yes|GrandMother|28216|Grandparents|$10,000 to $14,999|||Y|No||Neighbor/Friend|General Community|Amachi|RTBM|M|Black||55|28269||Married|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500010355|500187777|31|0|1|31|0|1|7|2|500003586||4|2|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500185842|500188911|500036911|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2624|Green||2004-12-02|2004-12-02|2012-02-08|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||86.2||1|1|1|1|M|Black||20||Mother|28206|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500008629|500187428|31|0|1|31|0|1|10|2|-2||4|1||-2||-1|0|10|||7464|9|||1|
501007512|501432962|500328182|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|125|Green|Amachi|2008-12-18|2009-01-08|2009-05-13|Child: Lost interest Child (or Parent): Does Not Like Vol|Child: Lost interest|Child (or Parent): Does Not Like Vol|4.1||1|1|1|1|F|Black||20||Mother|28215|One Parent: Female|Less than $10,000||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||63|28269|Some College|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500003657|501007785|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|5|||7464|9|||1|500000294
501680582|501457619|500375202|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|288|Red||2009-07-23|2009-07-28|2010-05-12|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||9.5||1|1|1|1|F|Black||20|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||43|28215|Some College|Single|Transport: Flight Attendant|32827|3|2|Self|Self|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500008629|501680920|31|0|2|31|0|2|10|2|||4|3||-2||-2|0|10|||7464|9|||1|
500801567|501834907|500391790|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1508|Green||2009-10-06|2009-10-26|2013-12-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||49.5||2|2|1|1|M|Black||20||Mother|28213|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||62|28078|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|500801835|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500801567|500814872|500167266|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|919|Green||2007-03-16|2007-03-20|2009-09-24|Volunteer: Moved|Volunteer: Moved||30.2||2|2|1|1|M|Black||20||Mother|28213|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||32|28205|Bachelors Degree|Single|Construction|28220|0|1|Recruitment Event|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500801835|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7460|12|||1|
500717519|500188838|500145722|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2456|Yellow||2006-12-05|2006-12-08|2013-08-29|Child: Lost interest|Child: Lost interest||80.7||1|1|2|2|M|Black||20||Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|No||School|General Community||Match Support|M|Black||37|28269|Bachelors Degree|Married|Education: Admin||0|0|Yahoo!|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011746|500717786|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|4|||32|2|||1|
500392858|501064465|500326650|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|745|Green||2008-12-15|2008-12-15|2010-12-30|Child/Family: Moved|Child/Family: Moved||24.5||3|3|2|2|M|Black||20||Aunt|28215|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community||Match Support|M|White||43|28227|High School Graduate|Married|Clergy||10|0|General|Other Big|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500393108|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|5|||6450|12|||1|
500186636|500452589|500102306|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1876|Green|Amachi|2006-06-27|2006-06-27|2011-08-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||61.6||2|2|1|1|F|Black||20||Mother|28208|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|F|Black||48|28277|Masters Degree|Married|Business: Sales||0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188037|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294
501217814|500995312|500265629|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|809|Green||2008-05-12|2008-05-19|2010-08-06|Volunteer: Moved|Volunteer: Moved||26.6||1|1|1|1|F|White||20|No|Mother|28027|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|F|White||29|28262|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501218090|1|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501228176|501279790|500279399|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1834|Red||2008-07-25|2008-08-05|2013-08-13|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||60.3||1|1|1|1|M|Black||20|No|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||33|28078|Masters Degree|Married|Finance: Auditor|28202|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|501228452|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
501072642|501204476|500322870|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|632|Yellow||2008-12-04|2008-12-15|2010-09-08|Child/Family: Time constraints|Child/Family: Time constraints||20.8||2|2|1|1|F|White||20|No|Mother|28134|One Parent: Female|$45,000 to $49,999||||No||Neighbor/Friend|General Community||Match Support|F|White||32|29732|Some College|Living w/ Significant Other|Business: Sales|28277|6|3|TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501072909|1|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|8|||130|1|||1|
500934359|500991215|500209165|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1139|Yellow|Amachi|2007-10-24|2007-11-08|2010-12-21|Volunteer: Time constraint|Volunteer: Time constraint||37.4||2|2|1|1|F|Black||20|Yes|Mother|28212|One Parent: Female|$10,000 to $14,999|||Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||35|28215|Bachelors Degree|Single|Business: Human Resources||3|0|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001281|500934629|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|0|9|||7671|13|||1|500000294
500472874|501179381|500278853|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1087|Red||2008-07-22|2008-08-06|2011-07-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.7||2|2|1|1|F|Black||20|No|Mother|28262|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||32|28262|Masters Degree|Single|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008062|500473122|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
502645489|502480739|500543463|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|369|Green|Project Big|2011-06-29|2011-06-30|2012-07-03|Child/Family: Moved|Child/Family: Moved||12.1||1|1|1|1|F|Black||20||Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||43|28214|Masters Degree|Married|Arts, Entertainment, Sports|28202|4|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502508948|31|0|2|31|0|2|10|2|500004641||4|1|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640
500763080|501173591|500250742|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|884|Green|Amachi|2008-03-06|2008-03-08|2010-08-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29||1|1|1|1|M|Black||20|No|Mother|28212|One Parent: Female|$20,000 to $24,999||||Yes||Faith Organization|General Community||Match Support|M|Hispanic||37|28202|Bachelors Degree|Single|Business: Engineer||1|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500763348|31|0|1|3|0|1|10|2|500003586||4|1||-2|500000294|-2|0|9|||46|2|||1|500000294
500186192|502323059|500490136|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1425|Green||2010-11-03|2010-11-18|2014-10-13|Child: Graduated|Child: Graduated||46.8||2|2|1|1|F|Black||20||Mother|28208|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||33|28208||Single|Service: Restaurant||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018987|500187762|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1|
500956278|501279041|500302301|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|698|Green||2008-10-21|2008-10-31|2010-09-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||22.9||1|1|1|1|F|Black||20|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|No||Neighbor/Friend|General Community||Match Support|F|White||35|28208|Juris Doctorate (JD)|Married|Law: Lawyer|28202|1|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500956548|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|0|8|||7464|9|||1|
500186101|500233328|500056732|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1311|Yellow||2005-11-14|2005-11-15|2009-06-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||43.1||2|2|1|1|M|White||20||Mother|28277|Other/Unknown|Unknown||||No||Self|General Community||Enrollment|M|White||44|28134|Some College|Married|Finance: Banking|28202|9|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500187695|1|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500747371|501279505|500329319|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|898|Yellow||2008-12-30|2008-12-31|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29.5||3|3|1|1|F|Black||20|No|Mother|28213|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|White||34|28025|Some College|Married|Business: Marketing|28262|11|0|Self|Self|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500008062|500747638|31|0|2|1|0|2|10|2|-2||4|2||-2|500000294|-2|0|4|||7464|9|||1|
500186791|500189594|500079732|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1420|Green|Amachi|2006-02-09|2006-02-09|2009-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||46.7||2|2|2|3|F|Multi-Race (None of the above)||20||Mother|28025|Other/Unknown|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|F|Black||38|28273|Bachelors Degree|Married|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188099|7|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
502552443|502471967|500537261|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1301|Green|Project Big|2011-05-20|2011-06-08|2014-12-30|Child: Graduated|Child: Graduated||42.7||1|1|1|1|F|Multi-race (Black & Hispanic)||20|No|GrandMother|28208|Grandparents|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28209|Bachelors Degree|Single|Medical|28209|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502552891|38|0|2|1|0|2|10|2|-2||4|1|500004640, 500005291|-2||-2|0|4|||7496|10|||1|500004640
500379986|500722764|500228460|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|846|Yellow||2007-12-10|2008-01-23|2010-05-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27.8||2|2|2|2|F|Black||20|Yes|Mother|28206|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Enrollment|F|Black||38|28217||Single|Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001281|500380236|31|0|2|31|0|2|5|2|-2||4|2||-2|500000294|-2|6854|8|||2238|7|||1|
500961015|501210561|500257073|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2365|Green|Amachi|2008-04-07|2008-04-11|2014-10-02|Child: Graduated|Child: Graduated||77.7||1|1|1|1|M|Black||20|Yes|Mother|28227|Two Parent|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||43|28104||Married|Tech: Computer/Programmer|29607|10|0|Relative|Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500934638|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||17161|11|||1|500000294
502646565|502528355|500543433|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|96|Green|Project Big, 2010-2012 OJJDP JJI|2011-06-29|2011-06-30|2011-10-04|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||3.2||1|1|2|2|M|Black||20|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502598113|31|0|1|1|0|1|10|2|500004641||4|1|500004640, 500005291|-2||-2|0|10|||132|8|||1|500004640, 500005291
501240369|501240602|500272039|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2282|Green|Amachi|2008-06-11|2008-07-10|2014-10-09|Child: Graduated|Child: Graduated||75||1|1|1|1|M|Black||20|Yes|Mother|28214|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|M|White||43|28269|Masters Degree|Single|Business: Mgt, Admin|28202|3|6|Radio|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501240645|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|3|||131|1|||1|500000294
502173811|500776552|500460247|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|416|Green|Amachi|2010-07-08|2010-07-13|2011-09-02|Volunteer: Moved|Volunteer: Moved||13.7||1|1|2|2|M|Black||20|Yes|Mother|28269|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|RTBM|M|Black||32|28202|Bachelors Degree|Single|Finance: Banking||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011184|502174240|31|0|1|31|0|1|7|2|500003586||4|1|500000294|-2||-2|7016|11|||46|2|||1|500000294
501676485|501684717|500369927|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|380|Red||2009-06-18|2009-07-13|2010-07-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.5||1|1|1|1|M|Black||20|No|Mother|28214|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|Black||43|28277|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501676823|31|0|1|31|0|1|5|2|||4|3||-2||-2|0|10|||7464|9|||1|
500261295|500188435|500073081|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4096|Green||2006-01-03|2005-12-21|2017-03-09|Child: Graduated|Child: Graduated||134.6||1|1|1|1|M|White||20||Mother|28104|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||60|28270|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Enrollment|1|0|0|1|277|60|598|500000170|500017732|500261310|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500320291|500516453|500121420|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1253|Yellow||2006-09-10|2006-09-26|2010-03-02|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||41.2||1|1|1|1|M|Black||20||Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||48|28205|Masters Degree|Single|Finance: Auditor|28202|3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500320412|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501070152|501052547|500224306|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1601|Yellow|Amachi|2007-11-28|2007-11-29|2012-04-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||52.6||1|1|2|2|M|Black||20|Yes|Mother|28212|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community|Amachi|Match Support|M|Black||45|28079|Bachelors Degree|Married|Business||13|6|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001281|501070425|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7671|13|||1|500000294
500780652|500189100|500164976|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1239|Green|Amachi|2007-03-05|2007-03-13|2010-08-03|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||40.7||1|1|3|3|F|Black||20|Yes|Mother|28208|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|Amachi|Match Support|F|Black||36|28269|Some College|Single|Customer Service||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500780920|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501164779|501159259|500251850|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1177|Green||2008-03-12|2008-03-27|2011-06-17|Volunteer: Moved|Volunteer: Moved||38.7||1|1|1|1|M|White||20|No|Mother|28210|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|White||40|22314|Bachelors Degree|Single|Business: Sales||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501165053|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500826592|501314246|500382768|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2567|Green||2009-09-04|2009-10-08|2016-10-18|Child: Graduated|Child: Graduated||84.3||3|3|1|1|F|Black||20|No|Mother|28226|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|F|White||33|28277|Bachelors Degree|Living w/ Significant Other|Unknown|28209|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|500826861|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|5|||7464|9|||1|
501012102|501519306|500348979|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|121|Green||2009-03-11|2009-03-17|2009-07-16|Child: Lost interest|Child: Lost interest||4||1|1|2|2|M|Black||20|No|Mother|28027|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500001262|501012375|31|0|1|1|0|1|10|2|-2||4|1||-2|500016374|-2|0|8|||7464|9|||1|
500896361|501276501|500291021|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1870|Yellow|Amachi|2008-09-24|2009-01-14|2014-02-27|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||61.4||2|2|1|1|F|Black||20|Yes|Mother|28208|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||51|28075||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500012459|500896631|31|0|2|31|0|2|10|2|-2||4|2|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501604440|501758365|500373108|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1945|Green||2009-07-08|2009-07-23|2014-11-19|Child: Graduated|Child: Graduated||63.9||1|1|1|1|M|Black||20|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Hispanic||38|28269||Married|Govt||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017732|501604760|31|0|1|3|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
500752612|500915297|500186913|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1400|Green||2007-08-02|2007-08-17|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||46||1|1|1|1|F|Black||20||Mother|28205|Foster Home|Unknown||||No||Self|General Community||Match Support|F|White||33|28207||Divorced|Consultant||5|0|TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500752880|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||130|1|||1|
501393942|501232528|500303603|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|138|Yellow||2008-10-23|2008-12-08|2009-04-25|Child (or Parent): Other Reason Vol: Other Reason|Child (or Parent): Other Reason|Vol: Other Reason|4.5||1|1|1|1|M|Black||20|No|Mother|28216|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||RTBM|M|White||30|28164|Some College|Single|Business: Sales||2|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|501394223|31|0|1|1|0|1|7|2|-2||4|2||-2||-2|0|8|||7464|9|||1|
501226817|501729866|500368063|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|307|Red|Amachi|2009-06-09|2009-07-09|2010-05-12|Volunteer: Time constraint|Volunteer: Time constraint||10.1||1|1|1|1|M|Black||20|Yes|Mother|28215|One Parent: Female|Unknown||||Yes||Relative|General Community|Amachi|Enrollment|M|Black||62|28269|Masters Degree|Married|Real Estate: Realtor||3|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501227093|31|0|1|31|0|1|5|2|-2||4|3|500000294|-2|500000294|-2|0|3|||2230|7|||1|500000294
500191424|502295287|500499432|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|379|Red|Amachi|2010-11-24|2010-12-16|2011-12-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12.5||3|3|2|2|F|Black||20|Yes|Mother|28031|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|White||47|28078|Juris Doctorate (JD)|Single|Law: Lawyer|28203|8|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011184|500191427|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2||-2|6854|8|||7464|9|||1|500000294
500191424|500998642|500222466|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1002|Yellow||2007-11-20|2007-12-11|2010-09-08|Volunteer: Moved|Volunteer: Moved||32.9||3|3|1|1|F|Black||20|Yes|Mother|28031|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Multi-Race (None of the above)||28|28035|Some College|Single|Student: College||0|0|Recruitment Event|College Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500191427|31|0|2|7|0|2|10|2|-2||4|2|500000294|-2||-2|6854|8|||7448|5|||1|
501042211|501089387|500251464|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|434|Green|Amachi|2008-03-11|2008-03-11|2009-05-19|Volunteer: Health|Volunteer: Health||14.3||1|1|1|1|M|White||20|Yes|Mother|28213|One Parent: Female|$10,000 to $14,999||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||66|28227|Associate Degree|Married|Tech: Production Line|28269|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501042484|1|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|34|2|||7464|9|||1|500000294
500186682|500887363|500184396|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2924|Green|Amachi|2007-07-13|2007-07-20|2015-07-22|Child: Graduated|Child: Graduated||96.1||3|4|1|1|M|Black||20|Yes|Mother|28227|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|Amachi|Match Support|M|Black||57|28262||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500188056|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502007951|502201951|500457933|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|120|Red||2010-06-23|2010-06-28|2010-10-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.9||1|1|1|1|M|Black||20|No|Mother|28216|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|M|Black||27|28215|Some College|Single|Student: College||4|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|502008350|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|8|||7464|9|||1|
502544191|502231024|500541173|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|930|Green|Amachi|2011-06-14|2011-06-21|2014-01-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||30.6||1|1|2|2|F|Black||20|Yes|Mother|28277|One Parent: Female|$50,000 to $59,999||||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||29|28277|Bachelors Degree|Single|Consultant|28204|0|11|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017777|502544644|31|0|2|1|0|2|10|2|-2||4|1|500000294|-2|500000294|-2|34|2|||46|2|||1|500000294
500185861|501357163|500360590|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|799|Green|Amachi|2009-04-30|2009-05-04|2011-07-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||26.3||3|4|1|1|F|Multi-Race (None of the above)||20|No|Mother|28211|Other/Unknown|Unknown||||No||School|General Community|Amachi|Enrollment|F|Black||53|28213|Some College|Single|Business: Sales||21|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500003657|501721919|7|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||7496|10|||1|500000294
500185601|501082220|500236473|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2733|Green||2008-01-09|2008-01-28|2015-07-23|Child: Graduated|Child: Graduated||89.8||2|2|1|1|M|Black||20||Mother|28210|Other/Unknown|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28078|High School Graduate|Single|Finance: Accountant|28202|0|4|Recruitment Event|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500012459|500187235|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|6854|8|||7458|9|||1|
500546821|500790181|500159910|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3128|Green||2007-02-13|2007-02-21|2015-09-15|Child: Graduated|Child: Graduated||102.8||1|1|3|3|M|Black||20|No|Mother|28083|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||52|28025||Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|1|0|0|1|277|60|598|500000170|500012459|500547073|31|0|1|31|0|1|10|2|-2||4|1||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7464|9|||1|
500185637|500189284|500073080|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3269|Green||2006-01-03|2005-12-29|2014-12-11|Child: Graduated|Child: Graduated||107.4||1|1|2|2|M|Black||20||Mother|28206|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|Black||55|28297|Masters Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500017732|500187271|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
500884730|500918341|500185843|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|798|Green||2007-07-24|2007-08-02|2009-10-08|Volunteer: Time constraint|Volunteer: Time constraint||26.2||1|1|1|1|M|White||20|No|Mother|28273|One Parent: Female|$45,000 to $49,999||||No|BBBS National Site|Web Link|General Community||Enrollment|M|White||38|29745|Bachelors Degree|Living w/ Significant Other|Business: Mgt, Admin|29732|4|7|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500884999|1|0|1|1|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
500186190|500189140|500037140|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3598|Yellow||2004-10-13|2004-10-13|2014-08-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||118.2||1|1|2|2|F|Black||20||Mother|28213|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|500187761|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501099098|500865864|500336493|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|61|Green|Amachi|2009-01-28|2009-02-20|2009-04-22|Vol: Lost Interest|Vol: Lost Interest||2||2|2|2|2|F|Black||20|Yes|Mother|28081|One Parent: Female|Unknown||||Yes||BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||35|28262||Single|Govt: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500002335|501099372|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|13|||2238|7|||1|500000294
501099098|502078407|500460269|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|138|Green||2010-07-08|2010-07-22|2010-12-07|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||4.5||2|2|2|2|F|Black||20|Yes|Mother|28081|One Parent: Female|Unknown||||Yes||BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||35|28083|Bachelors Degree|Single|Customer Service||5|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002335|501099372|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|13|||7464|9|||1|
502057399|502389976|500516780|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1127|Yellow|2010-2012 OJJDP JJI|2011-02-10|2011-02-28|2014-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||37||2|2|1|1|M|White||20|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||50|28078|Bachelors Degree|Single|Arts, Entertainment, Sports|28078|8|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502057823|1|0|1|1|0|1|10|2|-2||4|2|500005291|-2||-2|0|4|||7464|9|||1|500005291
502057399|502102663|500463696|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|164|Green||2010-07-30|2010-08-02|2011-01-13|Volunteer: Time constraint|Volunteer: Time constraint||5.4||2|2|1|1|M|White||20|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28031||Single|Finance||0|0|Recruitment Event|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011639|502057823|1|0|1|1|0|1|10|2|-2||4|1|500005291|-2|500000294|-2|0|4|||7458|9|||1|
500874765|502038804|500692473|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|833|Green||2013-04-11|2013-04-11|2015-07-23|Child: Graduated|Child: Graduated||27.4||4|4|2|2|F|Black||20|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|501755813|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|34|2|||7496|10|||1|
500874765|501587266|500356916|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|256|Green||2009-04-13|2009-04-24|2010-01-05|Volunteer: Time constraint|Volunteer: Time constraint||8.4||4|4|1|1|F|Black||20|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|White||34|28078|||Business: Marketing|28070|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501755813|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
500874765|502178791|500456682|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|426|Yellow||2010-06-14|2010-06-30|2011-08-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14||4|4|1|1|F|Black||20|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||29|28213|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501755813|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|34|2|||7464|9|||1|
502259491|501306527|500466849|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|782|Green||2010-08-24|2010-08-25|2012-10-15|Child: Lost interest|Child: Lost interest||25.7||1|1|4|5|F|White||20|No|Mother|28027|Two Parent|Unknown|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||31|28027|Some College|Married|Business: Clerical|28273|4|0|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Pending Match|0|1|1|0|277|60|598|500000170|500002335|502259924|1|0|2|1|0|2|10|2|-2||4|1||-2|500014681, 500016374|-2|0|5|||7464|9|||1|
500722500|500830633|500180184|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1589|Green||2007-06-14|2007-06-20|2011-10-26|Child/Family: Moved|Child/Family: Moved||52.2||2|2|1|1|F|White||20||Mother|28027||Unknown||||No||Service Organization|General Community||Match Support|F|White||34|28083|Bachelors Degree|Single|Education: Teacher Asst/Aid|28147|0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500722767|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|11|||7464|9|||1|
501287538|501420389|500336114|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|97|Green||2009-01-27|2009-01-27|2009-05-04|Child (or Parent): Other Reason|Child (or Parent): Other Reason||3.2||2|2|2|2|M|White||20|No|GrandMother|28025|Two Parent|Unknown||||No||Neighbor/Friend|General Community||RTBM|M|White||33|28107||Single|Law: Security Officer|28201|0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500002335|501287816|1|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
502142541|501905673|500455759|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1861|Green||2010-06-07|2010-06-18|2015-07-23|Child: Graduated|Child: Graduated||61.1||1|1|2|2|F|Black||20|No|Mother|28217|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|502142970|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1|
500934905|500915341|500185983|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|659|Green|Amachi|2007-07-25|2007-07-30|2009-05-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.7||1|1|1|1|F|Black||20|Yes|GrandMother|28216|One Parent: Female|Less than $10,000|||Y|No||Faith Organization|General Community|Amachi|Enrollment|F|Black||58|28262|Some College|Married|Retail: Mgt|28262|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500935173|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
500474486|500491064|500118168|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3282|Red||2006-08-16|2006-08-23|2015-08-18|Child: Graduated|Child: Graduated||107.8||1|1|1|1|M|Black||20||Mother|28214|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||38|28209|Bachelors Degree|Single|Construction|28247|0|2|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500474735|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|34|2|||7447|3|||1|
500845231|500360087|500320076|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|223|Yellow||2008-11-25|2008-12-02|2009-07-13|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.3||2|2|3|3|F|Black||20|No|Mother|28078|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Enrollment|F|Black||48|28070|Bachelors Degree|Single|Finance: Banking|28205|8|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500008629|500845500|31|0|2|31|0|2|5|2|-2||4|2||-2|500000294|-2|0|10|||2238|7|||1|
500969809|500940217|500230374|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|357|Red||2007-12-12|2008-02-07|2009-01-29|Agency: Concern with Volunteer re: child safety Volunteer: Moved|Agency: Concern with Volunteer re: child safety|Volunteer: Moved|11.7||1|1|1|1|M|Black||20||Mother|28205|Two Parent|Unknown||||No||Relative|General Community||Enrollment|M|White||59|28025|Bachelors Degree|Divorced|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500730811|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|3|||46|2|||1|
501860373|502078407|500505055|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|252|Green||2010-12-13|2010-12-16|2011-08-25|Volunteer: Time constraint|Volunteer: Time constraint||8.3||1|1|2|2|F|Black||20|No|GrandMother|28025|Grandparents|Unknown||||Yes|Brochure|Media|General Community||Match Support|F|Black||35|28083|Bachelors Degree|Single|Customer Service||5|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002335|501860746|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|51|1|||7464|9|||1|
501376516|501822933|500386771|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|303|Yellow|Amachi|2009-09-22|2009-09-30|2010-07-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||10||1|1|1|1|M|Black||20|Yes|Mother|28205|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Enrollment|M|White||34|28209|||Consultant||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|501376795|31|0|1|1|0|1|5|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
500186956|500189727|500037841|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3908|Green|Amachi|2004-06-21|2004-06-21|2015-03-04|Child: Graduated|Child: Graduated||128.4||1|1|1|1|M|Black||20||Mother|28213|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||54|28203|Bachelors Degree|Married|Law: Lawyer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500188141|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501099105|501033544|500458811|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|372|Green|Amachi|2010-06-28|2010-07-01|2011-07-08|Volunteer: Time constraint|Volunteer: Time constraint||12.2||2|2|2|2|F|Black||20|Yes|Mother|28081|One Parent: Female|Unknown||||Yes||Faith Organization|General Community|Amachi|Match Support|F|Some Other Race||35|28083|Some College|Divorced|Law: Police Officer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501099372|31|0|2|41|0|2|10|2|500003586||4|1|500000294|-2||-2|0|9|||2238|7|||1|500000294
501099105|501033544|500235298|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|847|Green|Amachi|2008-01-03|2008-01-11|2010-05-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27.8||2|2|2|2|F|Black||20|Yes|Mother|28081|One Parent: Female|Unknown||||Yes||Faith Organization|General Community|Amachi|Match Support|F|Some Other Race||35|28083|Some College|Divorced|Law: Police Officer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501099372|31|0|2|41|0|2|10|2|500003586||4|1|500000294|-2||-2|0|9|||2238|7|||1|500000294
502291098|500459674|500518681|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|236|Yellow|2010-2012 OJJDP JJI|2011-02-18|2011-03-03|2011-10-25|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.8||2|2|4|4|F|Black||20|No|Mother|28203|One Parent: Female|Unknown||||Yes|Brochure|Media|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||38|28219||Single|Finance: Banking|28273|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502291530|31|0|2|31|0|2|10|2|-2||4|2|500005291|-2|500000294|-2|51|1|||2238|7|||1|500005291
502291098|502597982|500575575|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|184|Yellow||2011-11-08|2011-11-23|2012-05-25|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||6||2|2|1|1|F|Black||20|No|Mother|28203|One Parent: Female|Unknown||||Yes|Brochure|Media|General Community|2010-2012 OJJDP JJI|Match Support|F|White||33|28273|Masters Degree|Single|Finance: Accountant|28202|4|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502291530|31|0|2|1|0|2|10|2|-2||4|2|500005291|-2||-2|51|1|||7464|9|||1|
502247430|502226106|500465539|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1255|Yellow||2010-08-12|2010-08-17|2014-01-23|Child: Lost interest|Child: Lost interest||41.2||1|1|1|1|F|Black||20|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||63|28078|Bachelors Degree|Married|Medical: Nurse||10|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|502247861|31|0|2|1|0|2|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1|
500408248|501258569|500359601|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|392|Green||2009-04-27|2009-04-27|2010-05-24|Volunteer: Time constraint|Volunteer: Time constraint||12.9||3|3|1|1|F|Black||20||Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|F|White||44|28203||Married|Law: Lawyer|28202|0|6|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002335|500187230|31|0|2|1|0|2|5|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
500408248|500725077|500206219|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|462|Red||2007-10-17|2007-10-25|2009-01-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||15.2||3|3|3|4|F|Black||20||Mother|28205|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|F|Black||34|28269|||Business: Marketing||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500187230|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|10|||46|2|||1|
500186106|500778380|500202993|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2856|Green||2007-10-11|2007-10-18|2015-08-13|Child: Graduated|Child: Graduated||93.8||2|2|1|1|F|Black||20||Mother|28217|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||35|28211|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018987|500187698|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500934903|500901552|500185986|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|729|Green|Amachi|2007-07-25|2007-07-30|2009-07-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24||1|1|1|1|F|Black||20|Yes|GrandMother|28216|One Parent: Female|Less than $10,000|||Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||36|28210|||Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500935173|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|9|||2238|7|||1|500000294
501114434|501315131|500324423|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1997|Red|Amachi|2008-12-09|2008-12-23|2014-06-12|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||65.6||1|1|1|1|M|Black||20|No|Uncle|28206|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||33|28207|Masters Degree|Single|Finance: Accountant|28244|0|0|TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501114708|31|0|1|1|0|1|10|2|-2||4|3|500000294|-2||-2|0|10|||130|1|11|3|1|500000294
500186435|500189358|500037395|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4411|Green||2003-07-23|2003-07-23|2015-08-20|Child: Graduated|Child: Graduated||144.9||1|1|1|1|M|Black||20||Mother|28216|One Parent: Female|Unknown||||No|Brochure|Media|General Community||Match Support|M|White||45|28226|Bachelors Degree|Married|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018987|500187988|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|51|1|||7496|10|||1|
502436202|502642999|500549046|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1410|Green||2011-08-08|2011-09-02|2015-07-13|Child: Graduated|Child: Graduated||46.3||1|1|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|Masters Degree|Single|Finance: Banking||0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502436645|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
500395038|500392006|500104016|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3125|Green||2006-07-06|2006-08-01|2015-02-20|Child: Graduated|Child: Graduated||102.7||1|1|1|1|M|White||20||Mother|28226|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||39|28211|Masters Degree|Married|Law: Lawyer|28204|2|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500395288|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
501626218|501587214|500350222|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2095|Green||2009-03-17|2009-03-24|2014-12-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||68.8||1|1|1|1|F|Black||20|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||30|11215|Bachelors Degree|Single|Consultant|11215|0|5|other|College Partner|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017732|501622822|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||7670|5|||1|
502278018|502813258|500597369|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|200|Red||2012-02-09|2012-02-12|2012-08-30|Child/Family: Moved|Child/Family: Moved||6.6||2|2|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||27|28212|Bachelors Degree|Single|Finance: Auditor|28262|0|4|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|502278450|31|0|1|1|0|1|10|2|||4|3||-2||-2|0|10|||7464|9|||1|
502278018|502227238|500477903|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|156|Yellow||2010-10-07|2010-10-25|2011-03-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.1||2|2|1|1|M|Black||20|No|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||26|28215|High School Graduate|Single|Unknown||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502278450|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
501522348|501223351|500349995|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1444|Red||2009-03-17|2009-03-17|2013-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||47.4||1|1|1|1|M|Multi-race (Black & White)||20|No|Mother|28031|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Single|Retail: Sales|28117|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501522640|36|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
501637367|501586552|500369810|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|315|Red||2009-06-17|2009-07-01|2010-05-12|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||10.3||2|2|1|1|F|Black||20||Mother|28214|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||32|28214|Associate Degree|Single|Student: College|28078|4|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501637690|31|0|2|1|0|2|10|2|||4|3||-2||-2|0|10|||7464|9|||1|
501637367|502606177|500555854|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|334|Green|Project Big|2011-09-19|2011-09-30|2012-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||11||2|2|1|1|F|Black||20||Mother|28214|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black|Other African|33|28209|Juris Doctorate (JD)|Single|Medical: Doctor, Provider|28012|1|0||Relative|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008629|501637690|31|0|2|31|31|2|10|2|-2||4|1||-2|500004640|-2|0|10|||0|11|||1|500004640
500566163|500989942|500236985|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1086|Green||2008-01-11|2008-01-23|2011-01-13|Volunteer: Time constraint|Volunteer: Time constraint||35.7||2|2|1|1|F|Black||20|No|Mother|28269|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Enrollment|F|Black||37|28213|Masters Degree|Single|Human Services: Social Worker||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500565754|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|34|2|||46|2|||1|
500876141|500899158|500183024|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1349|Yellow|Amachi|2007-07-05|2007-07-27|2011-04-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||44.3||1|1|1|1|M|Black||20|Yes|Mother|28216|One Parent: Female|$10,000 to $14,999|||Y|No||Faith Organization|General Community|Amachi|Match Support|M|Black||62|28216||Married|Clergy||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500876410|31|0|1|31|0|1|10|2|-2||4|2|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
500186432|501235725|500332721|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|669|Yellow||2009-01-14|2009-01-30|2010-11-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||22||4|4|1|1|F|Black||20||Mother|28212|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||34|28210|Masters Degree|Single|Medical: Healthcare Worker|28208|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|500187945|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501347056|501217000|500322327|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2495|Yellow||2008-12-03|2008-12-12|2015-10-12|Child: Graduated|Child: Graduated||82||1|1|1|1|M|Black||20|No|Mother|28217|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28226|Bachelors Degree|Married|Tech: Engineer|28202|2|8|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017777|501347335|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|34|2|||7446|3|||1|
502861544|502817316|500588737|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|318|Red||2011-12-22|2012-01-03|2012-11-16|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||10.4||1|1|1|1|M|Black||20|No|Mother|28205|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|Black||45|28210|Some College|Married|Tech: Production Line||8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502862935|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|4|||7496|10|||1|
500997812|501429055|500329285|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1404|Green||2008-12-30|2009-01-12|2012-11-16|Child/Family: Moved|Child/Family: Moved||46.1||1|1|1|1|M|Black||20|No|Mother|28266|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|M|White||40|28203|Bachelors Degree|Single|Transport: Pilot||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011746|500998085|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7496|10|||1|
502249063|502266549|500468039|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|136|Yellow||2010-08-30|2010-09-17|2011-01-31|Volunteer: Time constraint|Volunteer: Time constraint||4.5||1|1|1|1|M|White||19|No|Mother|28277|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||49|28277|Bachelors Degree|Married|Self-Employed, Entrepreneur|28277|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|502249494|1|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
500838847|501647679|500364921|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|724|Green||2009-05-21|2009-06-15|2011-06-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||23.8||2|2|1|1|M|Black||19|No|Mother|28278|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|M|Black||37|28226|||Finance: Accountant|28110|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|500839116|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501792675|501664548|500386328|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|721|Green||2009-09-21|2009-09-30|2011-09-21|Volunteer: Moved|Volunteer: Moved||23.7||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||31|19085|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501793030|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502590656|502578640|500538729|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|132|Red|Project Big, 2010-2012 OJJDP JJI|2011-05-26|2011-06-30|2011-11-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.3||1|1|1|1|F|Black||19|No|Mother|28213|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|RTBM|F|Black||34|28262|Bachelors Degree|Single|Medical: Nurse|28262|1|6|TV|Media|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502591168|31|0|2|31|0|2|7|2|500004641||4|3|500004640, 500005291|-2|500004640|-2|0|4|||130|1|||1|500004640, 500005291
502045254|502171015|500454926|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1949|Yellow||2010-05-28|2010-06-08|2015-10-09|Child: Graduated|Child: Graduated||64||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||27|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017777|502045664|31|0|2|31|0|2|10|2|-2||4|2||-2|500007920, 500011315, 500011316|-2|0|10|||7496|10|||1|
500186434|500338442|500088982|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1419|Green||2006-04-19|2006-04-23|2010-03-12|Volunteer: Time constraint|Volunteer: Time constraint||46.6||2|2|1|1|M|Black||19||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|White||37|28210|Bachelors Degree|Single|Journalist/Media|28217|0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500187978|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500771298|500953236|500206613|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1454|Yellow||2007-10-17|2007-11-02|2011-10-26|Volunteer: Time constraint|Volunteer: Time constraint||47.8||1|1|1|1|M|Black||19||Mother|28105|One Parent: Female|$35,000 to $39,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28110|||Finance: Banking||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500771566|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|34|2|||46|2|||1|
500191820|500191501|500044434|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2890|Red|Amachi|2005-09-30|2005-09-30|2013-08-29|Child: Lost interest|Child: Lost interest||94.9|Y|2|2|2|2|M|Black||19||Mother|28227||Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||72|28214||Married|Retired||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500191823|31|0|1|31|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500186963|500189733|500037847|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2017|Green|Amachi|2005-05-04|2005-05-04|2010-11-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||66.3||1|1|1|1|F|Black||19||Mother|28269|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||69|28216|Bachelors Degree|Single|Arts, Entertainment, Sports|28237|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500010355|500188165|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502860019|502873149|500596129|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|733|Green||2012-02-06|2012-02-22|2014-02-24|Volunteer: Time constraint|Volunteer: Time constraint||24.1||1|1|1|1|F|Hispanic||19|No|Mother|28213|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||36|28205|Bachelors Degree||Tech: Engineer|28204|1|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502861418|3|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502601023|502546883|500550809|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1807|Green|2010-2012 OJJDP JJI|2011-08-18|2011-08-31|2016-08-11|Child: Graduated|Child: Graduated||59.4||1|1|1|1|F|Black||19||Mother|28216|Two Parent|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||51|28277|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|502601540|31|0|2|1|0|2|10|2|-2||4|1|500005291|-2||-2|6854|8|||7464|9|||1|500005291
501390340|501869291|500421297|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|217|Green|Amachi|2009-12-14|2010-01-07|2010-08-12|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.1||2|2|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||38|28208|||Law: Lawyer||0|0|Self|Self|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500010355|501390617|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501390340|501386074|500328396|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|252|Green|Amachi|2008-12-19|2009-01-29|2009-10-08|Volunteer: Moved|Volunteer: Moved||8.3||2|2|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||37|28205||Divorced|Medical: Doctor, Provider|28025|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501390617|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501390336|501554452|500334574|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|634|Green|Amachi|2009-01-21|2009-01-29|2010-10-25|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||20.8||1|1|1|1|M|Black||19|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|RTBM|M|White||37|28203|Some College|Single|Construction|28203|8|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|501390617|31|0|1|1|0|1|7|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501498116|501289204|500309404|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|104|Green||2008-11-03|2008-11-04|2009-02-16|Child (or Parent): Other Reason|Child (or Parent): Other Reason||3.4||1|1|2|2|F|Black||19|No|Mother|28208|One Parent: Female|Unknown|||Y|Yes||Neighbor/Friend|General Community||Match Support|F|Black||32|28214|Some College|Single|Tech: Production Line||1|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001281|501498402|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|8|||46|2|||1|
501234604|501165150|500278984|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1506|Yellow||2008-07-23|2008-07-23|2012-09-06|Child: Severity of challenges|Child: Severity of challenges||49.5||1|1|1|1|F|Black||19|No|Mother|28215|Grandparents|Unknown||||No||Self|General Community||Match Support|F|Black||38|28213|Masters Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501234880|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
501561536|501651672|500361623|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|362|Red||2009-05-06|2009-05-15|2010-05-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.9||1|1|1|1|M|Black||19|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||33|28209|Bachelors Degree|Single|Finance: Banking|28204|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501561821|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502824908|502891382|500596373|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1247|Green||2012-02-06|2012-02-21|2015-07-22|Child: Graduated|Child: Graduated||41||1|1|1|1|F|Black||19|No|Mother|28226|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community||Match Support|F|White||34|28226|Bachelors Degree|Married|Unknown|29715|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502826191|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501015201|500953684|500208541|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1255|Yellow||2007-10-23|2007-11-13|2011-04-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||41.2||1|1|1|1|F|Black||19|No|Mother|28227|One Parent: Female|Less than $10,000||||No|AARTF|Neighbor/Friend|General Community||Enrollment|F|White||36|28211|Bachelors Degree|Single|Finance: Auditor||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011639|501015474|31|0|2|1|0|2|5|2|-2||4|2||-2||-2|6855|8|||46|2|||1|
500185907|500697782|500134557|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3034|Red|Amachi|2006-10-29|2006-10-29|2015-02-18|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||99.7||2|3|1|1|F|Black||19|Yes|Mother|28262|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||48|28212||Single|Medical: Healthcare Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500187470|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500514447|500807371|500174451|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|926|Red||2007-04-30|2007-04-30|2009-11-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||30.4||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|$20,000 to $24,999||||Yes||Neighbor/Friend|General Community||Match Support|M|White||44|28204|Bachelors Degree|Living w/ Significant Other|Finance: Banking||5|0|Superbowl 41|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500514698|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|8|||4178|1|||1|
500930976|501176751|500280106|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1717|Green||2008-07-31|2008-08-13|2013-04-26|Child: Lost interest|Child: Lost interest||56.4||1|1|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|||Y|No||Service Organization|General Community||Match Support|F|Black||66|28205|Masters Degree|Single|Self-Employed, Entrepreneur||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500931243|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|11|||46|2|||1|
500459684|500773055|500161728|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1134|Red||2007-02-20|2007-02-27|2010-04-06|Child/Family: Moved|Child/Family: Moved||37.3||1|1|2|2|M|Black||19|No|Mother|28211|One Parent: Female|Unknown||||No|Hampton Crest|Service Organization|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500459932|31|0|1|3|14|1|10|2|-2||4|3||-2||-2|7295|11|||46|2|||1|
502671406|502885637|500597397|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|933|Yellow||2012-02-09|2012-02-14|2014-09-04|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||30.7||1|1|1|1|F|Black||19|No|Mother|28210|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||34|28226|PHD|Single|Medical: Healthcare Worker|28207|3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502672234|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500898048|501141032|500248589|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|342|Green||2008-02-27|2008-03-07|2009-02-12|Child/Family: Time constraints|Child/Family: Time constraints||11.2||1|1|1|1|M|Black||19|No|Mother|28262|One Parent: Female|$30,000 to $34,999||||No||Relative|General Community||Match Support|M|Hispanic||37|28269||Single|Finance: Accountant|28164|0|0|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500001281|500898318|31|0|1|3|0|1|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
501741559|502213067|500464036|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|426|Yellow||2010-08-03|2010-08-13|2011-10-13|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||32|28208|Bachelors Degree|Married|Tech: Production Line||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|501741899|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501687515|501284245|500361402|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|558|Green||2009-05-05|2009-05-21|2010-11-30|Volunteer: Moved|Volunteer: Moved||18.3||1|1|1|1|M|White||19|No|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||36|28078|Bachelors Degree|Single|Tech: Support, Writing|28204|2|0|General|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501687853|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||6450|12|||1|
502893765|502874079|500599963|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1159|Green||2012-02-23|2012-03-08|2015-05-11|Child: Graduated|Child: Graduated||38.1||1|1|1|1|F|Black||19|No|Mother|28213|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||32|28262|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502895172|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502431164|502850528|500606503|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1291|Green||2012-03-27|2012-03-30|2015-10-12|Child: Graduated|Child: Graduated||42.4||1|1|1|1|M|Black||19|No|GrandMother|28208|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community||Match Support|M|White||59|28277|Masters Degree|Single|Tech: Computer/Programmer|28203|3|4|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502431607|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|5|||7439|1|||1|
500408135|500189709|500099932|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3172|Green|Amachi|2006-05-25|2006-05-25|2015-01-30|Child: Graduated|Child: Graduated||104.2||1|1|4|4|F|Black||19|Yes|Mother|28083|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500008321|500408385|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294, 500016374|-2|6854|8|||2230|7|||1|500000294
500360893|500382815|500091022|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1042|Green|Amachi|2006-04-28|2006-04-28|2009-03-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.2||1|1|1|1|M|Black||19|Yes|Mother|28210|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|M|Black||72|28222|Some College|Single|Business: Clerical|28203|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|RTBM|1|0|1|0|277|60|598|500000170|500003657|500361143|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294
501181241|502196362|500460441|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|98|Green|Amachi|2010-07-09|2010-07-20|2010-10-26|Child: Severity of challenges|Child: Severity of challenges||3.2||2|2|1|1|F|Black||19|Yes|GrandMother|28205|Two Parent|$25,000 to $29,999||||Yes||Self|General Community|Amachi|Match Support|F|White||45|28205|Masters Degree|Married|Retail: Mgt||2|0|Self|Self|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500003657|501181515|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501181241|501228929|500281828|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|675|Green|Amachi|2008-08-13|2008-08-22|2010-06-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||22.2||2|2|1|1|F|Black||19|Yes|GrandMother|28205|Two Parent|$25,000 to $29,999||||Yes||Self|General Community|Amachi|Match Support|F|White||35|28205|Bachelors Degree|Single|Business: Mgt, Admin|28211|0|9|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501181515|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||2238|7|||1|500000294
502765606|502842142|500607132|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|904|Red||2012-03-29|2012-04-03|2014-09-24|Volunteer: Moved|Volunteer: Moved||29.7||1|1|1|1|F|Black||19|No|Mother|28105|One Parent: Female|$15,000 to $19,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28209|Some College|Single|Finance: Accountant|28232|0|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502766519|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|6854|8|||7462|13|||1|
502011780|501828625|500516418|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|208|Green|2010-2012 OJJDP JJI|2011-02-09|2011-02-10|2011-09-06|Child: Lost interest|Child: Lost interest||6.8||2|2|2|2|F|White||19|No|Mother|28081|Two Parent|Unknown||||No||School|General Community|2010-2012 OJJDP JJI|Match Support|F|Asian||40|28027|Masters Degree|Married|Govt: Mgmt/Admin|28082|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|502012179|1|0|2|4|0|2|10|2|-2||4|1|500005291|-2||-2|0|4|||7464|9|||1|500005291
500186260|500189139|500037139|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4066|Yellow||2004-10-29|2004-10-29|2015-12-17|Child: Graduated|Child: Graduated||133.6||3|3|1|1|M|Black||19|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Site||Match Support|M|Black||42|28025|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500002335|500187857|31|0|1|31|0|1|10|2|-2||4|2||-1||-2|0|10|||7464|9|||1|
501603874|501671842|500355825|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|235|Green||2009-04-07|2009-04-09|2009-11-30|Volunteer: Time constraint|Volunteer: Time constraint||7.7||1|1|1|1|M|Black||19|No|Mother|28213|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||35|28202|||Business: Engineer|29715|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501604194|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
501299214|501186582|500283997|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|120|Red||2008-08-27|2008-09-22|2009-01-20|Child/Family: Moved|Child/Family: Moved||3.9||1|1|1|1|F|White||19|No|Father|28214|One Parent: Male|Unknown||||No||Therapist/Counselor|General Community||Match Support|F|White||60|28120|High School Graduate|Married|Law: Legal Secretary|28280|7|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500001267|501299492|1|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|5|||7446|3|||1|
501516900|501438601|500332399|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2402|Green||2009-01-13|2009-01-28|2015-08-27|Child: Graduated|Child: Graduated||78.9||1|1|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||39|28212|Bachelors Degree|Single|Medical: Healthcare Worker|28210|1|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|501517192|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|6854|8|||7462|13|||1|
501194371|501062230|500262721|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|647|Red||2008-04-24|2008-05-27|2010-03-05|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||21.3||2|2|1|1|F|Multi-race (Black & White)||19|No|Mother|28216|Two Parent|$15,000 to $19,999||||Yes||Therapist/Counselor|General Community||Match Support|F|Black||32|28216|Bachelors Degree|Single|Insurance||4|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501194645|36|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|5|||7446|3|||1|
501194371|502143351|500463829|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|41|Red||2010-08-02|2010-08-26|2010-10-06|Child: Lost interest|Child: Lost interest||1.3||2|2|2|2|F|Multi-race (Black & White)||19|No|Mother|28216|Two Parent|$15,000 to $19,999||||Yes||Therapist/Counselor|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Law|28273|5|0|Relative|Relative|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500009007|501194645|36|0|2|1|0|2|10|2|-2||4|3||-2|500000294|-2|0|5|||17161|11|||1|
501204263|500710082|500263390|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|262|Green||2008-04-28|2008-04-29|2009-01-16|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||8.6||1|1|2|2|M|White||19|No|Mother|28078|One Parent: Female|Unknown||||No|Radio|Media|General Community||Enrollment|M|White||51|28078||Single|Business: Sales||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501204537|1|0|1|1|0|1|5|2|-2||4|1||-2||-2|55|1|||46|2|||1|
501204266|501077703|500263389|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|694|Red||2008-04-28|2008-04-29|2010-03-24|Volunteer: Time constraint|Volunteer: Time constraint||22.8||1|1|1|1|F|White||19|No|Mother|28078|One Parent: Female|Unknown||||No|Radio|Media|General Community||Enrollment|F|White||31|28216|Bachelors Degree|Single|Business: Marketing||0|4|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501204540|1|0|2|1|0|2|5|2|-2||4|3||-2||-2|55|1|||46|2|||1|
500539341|500191356|500123020|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1951|Green|Amachi|2006-09-21|2006-09-24|2012-01-27|Child: Family structure changed|Child: Family structure changed||64.1||1|1|2|2|M|White||19|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||44|28205||Single|Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001281|500539592|1|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
500186960|500738970|500186719|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2207|Red|Amachi|2007-07-31|2007-07-31|2013-08-15|Volunteer: Time constraint|Volunteer: Time constraint||72.5||2|2|1|1|M|White||19|Yes|Mother|28227|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||40|28105|Some College|Married|Military|28112|11|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500188147|1|0|1|1|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|6854|8|||2238|7|||1|500000294
501224287|501343190|500298289|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1911|Red|Amachi|2008-10-13|2008-10-30|2014-01-23|Child: Lost interest|Child: Lost interest||62.8||1|1|1|1|M|Black||19|Yes|Mother|28270|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||43|28262|Bachelors Degree|Married|Customer Service|28211|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501224558|31|0|1|31|0|1|10|2|-2||4|3|500000294|-2|500000294|-2|5635|9|||2230|7|||1|500000294
501994951|502048623|500455478|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1556|Yellow||2010-06-03|2010-06-15|2014-09-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||51.1||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|Unknown||||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||36|28078||Single|Customer Service||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|501843047|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|7294|13|||7464|9|||1|
500417506|500640012|500136537|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1090|Green||2006-11-01|2006-11-03|2009-10-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.8||1|1|1|1|M|Multi-Race (None of the above)||19||Mother|28215|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community||RTBM|M|Black||58|28205||Separated|Business: Sales|28212|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|500417756|7|0|1|31|0|1|7|2|-2||4|1||-2||-2|0|5|||7464|9|||1|
502966254|502895517|500609631|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1048|Yellow||2012-04-12|2012-05-04|2015-03-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.4||1|1|1|1|F|Black||19|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|F|Black||48|28217|Bachelors Degree|Divorced|Medical: Admin|28232|11|5|Local TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|500784955|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7438|1|||1|
501852702|501637271|500458675|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|431|Red||2010-06-25|2010-06-25|2011-08-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.2||1|1|1|1|F|Black||19|No|Mother|28216|Two Parent|Unknown||||No||Self|General Community||Match Support|F|White||33|28205||Single|Consultant|28205|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501853073|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500915359|501189280|500311316|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1094|Green||2008-11-06|2008-11-10|2011-11-09|Volunteer: Time constraint|Volunteer: Time constraint||35.9||3|3|1|1|F|Black||19|No|Mother|28227|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|F|White||38|28105|PHD|Married|Human Services: Non-Profit|28110|0|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500915629|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
500915359|503044413|500622861|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|860|Yellow||2012-07-05|2012-08-10|2014-12-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.3||3|3|1|1|F|Black||19|No|Mother|28227|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28204|Bachelors Degree|Single|Medical: Nurse||0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|500915629|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|34|2|||7496|10|||1|
502426852|502437756|500525086|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|373|Yellow||2011-03-14|2011-03-22|2012-03-29|Child/Family: Time constraints|Child/Family: Time constraints||12.3||1|1|1|1|F|Black||19|No|Mother|28278|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||61|28215|Bachelors Degree|Divorced|Self-Employed, Entrepreneur||0|0|TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502427295|31|0|2|31|0|2|10|2|-2||4|2|500000294|-2||-2|0|10|||130|1|||1|
502241349|502240986|500461089|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1140|Green||2010-07-15|2010-07-22|2013-09-04|Child/Family: Moved|Child/Family: Moved||37.5||1|1|2|2|M|Black||19|No|Aunt|28081|Two Parent|Unknown||||No|Other|Faith Organization|General Community||Match Support|M|Black||54|28025||Married|Clergy|28025|23|0|Other|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500002335|502241780|31|0|1|31|0|1|10|2|-2||4|1||-2|500016374|-2|5635|9|||7671|13|||1|
502714405|502764673|500577475|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1337|Green||2011-11-11|2011-12-08|2015-08-06|Child: Graduated|Child: Graduated||43.9||1|1|1|1|M|Black||19|No|Mother|28206|One Parent: Female|Less than $10,000|||Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||33|28213|Associate Degree|Single|Transport: Driver|28205|5|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500017732|502715293|31|0|1|31|0|1|10|2|-2||4|1|500005291|-2||-2|56|1|||7446|3|||1|
502142129|502926748|500605216|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|413|Red||2012-03-20|2012-04-04|2013-05-22|Volunteer: Time constraint|Volunteer: Time constraint||13.6||1|1|1|1|F|Some Other Race||19|No|Father|28214|One Parent: Male|Unknown||||No||Self|General Community||Match Support|F|White||45|28209|Bachelors Degree|Single|Tech: Engineer|2494|14|0||Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502142558|41|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||0|11|||1|
500191327|500547393|500144146|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2099|Green||2006-11-29|2006-12-07|2012-09-05|Child: Family structure changed|Child: Family structure changed||69||2|2|1|1|M|Black||19||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||42|28212||Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500191330|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502136043|502459922|500517447|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|836|Green|2010-2012 OJJDP JJI|2011-02-14|2011-02-21|2013-06-06|Child/Family: Moved|Child/Family: Moved||27.5||1|1|2|2|M|Black||19|No|GrandMother|28227|Other Relative|Unknown||||Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502136472|31|0|1|1|0|1|10|2|-2||4|1|500005291|-2|500004640|-2|56|1|||7464|9|||1|500005291
500740293|500876177|500179697|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2586|Yellow||2007-06-11|2007-06-12|2014-07-11|Child: Lost interest|Child: Lost interest||85||1|1|1|1|M|Black||19||Mother|28216|One Parent: Female|$20,000 to $24,999||||No||Therapist/Counselor|General Community||Match Support|M|Black||39|28216||Single|Transport: Pilot||3|0|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500740560|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|5|||6450|12|||1|
501349143|501637748|500363970|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|148|Yellow||2009-05-15|2009-05-27|2009-10-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.9||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||||Yes||Relative|General Community||RTBM|M|White||26|28031|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501349422|31|0|1|1|0|1|7|2|-2||4|2||-2||-2|0|3|||7464|9|||1|
500577810|500648158|500154518|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1359|Red||2007-01-24|2007-02-05|2010-10-26|Volunteer: Moved|Volunteer: Moved||44.6||1|1|1|1|F|Black||19||Mother|28273|One Parent: Female|$30,000 to $34,999||||No|BBBS National Site|Web Link|General Community||Match Support|F|Black||36|28273|Bachelors Degree|Single|Tech: Sales, Mktg|28608|1|6|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500578062|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|34|2|||6450|12|||1|
501285234|501463291|500329314|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|686|Yellow||2008-12-30|2009-01-13|2010-11-30|Volunteer: Time constraint|Volunteer: Time constraint||22.5||1|1|1|1|M|Multi-race (Black & Hispanic)||19|No|Mother|28269|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|White||32|28262|Bachelors Degree|Single|Service: Restaurant|28025|0|1|Recruitment Event|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|501285512|38|0|1|1|0|1|10|2|-2||4|2||-2|500000294|-2|0|8|||7460|12|||1|
503158441|503130365|500631432|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|657|Red||2012-08-29|2012-09-14|2014-07-03|Volunteer: Moved|Volunteer: Moved||21.6||1|1|1|1|F|Black||19|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||27|28202|Bachelors Degree|Single|Business||1|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|503160119|31|0|2|1|0|2|10|2|-2||4|3||-2|500000294|-2|0|5|||7464|9|||1|
501609864|501611087|500351248|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|255|Green||2009-03-23|2009-03-23|2009-12-03|Volunteer: Time constraint|Volunteer: Time constraint||8.4||1|1|1|1|M|Black||19|No||28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||30|28262|Bachelors Degree|Single|Finance: Banking|28262|0|7|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501610184|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7438|1|||1|
501209692|501267614|500278985|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|623|Red||2008-07-23|2008-07-23|2010-04-07|Volunteer: Time constraint|Volunteer: Time constraint||20.5||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||||Yes|Brochure|Media|General Community||Enrollment|M|Black||39|28209|Masters Degree|Married|Finance: Banking|28288|0|2||Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501209966|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|51|1|||0|11|||1|
501092911|501176101|500261235|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2665|Red||2008-04-16|2008-05-01|2015-08-18|Child: Graduated|Child: Graduated||87.6||1|1|1|1|M|Black||19||Mother|28226|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|White||37|28210|Some College|Single|Business: Mgt, Admin||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501064244|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|4|||46|2|||1|
500399525|500416787|500099891|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2267|Green||2006-05-25|2006-06-15|2012-08-29|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||74.5||1|1|1|1|F|Black||19||Mother|28214|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|Black||46|28217|Some College|Single|Finance: Accountant|28208|0|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500399775|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
502697677|502590370|500550704|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|572|Yellow||2011-08-18|2011-09-02|2013-03-27|Volunteer: Moved|Volunteer: Moved||18.8||1|1|1|1|F|Hispanic||19|No|Mother|28027|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|White||32|28027|Bachelors Degree|Single|Business: Marketing|28075|3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502605848|3|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501488008|501580288|500349241|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|120|Green||2009-03-12|2009-03-25|2009-07-23|Volunteer: Moved|Volunteer: Moved||3.9||1|1|1|1|F|Black||19|No|Mother|28213|One Parent: Female|Unknown||||Yes||Service Organization|General Community||Match Support|F|Some Other Race||39|28203|Masters Degree|Single|Business: Marketing|27101|2|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501488294|31|0|2|41|0|2|10|2|-2||4|1||-2||-2|0|11|||7464|9|||1|
501228477|501317923|500286344|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1009|Green||2008-09-05|2008-09-11|2011-06-17|Child/Family: Moved|Child/Family: Moved||33.1||1|1|1|1|M|Black||19|No|Mother|28105|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|M|White||59|28227|Some College|Married|Insurance|28211|0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501228753|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
500636603|500842825|500168014|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1549|Red||2007-03-21|2007-03-21|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||50.9||2|4|1|1|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|F|White||38|28226|Bachelors Degree|Married|Homemaker||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500636863|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|8|||7671|13|||1|
500186784|500909789|500184677|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1031|Green|Amachi|2007-07-17|2007-07-24|2010-05-20|Volunteer: Time constraint|Volunteer: Time constraint||33.9||2|2|1|1|F|Black||19|Yes|GrandMother|28205|Other Relative|Unknown|||Y|No||Self|General Community|Amachi|Enrollment|F|Black||33|28262|Bachelors Degree|Single|Education: Teacher||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500010355|500188096|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501765404|501958658|500443642|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1227|Yellow||2010-03-25|2010-04-20|2013-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||40.3||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Multi-race (Black & White)||28|28262||Single|Student: College|28262|3|0|UNCC|College Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501765751|31|0|1|36|0|1|10|2|-2||4|2||-2||-2|0|10|||9221|5|||1|
501190091|501262221|500289240|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|109|Green||2008-09-18|2008-09-29|2009-01-16|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.6||1|1|1|1|F|Black||19||Aunt|28215|Two Mothers|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|F|Black||38|28215||Married|Business: Clerical|28202|0|0||Relative|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008062|501190365|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|34|2|||0|11|||1|
501189685|501263133|500289237|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|109|Green||2008-09-18|2008-09-29|2009-01-16|Vol: Does Not Like Child or Parent|Vol: Does Not Like Child or Parent||3.6||1|1|1|1|M|Black||19|No|Aunt|28215|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|M|Black||35|28215|Masters Degree|Married|Tech: Engineer|28204|0|2||Relative|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500008062|501190365|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|3|||0|11|||1|
500799303|500798390|500167062|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3433|Red||2007-03-15|2007-03-27|2016-08-19|Child: Graduated|Child: Graduated||112.8||1|1|1|1|M|White||19|No|Mother|28081|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||46|28202||Single|Business: Sales||0|4|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500020753|500799571|1|0|1|1|0|1|10|2|-2||4|3|500016374|-2|500016374|-2|34|2|||7464|9|||1|
500186905|500189677|500037790|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3919|Red|Amachi|2005-02-10|2005-02-10|2015-11-04|Child: Graduated|Child: Graduated||128.8||1|1|1|1|F|Black||19|Yes|Mother|28205|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Match Support|F|Black||50|28215|Some College|Single|Finance: Banking||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500188151|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||7453|7|||1|500000294
501300101|500346193|500281421|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2461|Yellow|Amachi|2008-08-11|2008-08-14|2015-05-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||80.9||1|1|4|4|F|Black||19|Yes|GrandMother|28273|Grandparents|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||46|28278|Masters Degree|Single|Education: Teacher|28278|7|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501300379|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2||-2|7294|13|||46|2|||1|500000294
502063943|502890782|500617038|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|133|Red||2012-05-30|2012-06-20|2012-10-31|Child: Severity of challenges|Child: Severity of challenges||4.4||1|1|1|1|M|White||19|No|Mother|28213|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community||Match Support|M|White||62|28209|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Local Print|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502064367|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|5|||7439|1|1209|1|1|
500876118|500867392|500176228|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1163|Red||2007-05-09|2007-05-16|2010-07-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38.2||1|1|1|1|F|Black||19|No|Mother|28203|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||38|28207||Married|Business: Sales||2|0|Recruitment Event|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500876387|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7460|12|||1|
501776333|501832599|500381636|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1416|Green||2009-08-31|2009-09-08|2013-07-25|Volunteer: Moved|Volunteer: Moved||46.5||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||39|28210|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011746|501776688|31|0|1|31|0|1|10|2|-2||4|1||-2|500000294|-2|34|2|||7464|9|||1|
501124034|501543908|500337028|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|222|Green||2009-01-29|2009-02-19|2009-09-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.3||2|2|1|1|F|Black||19|No|Mother|28269|One Parent: Female|Less than $10,000||||Yes||Therapist/Counselor|General Community||Match Support|F|Black||33|28269|Bachelors Degree|Single|Tech: Research/Design|28285|0|5|Local Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009242|501124308|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|5|||7437|1|||1|
500465790|500398217|500153025|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Green||2007-01-18|2007-01-23|2009-06-23|Child/Family: Infraction of match rules/agency policies Volunteer: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies|29||1|1|2|2|M|Black||19||Mother|28212|One Parent: Female|Unknown||||No|Brochure|Media|General Community||Match Support|M|Black||56|28213|Bachelors Degree|Single|Finance: Banking||0|6|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500466041|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|51|1|||7458|9|||1|
501714939|501584958|500365824|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1299|Yellow|Amachi|2009-05-27|2009-06-03|2012-12-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||42.7||1|1|1|1|M|Black||19|Yes|Mother|28105|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||34|28277||Single|Business: Sales|28206|0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|501715277|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
500733695|500307108|500150172|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2989|Red|Amachi|2006-12-26|2006-12-26|2015-03-03|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||98.2||1|1|1|1|F|Black||19|Yes|GrandMother|28217|Grandparents|Less than $10,000|||Y|No|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||34|28210|Bachelors Degree|Married|Finance: Accountant|28202|0|2|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|500733962|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2||-2|7294|13|||2238|7|||1|500000294
501097437|500967534|500241097|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|345|Green||2008-01-30|2008-02-06|2009-01-16|Child: Severity of challenges Vol: Other Reason|Child: Severity of challenges|Vol: Other Reason|11.3||1|1|1|1|F|White||19|No|GrandMother|28078|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||46|28078|Some College|Married|Business: Mgt, Admin|28202|5|6|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500001281|501097711|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501431685|501556970|500338061|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|779|Green|Amachi|2009-02-03|2009-02-10|2011-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25.6||1|1|1|1|M|Black||19|Yes|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||35|28215|High School Graduate|Married|Service: Restaurant|28105|0|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501431970|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501572942|500981458|500349208|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|80|Green||2009-03-12|2009-05-01|2009-07-20|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||2.6||1|1|2|2|F|Black||19|No|Foster Parent|28027|Foster Home|Unknown||||Yes||Self|General Community||Match Support|F|Black||40|28075|Masters Degree|Married|Finance: Banking||8|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001262|501012375|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||2238|7|||1|
501309737|501347994|500302521|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|109|Green|Amachi|2008-10-21|2008-10-31|2009-02-17|Volunteer: Changed workplace/school partnership Child/Family: Moved|Volunteer: Changed workplace/school partnership|Child/Family: Moved|3.6||2|2|1|1|F|Black||19|Yes|Mother|28208|One Parent: Female|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Enrollment|F|Black||37|28269|Some College|Married|Human Services: Social Worker|28269|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500007521|501310015|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2||-2|7294|13|||7464|9|||1|500000294
501309737|501289204|500359681|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|516|Green|Amachi|2009-04-27|2009-05-01|2010-09-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||17||2|2|2|2|F|Black||19|Yes|Mother|28208|One Parent: Female|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Enrollment|F|Black||32|28214|Some College|Single|Tech: Production Line||1|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501310015|31|0|2|31|0|2|5|2|-2||4|1|500000294|-2|500000294|-2|7294|13|||46|2|||1|500000294
501073858|501184292|500255133|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|859|Green|Amachi|2008-03-26|2008-03-27|2010-08-03|Volunteer: Moved|Volunteer: Moved||28.2||1|1|1|1|M|Black||19|Yes|Mother|28205|One Parent: Female|Less than $10,000||||Yes||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||33|28203|Bachelors Degree|Single|Finance: Banking|28255|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501074131|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|8|||46|2|||1|500000294
502316483|502428948|500518256|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|580|Yellow|Project Big AND Amachi|2011-02-17|2011-02-25|2012-09-27|Child: Lost interest|Child: Lost interest||19.1||1|1|1|1|M|Black||19|Yes|Mother|28208|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|M|Black||32|28269|Bachelors Degree|Single|Medical: Pharmacist|27511|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011746|501467438|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|4|||7496|10|||1|500004901
500185723|501310677|500284133|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2484|Red||2008-08-27|2008-09-05|2015-06-25|Child: Graduated|Child: Graduated||81.6||2|2|1|1|M|Black||19||Mother|28214|One Parent: Female|Unknown||||No|AARTF|Neighbor/Friend|General Community||Match Support|M|Black||36|28214|Bachelors Degree|Single|Tech: Computer/Programmer|28147|0|3|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500187335|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|6855|8|||7464|9|||1|
501872495|501891059|500418064|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|316|Red||2009-12-03|2009-12-14|2010-10-26|Child/Family: Moved|Child/Family: Moved||10.4||1|1|1|1|M|Black||19|No|Non-Relative: Other|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|Some Other Race||37|28209|PHD|Single|Medical: Doctor, Provider||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501872868|31|0|1|41|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501342393|501210017|500293459|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2053|Green||2008-09-30|2008-10-22|2014-06-06|Child: Lost interest|Child: Lost interest||67.4||1|1|1|1|F|White||19|No|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||31|28209|Bachelors Degree|Single|Business: Sales||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500017732|501342672|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501064559|501479598|500344055|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|111|Green||2009-02-23|2009-02-25|2009-06-16|Child (or Parent): Other Reason|Child (or Parent): Other Reason||3.6||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|$40,000 to $44,999||||Yes||Neighbor/Friend|General Community||Match Support|M|White||34|28269|Bachelors Degree|Married|Finance: Accountant|28202|3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501064832|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
502072733|502080569|500456384|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|79|Green||2010-06-10|2010-06-15|2010-09-02|Child: Lost interest|Child: Lost interest||2.6||1|1|2|2|F|Black||19|No|GrandMother|28216|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||33|28078|High School Graduate|Single|Self-Employed, Entrepreneur|28269|0|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|502073157|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502926905|503096831|500635818|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|687|Yellow||2012-09-17|2012-10-31|2014-09-18|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||22.6||1|1|1|1|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||32|28216|Bachelors Degree|Single|Tech: Support, Writing|28117|1|9|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502928325|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|7294|13|||7438|1|||1|
501060196|501036081|500223215|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2807|Green||2007-11-26|2007-11-26|2015-08-03|Child/Family: Moved|Child/Family: Moved||92.2||1|1|1|1|M|Black||19|No|Mother|28205|One Parent: Female|$15,000 to $19,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28226|Masters Degree|Single|Finance: Accountant||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500011349|501060469|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
501214257|501075530|500258621|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|578|Green||2008-04-11|2008-04-11|2009-11-10|Volunteer: Time constraint|Volunteer: Time constraint||19||1|1|1|1|F|Black||19|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|White||37|28207|Bachelors Degree|Married|Business: Marketing||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501214533|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500923444|500824500|500182563|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|988|Green|Amachi|2007-06-29|2007-08-13|2010-04-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||32.5|Y|1|1|1|1|M|Black||19|No|Mother|28083|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|RTBM|F|Black||51|28027||Married|Medical: Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500002335|500923714|31|0|1|31|0|2|7|2|500003586||4|1|500005291|-2|500000294|-2|5635|9|||2238|7|||1|500000294
501614044|501315493|500349169|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|837|Yellow||2009-03-12|2009-04-06|2011-07-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27.5||1|1|1|1|F|Hispanic||19|No|Mother|28273|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||41|28273|Bachelors Degree|Single|Tech: Research/Design|28217|0|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501614360|3|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502173445|502266833|500532710|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|857|Red|Amachi|2011-04-21|2011-05-23|2013-09-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.2||1|1|1|1|F|Black||19|Yes|Mother|28214|One Parent: Female|Unknown||||Yes||Service Organization|General Community|Amachi|Match Support|F|White||28|28206|Bachelors Degree|Single|Education: Teacher||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502173869|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2||-2|0|11|||7464|9|||1|500000294
502743091|503079983|500623169|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|778|Yellow||2012-07-09|2012-07-18|2014-09-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25.6||1|1|1|1|M|Black||19|No|Mother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||39|28203|Bachelors Degree|Single|Unemployed||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502743998|31|0|1|1|0|1|10|2|-2||4|2|500005291|-2||-2|6854|8|||7496|10|||1|
501401872|501721615|500433383|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|239|Green||2010-02-09|2010-05-05|2010-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.9||2|2|2|2|M|Black||19|No|Mother|28215|One Parent: Female|Unknown||||Yes||Service Organization|General Community||Enrollment|M|Hispanic||47|28215||Married|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501402157|31|0|1|3|0|1|5|2|-2||4|1||-2||-2|0|11|||46|2|||1|
501401872|500783871|500323014|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|336|Green||2008-12-04|2008-12-10|2009-11-11|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11||2|2|2|2|M|Black||19|No|Mother|28215|One Parent: Female|Unknown||||Yes||Service Organization|General Community||Enrollment|M|Black||42|28205|||Education: Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|501402157|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|11|||46|2|||1|
501791428|501726049|500374912|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1135|Green||2009-07-21|2009-07-29|2012-09-06|Volunteer: Moved|Volunteer: Moved||37.3||1|1|1|1|M|Black||19|No|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Multi-Race (None of the above)||33|28273|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501163776|31|0|1|7|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500881720|501165156|500260861|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1158|Green||2008-04-15|2008-04-15|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38||1|1|1|1|M|Black||19|No|Mother|28269|One Parent: Female|$10,000 to $14,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|Black||33|28269|Bachelors Degree|Single|Finance: Banking||0|5|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500881989|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
501330628|501245666|500287591|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|913|Green|Amachi|2008-09-11|2008-09-29|2011-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||30||1|1|2|2|F|Black||19|Yes|Mother|28208|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||33|28215|Bachelors Degree|Single|Tech: Support, Writing|28204|6|0|Other|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|1|0|1|0|277|60|598|500000170|500003657|501330906|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500014506|-2|34|2|||7671|13|||1|500000294
502217445|502685222|500573483|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|352|Red||2011-11-02|2011-11-14|2012-10-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.6||1|1|1|1|M|Black||19|No|Mother|28226|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||42|28277|Some College|Single|Self-Employed, Entrepreneur||5|0|Local Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502217876|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7437|1|||1|
500968246|501179573|500251681|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2557|Green||2008-03-11|2008-04-29|2015-04-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||84||1|1|1|1|M|Black||19|No|Aunt|28269|One Parent: Female|$10,000 to $14,999|||Y|No||Therapist/Counselor|General Community||Match Support|M|Black||35|28213|Bachelors Degree|Single|Business: Sales||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500968516|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|5|||46|2|||1|
500185571|500188438|500089543|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3360|Red||2006-04-25|2006-05-02|2015-07-14|Child: Graduated|Child: Graduated||110.4||1|1|1|1|M|Black||19||Mother|28215|Other/Unknown|Unknown||||No|Other|Faith Organization|General Community||Match Support|M|Black||49|28213|Bachelors Degree|Married|Finance: Banking|28288|4|6|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500187198|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|5635|9|||7464|9|||1|
502527850|502598777|500541242|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|462|Yellow|2010-2012 OJJDP JJI|2011-06-15|2011-06-30|2012-10-04|Child: Lost interest|Child: Lost interest||15.2||1|1|2|2|F|Black||19|No|Mother|28027|One Parent: Female|Less than $10,000||||Yes|Brochure|Media|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||42|28213|Bachelors Degree|Single|Finance: Banking|28202|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|502528298|31|0|2|31|0|2|10|2|-2||4|2|500005291|-2|500016374|-2|51|1|||7464|9|||1|500005291
500969479|500955544|500274110|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|379|Red||2008-06-19|2008-07-22|2009-08-05|Volunteer: Time constraint|Volunteer: Time constraint||12.5||1|1|1|1|F|Black||19|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|No||Therapist/Counselor|General Community||Enrollment|F|Black||47|28217|Bachelors Degree||Education: Teacher||3|0|Essence Magazine|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500969749|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|5|||3892|1|||1|
501146326|501247637|500269664|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|689|Green||2008-06-03|2008-06-17|2010-05-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||22.6||1|1|1|1|M|Black||19||Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||32|28269|Bachelors Degree|Married|Finance: Banking|28262|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501146600|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500186282|500189220|500037220|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1710|Green||2005-08-10|2005-08-10|2010-04-16|Volunteer: Time constraint|Volunteer: Time constraint||56.2||1|1|1|1|F|Black||19||Mother|28227|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|Black||38|28078|Bachelors Degree||Medical: Healthcare Worker||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500187881|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500185806|501043306|500262116|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1094|Yellow||2008-04-22|2008-04-22|2011-04-21|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||35.9||4|4|1|1|F|Black||19||Mother|28203|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|Black||40|28211|Masters Degree|Single|Finance: Banking||0|3|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500009007|500187395|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
500185865|500189140|500326656|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2074|Yellow||2008-12-15|2008-12-15|2014-08-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||68.1||2|2|2|2|F|Black||19||Mother|28213|Other/Unknown|Unknown||||No||Self|General Community||Match Support|F|Black||40|28273|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|500187761|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501641322|501400426|500366881|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|118|Green||2009-06-01|2009-06-24|2009-10-20|Volunteer: Time constraint|Volunteer: Time constraint||3.9||2|2|1|1|F|Black||19||Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Hispanic||37|28262|Bachelors Degree|Divorced|Journalist/Media|28262|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501641645|31|0|2|3|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501641322|500892262|500419238|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|117|Red|Amachi|2009-12-08|2010-01-15|2010-05-12|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||3.8||2|2|2|2|F|Black||19||Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black|Other African|36|28105||Single|Consultant|28244|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501641645|31|0|2|31|31|2|10|2|||4|3||-2||-2|0|10|||46|2|||1|500000294
501641337|500835981|500373972|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2044|Green||2009-07-14|2009-08-07|2015-03-13|Volunteer: Moved|Volunteer: Moved||67.2||1|1|2|2|F|Black||19|No|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||31|28269|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500011349|501641648|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2|500000294|-2|0|10|||46|2|||1|
501226826|501293480|500310244|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1056|Red|Amachi|2008-11-04|2008-11-07|2011-09-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.7||1|1|1|1|M|Black||19|Yes|Mother|28215|One Parent: Female|Unknown||||Yes||Relative|General Community|Amachi|Match Support|M|White||33|28202|Masters Degree|Single|Finance: Economist||0|8|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501227093|31|0|1|1|0|1|10|2|-2||4|3|500000294|-2||-2|0|3|||7447|3|||1|500000294
501365520|500868727|500454745|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|427|Green||2010-05-27|2010-05-28|2011-07-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||14||1|1|4|4|F|Black||19||Mother|28203|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||38|28214|Bachelors Degree|Single|Business: Clerical|28273|2|3|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|501365799|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
501506214|501588885|500351462|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2644|Green||2009-03-23|2009-03-28|2016-06-23|Child: Graduated|Child: Graduated||86.9||1|1|1|1|M|Black||19|No|Mother|28105|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||55|28173|||Unknown|28203|0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|501506506|31|0|1|31|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
502526973|503037794|500623286|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|217|Green||2012-07-09|2012-07-19|2013-02-21|Volunteer: Moved|Volunteer: Moved||7.1||1|1|1|1|M|Hispanic||19|No|Mother|28210|One Parent: Female|Less than $10,000||||Yes||Relative|General Community||Match Support|M|Hispanic||27|28202|Bachelors Degree|Single|Finance|28255|0|11|Coworker|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502527426|3|0|1|3|0|1|10|2|-2||4|1||-2||-2|0|3|||7447|3|||1|
500186570|500189615|500037719|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|2373|Yellow||2004-10-05|2004-10-05|2011-04-05|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||78||2|2|1|1|F|Black||19||Mother|28269|Other/Unknown|Unknown||||No||Self|General Community||RTBM|F|Black||37|28213|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500188168|31|0|2|31|0|2|7|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
501313839|501788563|500396680|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1315|Yellow||2009-10-19|2009-11-11|2013-06-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||43.2||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||36|28204|Bachelors Degree|Single|Consultant||4|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|501314117|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500186768|500189734|500037848|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1643|Yellow|Amachi|2005-04-07|2005-04-07|2009-10-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||54||2|2|1|1|M|Black||19||Mother|28213|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||39|28202|Bachelors Degree|Single|Business: Sales|28262|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500188084|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501645192|501519306|500374818|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2586|Red||2009-07-21|2009-07-21|2016-08-19|Child: Graduated|Child: Graduated||85||1|1|2|2|M|Hispanic||19|No|Mother|28025|One Parent: Female|Unknown||||Yes||Self|General Community|Cabarrus County|Match Support|M|White||63|28075||Married|Unknown||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500020753|501645515|3|0|1|1|0|1|10|2|-2||4|3|500016374|-2|500016374|-2|0|10|||7464|9|||1|
500796688|500578813|500155138|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|742|Green|Amachi|2007-01-28|2007-02-05|2009-02-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.4||1|1|1|1|M|Black||19|Yes|Mother|28216|Other/Unknown|Unknown||||No||Self|General Community|Amachi|RTBM|M|Black||49|28204||Single|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188072|31|0|1|31|0|1|7|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502205848|502624702|500549350|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2037|Green|2010-2012 OJJDP JJI|2011-08-10|2011-08-18|NaT||||66.9||1|1|1|1|M|Black||19|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Juris Doctorate (JD)|Single|Student: College|28208|0|0||Law Student Association|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502206277|31|0|1|1|0|1|10|2|-2||2|1|500005291|-2||-2|0|10|||0|15|||1|500005291
500186990|500189496|500339895|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1837|Red|Amachi|2009-02-10|2009-02-17|2014-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||60.4||2|2|3|3|M|Black||19|Yes|Mother|28269|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||51|28269|Bachelors Degree|Married|Unknown|28202|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|500188170|31|0|1|31|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501868921|501220647|500398441|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|417|Yellow||2009-10-22|2009-10-30|2010-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.7||2|2|1|1|F|Black||19|No|Mother|28211|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||34|28217|Juris Doctorate (JD)|Married|Law: Lawyer|28204|0|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501869291|31|0|2|31|0|2|10|2|-2||4|2|500005291|-2||-2|0|10|||7464|9|||1|
501868921|501382633|500524206|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1947|Green|2010-2012 OJJDP JJI|2011-03-09|2011-03-31|2016-07-29|Child/Family: Moved|Child/Family: Moved||64||2|2|2|2|F|Black||19|No|Mother|28211|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28211||Married|Finance: Banking|28255|0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501869291|31|0|2|1|0|2|10|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|500005291
502537477|500189507|500535475|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1890|Green|Project Big, 2010-2012 OJJDP JJI|2011-05-09|2011-05-12|2016-07-14|Child: Graduated|Child: Graduated||62.1||1|1|3|4|F|Black||19||Mother|28208|Two Parent|$15,000 to $19,999||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||48|28214|Bachelors Degree|Single|Tech: Management|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Project Big|Enrollment|0|1|0|1|277|60|598|500000170|500017732|502537922|31|0|2|31|0|2|10|2|-2||4|1|500004640, 500005291|-2|500000294, 500004640|-2|0|4|||2238|7|||1|500004640, 500005291
500911250|500911214|500183000|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|595|Green|Amachi|2007-07-05|2007-07-19|2009-03-05|Child/Family: Moved|Child/Family: Moved||19.5||1|1|1|1|F|Black||19|Yes|Mother|28075|One Parent: Female|$15,000 to $19,999|||Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||75|28212||Widowed|Business: Clerical||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|RTBM|1|0|1|0|277|60|598|500000170|500003657|500911515|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||7453|7|||1|500000294
501877268|501942543|500429020|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|625|Red||2010-01-22|2010-01-26|2011-10-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.5||1|1|1|1|M|Black||19|No|Mother|28213|One Parent: Female|Unknown|||Y|Yes|Radio|Media|General Community||Match Support|M|White||33|28269|||Construction||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|501877641|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|55|1|||7447|3|||1|
501669649|501818546|500388262|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|887|Red||2009-09-25|2009-10-26|2012-03-31|Volunteer: Time constraint|Volunteer: Time constraint||29.1||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Enrollment|M|Black||67|28262||Married|Business: Mgt, Admin||32|0|Mayfield Memorial|Faith Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013709|501669987|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|6854|8|||9212|7|||1|
501184645|500781896|500245777|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1260|Green||2008-02-18|2008-02-22|2011-08-05|Volunteer: Moved|Volunteer: Moved||41.4||1|1|2|2|M|Multi-race (Black & White)||19|No|Mother|28081|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||37|28027|Bachelors Degree|Married|Business: Sales|27263|4|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501184919|36|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501631547|502170945|500528464|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1947|Green|Project Big, 2010-2012 OJJDP JJI|2011-03-30|2011-03-31|2016-07-29|Child: Graduated|Child: Graduated||64||2|2|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||38|28277|Bachelors Degree|Single|Arts, Entertainment, Sports|28203|3|6|UnitedMethodistChrch|Faith Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501631870|31|0|1|1|0|1|10|2|500004641||4|1|500004640, 500005291|-2||-2|0|10|||8529|7|||1|500004640, 500005291
501631547|501645587|500388261|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|447|Yellow|Project Big|2009-09-25|2009-09-30|2010-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.7||2|2|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||32|28202|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501631870|31|0|1|1|0|1|10|2|500004641||4|2|500004640, 500005291|-2||-2|0|10|||7464|9|||1|500004640
500871683|500933829|500199601|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3066|Green|Amachi|2007-10-01|2007-10-01|2016-02-22|Child: Graduated|Child: Graduated||100.7||1|1|1|1|M|Black||19|Yes|Aunt|28208|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Match Support|M|White||46|28209|Masters Degree|Single|Self-Employed, Entrepreneur|28209|4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500871952|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501572413|501528066|500348882|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|742|Green|Amachi|2009-03-11|2009-03-25|2011-04-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.4||1|1|1|1|M|Black||19|Yes|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|M|White||46|28269|Bachelors Degree|Living w/ Significant Other|Medical: Nurse|28232|1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501572709|31|0|1|1|0|1|5|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
502265907|501332017|500512367|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|387|Red|Amachi|2011-01-21|2011-01-31|2012-02-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.7||1|1|1|1|F|Black||19|Yes|Mother|28210|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||37|28209|PHD|Single|Medical: Doctor, Provider|28210|2|3|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|502266339|31|0|2|1|0|2|10|2|-2||4|3|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501724491|501852487|500397005|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|517|Green||2009-10-20|2009-10-29|2011-03-30|Volunteer: Moved|Volunteer: Moved||17||1|1|1|1|M|Multi-race (Black & Asian)||19|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||42|28216||Divorced|Medical|28078|1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501724831|39|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501811385|502460013|500524684|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1976|Red|2010-2012 OJJDP JJI, Cabarrus County|2011-03-11|2011-03-23|2016-08-19|Child: Graduated|Child: Graduated||64.9||2|2|1|1|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||43|28075|Bachelors Degree|Married|Business: Mgt, Admin||7|0|Recruitment Event|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500020753|501811730|31|0|2|31|0|2|10|2|-2||4|3|500016374|-2|500016374|-2|6854|8|||7459|10|||1|500005291, 500016374
501811385|500981458|500374643|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|589|Green||2009-07-20|2009-07-27|2011-03-08|Volunteer: Time constraint|Volunteer: Time constraint||19.4||2|2|2|2|F|Black||19|No|Mother|28027|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||40|28075|Masters Degree|Married|Finance: Banking||8|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002335|501811730|31|0|2|31|0|2|10|2|-2||4|1|500016374|-2|500000294|-2|6854|8|||2238|7|||1|
501394968|501322428|500310512|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|859|Green||2008-11-05|2008-11-21|2011-03-30|Volunteer: Moved|Volunteer: Moved||28.2||1|1|1|1|M|Black||19|No|Mother|28278|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||44|28277|Masters Degree|Single|Business: Mgt, Admin|28277|0|2|BFKS|Special Event|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500010765|501395249|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7454|8|||1|
500186742|502397541|500501282|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2031|Green|Amachi|2010-12-02|2010-12-08|2016-06-30|Child: Graduated|Child: Graduated||66.7||4|4|1|1|M|Black||19|Yes|Mother|28227|One Parent: Female|Unknown|||Y|No||School|General Community|Amachi|Match Support|M|Black||52|28227|Masters Degree|Married|Education: Teacher|28227|2|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500013781|500188056|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294, 500004640|-2|0|4|||12183|14|635|1|1|500000294
500186742|500757564|500192033|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1071|Green|Amachi|2007-08-21|2007-08-23|2010-07-29|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||35.2||4|4|3|3|M|Black||19|Yes|Mother|28227|One Parent: Female|Unknown|||Y|No||School|General Community|Amachi|Match Support|M|Black||51|28216||Married|Craftsman||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188056|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294
501185594|501153366|500248756|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3029|Green||2008-02-28|2008-02-29|2016-06-15|Child: Graduated|Child: Graduated||99.5||1|1|1|1|M|Multi-race (Black & White)||19|No|Mother|28227|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Consultant|28226|0|8|Other|Service Organization|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501185866|36|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||7452|6|||1|
500186946|500865596|500181565|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1891|Red|Amachi|2007-06-19|2007-06-20|2012-08-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||62.1||2|2|1|1|F|Black||19|Yes|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||36|28262||Single|Education: Teacher||4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500188139|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500956242|500189847|500259433|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1781|Red||2008-04-14|2008-04-14|2013-02-28|Child/Family: Moved|Child/Family: Moved||58.5||1|1|2|2|M|Multi-Race (None of the above)||19|No|Mother|28210|One Parent: Female|$20,000 to $24,999||||Yes||Therapist/Counselor|General Community||Match Support|M|White||38|28210|||Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500956512|7|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|5|||7464|9|||1|
502312421|502402041|500510430|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|589|Green|Amachi|2011-01-12|2011-01-18|2012-08-29|Volunteer: Moved|Volunteer: Moved||19.4||1|1|1|1|M|Black||19|Yes|Mother|28211|One Parent: Female|Unknown||||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||33|28210|Bachelors Degree|Single|Construction|28269|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502312845|31|0|1|1|0|1|10|2|-2||4|1|500000294|-2||-2|7295|11|||7496|10|||1|500000294
501965241|502081691|500457757|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|763|Green||2010-06-22|2010-06-29|2012-07-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||25.1||1|1|1|1|M|Black||19||Mother|28208|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|M|Black||37|28210||Single|Law||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501578929|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
502934500|503123393|500676924|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|254|Red||2013-01-24|2013-02-19|2013-10-31|Volunteer: Time constraint|Volunteer: Time constraint||8.3||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|M|Black||43|28216|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502935923|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|3|||7464|9|||1|
503108699|503106216|500631547|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|696|Red||2012-08-30|2012-09-14|2014-08-11|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||22.9||1|1|1|1|M|White||19|No|Mother|28031|One Parent: Female|$30,000 to $34,999|||Y|No||Self|General Community||Match Support|M|White||37|28036|Bachelors Degree|Single|Business: Sales|28117|8|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503110361|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502165495|502087652|500460127|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|595|Green||2010-07-07|2010-07-13|2012-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.5||1|1|1|1|F|Black||19|No|Mother|28208|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community||Enrollment|F|White||33|28203|Bachelors Degree|Single|Retail: Sales||2|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502165924|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|5635|9|||7464|9|||1|
501394276|501358317|500311375|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1087|Yellow||2008-11-06|2008-11-19|2011-11-11|Volunteer: Health|Volunteer: Health||35.7||1|1|1|1|F|Black||19|No|Mother|28206|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community||Enrollment|F|White||33|28202|Bachelors Degree|Single|Arts, Entertainment, Sports||2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501394557|31|0|2|1|0|2|5|2|-2||4|2||-2||-2|7016|11|||7464|9|||1|
502462646|502431913|500520035|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|713|Red|2010-2012 OJJDP JJI|2011-02-24|2011-03-18|2013-02-28|Child: Lost interest|Child: Lost interest||23.4||1|1|1|1|F|Black||19|No|Mother|28262|One Parent: Female|$25,000 to $29,999||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||36|28269|PHD|Living w/ Significant Other|Medical: Pharmacist|28217|4|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502463093|31|0|2|31|0|2|10|2|-2||4|3|500005291|-2||-2|0|10|||7464|9|||1|500005291
500186692|501022332|500251970|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|388|Green||2008-03-12|2008-03-17|2009-04-09|Volunteer: Moved|Volunteer: Moved||12.7||7|8|1|1|F|Black||19|No|Mother|28270|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|White||53|28134|Bachelors Degree|Divorced|Construction||5|9|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500188059|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186692|501582415|500381441|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1023|Red||2009-08-28|2009-09-11|2012-06-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||33.6||7|8|1|1|F|Black||19|No|Mother|28270|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|White||50|28270|Some College|Single|Finance: Banking|28217|1|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|500188059|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502307481|502212397|500501813|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|392|Red|Project Big|2010-12-03|2010-12-31|2012-01-27|Volunteer: Time constraint|Volunteer: Time constraint||12.9||1|1|1|1|M|Black||19|No|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|RTBM|M|White||38|28205|Bachelors Degree|Married|Business: Sales||4|0|Other|Service Organization|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500013709|502307910|31|0|1|1|0|1|7|2|500004641||4|3|500004640|-2|500004640|-2|0|4|||7452|6|||1|500004640
500186133|500188930|500036930|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4275|Green||2004-10-14|2004-10-14|2016-06-28|Child: Graduated|Child: Graduated||140.5||1|1|1|1|M|White||18||Mother|28273|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||51|28262|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500187724|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500549982|500917920|500183219|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1161|Green||2007-07-09|2007-08-16|2010-10-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||38.1||1|1|1|1|M|Multi-Race (None of the above)||18||Mother|28027|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||46|28107|Masters Degree|Single|Law: Police Officer|28203|13|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500550234|7|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
501626226|501420794|500350473|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|420|Green||2009-03-18|2009-03-24|2010-05-18|Volunteer: Moved|Volunteer: Moved||13.8||2|2|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||33|28211|||Medical: Admin|28262|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501622822|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501626226|502036832|500457771|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2449|Green||2010-06-22|2010-06-30|2017-03-14|Child: Graduated|Child: Graduated||80.5||2|2|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||33|28203|High School Graduate|Single|Retail: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501622822|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501788773|501845020|500393644|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|975|Green|Amachi|2009-10-12|2009-10-27|2012-06-28|Volunteer: Moved|Volunteer: Moved||32||1|1|1|1|M|Black||18|Yes|Mother|28214|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|RTBM|M|White||33|28202|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501789128|31|0|1|1|0|1|7|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501688212|501814209|500381738|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|320|Red||2009-08-31|2009-09-03|2010-07-20|Child/Family: Moved|Child/Family: Moved||10.5||1|1|1|1|M|Black||18|No|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||34|28202|||Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501688550|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501197292|501240286|500269444|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1394|Green||2008-06-02|2008-06-06|2012-03-31|Volunteer: Moved|Volunteer: Moved||45.8||1|1|1|1|M|White||18|No|Mother|28110|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||50|28112|High School Graduate|Married|Business: Marketing|28105|0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501197566|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500997880|500990660|500237316|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3083|Green||2008-01-14|2008-02-19|2016-07-29|Child: Graduated|Child: Graduated||101.3||1|1|1|1|M|Black||18|No|Mother|28204|Two Parent|$40,000 to $44,999||||Yes||Self|General Community||Match Support|M|White||33|28202|Bachelors Degree|Married|Business: Marketing||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500998153|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502588461|502636478|500546741|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1743|Red|2010-2012 OJJDP JJI|2011-07-19|2011-07-22|2016-04-29|Child: Graduated|Child: Graduated||57.3||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999||||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||46|28278|Bachelors Degree|Separated|Transport: Pilot|28208|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502588977|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2||-2|6854|8|||46|2|||1|500005291
500186910|501091438|500251869|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|438|Green|Amachi|2008-03-12|2008-04-10|2009-06-22|Vol: Other Reason|Vol: Other Reason||14.4||2|2|1|1|F|Black||18|Yes|GrandMother|28208|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Enrollment|F|Black||40|28273|Bachelors Degree|Single|Retail: Mgt||1|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188123|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500186908|501161246|500258298|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|400|Green|Amachi|2008-04-10|2008-04-10|2009-05-15|Volunteer: Moved Vol: Other Reason|Volunteer: Moved|Vol: Other Reason|13.1||2|2|1|1|F|Black||18|Yes|GrandMother|28208|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Enrollment|F|Asian||33|28277|Bachelors Degree|Single|Finance: Economist||0|7|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500188123|31|0|2|4|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
500882189|501535504|500360654|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|678|Green|Amachi|2009-04-30|2009-05-22|2011-03-31|Volunteer: Moved|Volunteer: Moved||22.3||2|2|1|1|F|Black||18|Yes|Mother|28216|One Parent: Female|$20,000 to $24,999||||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Multi-race (Hispanic & White)||34|28211|Bachelors Degree|Single|Business: Human Resources|28280|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501616314|31|0|2|35|0|2|10|2|500003586||4|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
502638767|502570705|500565299|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|246|Red|Project Big, 2010-2012 OJJDP JJI|2011-10-13|2011-10-27|2012-06-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||8.1||1|1|1|1|M|Black||18|No||28206|One Parent: Female|$60,000 to $74,999||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||47|28205||Divorced|Retired||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502639463|31|0|1|1|0|1|10|2|-2||4|3|500005291|-2||-2|0|10|||7464|9|||1|500004640, 500005291
502631914|502581901|500546271|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1127|Red||2011-07-14|2011-07-28|2014-08-28|Volunteer: Moved|Volunteer: Moved||37||1|1|1|1|F|Black||18|No|Mother|28215|One Parent: Female|$20,000 to $24,999||||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|White||37|28205|Associate Degree|Single|Medical: Healthcare Worker|28205|7|10|Local Print|Media|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500013781|502632569|31|0|2|1|0|2|10|2|-2||4|3|500005291|-2|500004640|-2|6854|8|||7439|1|||1|
503469094|501717376|500696470|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1085|Green||2013-05-10|2013-05-10|2016-04-29|Volunteer: Moved|Volunteer: Moved||35.6||1|1|1|1|F|Black||18|No|Mother|28216|Two Parent|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||33|28269|Bachelors Degree|Single|Human Services: Non-Profit|28202|0|8|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|503470960|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|6854|8|||7464|9|||1|
501201377|501497622|500331903|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2764|Red||2009-01-12|2009-01-31|2016-08-26|Child: Graduated|Child: Graduated||90.8||1|1|1|1|F|Hispanic||18|No|Mother|28212|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community||Match Support|F|Hispanic||65|28269|Masters Degree|Single|Medical: Admin|28262|8|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500017777|501201651|3|0|2|3|0|2|10|2|-2||4|3||-2||-2|7016|11|||7446|3|||1|
502070483|502087592|500457368|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|63|Green||2010-06-18|2010-06-22|2010-08-24|Child/Family: Moved|Child/Family: Moved||2.1||1|1|3|3|M|Black||18|Yes|Mother|28269|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|M|Black||45|28262|Bachelors Degree|Married|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500010355|502070907|31|0|1|31|0|1|5|2|500003586||4|1|500000294|-2|500014505, 500015184|-1|34|2|||7462|13|||1|
500185778|500188776|500036776|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4389|Green||2004-06-17|2004-06-17|2016-06-23|Child: Graduated|Child: Graduated||144.2||1|1|1|1|M|Black||18||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||42|27514||Married|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500187368|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500185546|500697858|500150181|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1465|Green|Amachi|2006-12-26|2006-12-26|2010-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||48.1|Y|1|1|1|1|M|Hispanic||18|Yes|Mother|28078|One Parent: Female|Unknown|||Y|No||Faith Organization|General Community|Amachi|Match Support|F|Black||46|28269||Married|Education: Teacher||3|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500187171|3|0|1|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
500417525|500755435|500151964|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2144|Green|Project Big|2007-01-10|2007-01-17|2012-11-30|Volunteer: Time constraint|Volunteer: Time constraint||70.4||1|1|1|1|M|Black||18||Mother|28208|One Parent: Female|Unknown||||No|TV|Media|General Community|Project Big|Match Support|M|White||37|28202|||Medical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500417775|31|0|1|1|0|1|10|2|500004641||4|1|500004640|-2||-2|56|1|||46|2|||1|500004640
502099440|502104508|500460403|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|670|Green||2010-07-09|2010-07-23|2012-05-23|Child/Family: Moved|Child/Family: Moved||22||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|F|Black||26|28262||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|502099867|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|3|||7496|10|||1|
501877073|502035292|500447499|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|124|Yellow||2010-04-15|2010-04-30|2010-09-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||4.1||1|1|2|2|M|Black||18|No|Mother|28215|One Parent: Female|Unknown||||Yes|Radio|Media|General Community||Enrollment|M|Black||40|28215|Some College|Married|Transport: Driver||3|0|Michael Baisden|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|501877446|31|0|1|31|0|1|5|2|-2||4|2||-2||-2|55|1|||11146|1|||1|
501222378|501141328|500261017|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|663|Red||2008-04-15|2008-04-23|2010-02-15|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||21.8||1|1|1|1|M|Black||18|No|Mother|28213|One Parent: Female|$40,000 to $44,999|||Y|Yes|A Child's Place|Service Organization|General Community||Enrollment|M|White||33|28211|Bachelors Degree|Single|Business: Clerical|28211|0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501222654|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|7016|11|||7464|9|||1|
500863413|502632871|500551916|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|524|Red||2011-08-25|2011-09-23|2013-02-28|Volunteer: Moved|Volunteer: Moved||17.2||2|2|2|2|M|White||18|No|Mother|28227|One Parent: Female|$25,000 to $29,999||||No||School|General Community||Match Support|M|White||36|28226|Some College|Single|Business: Marketing||2|4|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|500863682|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|4|||46|2|||1|
500863413|501292217|500281316|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1020|Green||2008-08-11|2008-08-31|2011-06-17|Volunteer: Time constraint|Volunteer: Time constraint||33.5||2|2|1|1|M|White||18|No|Mother|28227|One Parent: Female|$25,000 to $29,999||||No||School|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Finance: Economist||0|6|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500863682|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||7447|3|||1|
502908460|502938939|500616222|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|819|Yellow||2012-05-24|2012-06-07|2014-09-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||26.9||1|1|1|1|F|Hispanic||18|No|Mother|28227|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||40|28079|Bachelors Degree|Single|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502909871|3|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502863781|503002010|500621061|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|913|Red||2012-06-22|2012-07-31|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||30||1|1|1|1|M|Black||18|No|Mother|28031|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|White||26|28031|High School Graduate|Single|Personal Trainer/Coach|28117|0|4|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502865175|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||17161|11|||1|
500865533|500858196|500176255|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|947|Green||2007-05-09|2007-05-14|2009-12-16|Volunteer: Time constraint|Volunteer: Time constraint||31.1||1|1|1|1|M|Black||18|No|Mother|28205|One Parent: Female|$40,000 to $44,999||||No||BBBS Board/Staff|General Community||Match Support|M|Black||32|28212||Single|Student: College||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500865802|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|13|||7462|13|||1|
501226882|500914929|500259581|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1873|Green|Amachi|2008-04-14|2008-04-21|2013-06-07|Volunteer: Time constraint|Volunteer: Time constraint||61.5||1|1|2|2|M|Black||18|Yes|GrandMother|28027|Grandparents|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||52|28027|Bachelors Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|501227158|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||2238|7|||1|500000294
501402710|501728845|500368860|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2189|Green||2009-06-15|2009-06-19|2015-06-17|Child/Family: Moved|Child/Family: Moved||71.9||1|1|1|1|M|Black||18|No|Mother|30058|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||34|28215||Married|Consultant|28285|0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501402995|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501777213|501897253|500417596|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|400|Green||2009-12-02|2009-12-15|2011-01-19|Volunteer: Moved|Volunteer: Moved||13.1||2|2|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||37|28217|Bachelors Degree|Single|Unemployed||0|0|Yahoo!|Web Link|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011639|501777568|31|0|1|31|0|1|5|2|-2||4|1|500005291|-2||-2|0|10|||32|2|||1|
501777213|502475369|500527844|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|414|Green|2010-2012 OJJDP JJI|2011-03-28|2011-04-04|2012-05-22|Volunteer: Moved|Volunteer: Moved||13.6||2|2|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||33|28202|Bachelors Degree|Single|Finance: Banking|28255|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500011746|501777568|31|0|1|31|0|1|5|2|-2||4|1|500005291|-2|500005291|-2|0|10|||7496|10|1202|1|1|500005291
501749652|501645507|500464305|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1163|Yellow||2010-08-05|2010-09-01|2013-11-07|Child/Family: Moved|Child/Family: Moved||38.2||1|1|2|2|M|Black||18||Mother|28213|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|Black||52|28107|Some College|Divorced|Tech: Engineer|28262|3|0|Local Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|501749994|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7437|1|||1|
500730385|500761242|500166676|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1555|Red||2007-03-13|2007-03-15|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||51.1||1|1|1|1|F|Black||18||Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||Match Support|F|Black||38|28217|Bachelors Degree|Single|Finance: Banking|29715|5|0|Recruitment Event|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500730652|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7460|12|||1|
501174643|501687908|500358149|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1282|Red||2009-04-20|2009-05-06|2012-11-08|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||42.1||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|Black||34|28214||Married|Business: Sales|28210|0|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|501174917|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7446|3|||1|
502698998|502692148|500564380|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|853|Yellow||2011-10-12|2011-11-11|2014-03-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||28||1|1|1|1|F|Black||18|No|GrandMother|28211|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28203|Masters Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500012459|502699843|31|0|2|1|0|2|10|2|-2||4|2|500005291|-2||-2|0|4|||7464|9|||1|
501639256|502626656|500612984|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|327|Red||2012-05-02|2012-05-30|2013-04-22|Volunteer: Moved|Volunteer: Moved||10.7||2|2|1|1|M|Multi-Race (None of the above)||18|No|Mother|28211|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||46|28104|Some College|Single|Tech: Support, Writing|28104|3|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501639579|7|0|1|1|0|1|10|2|-2||4|3|500000294|-2||-2|0|10|||7464|9|||1|
501639256|501721160|500360117|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|961|Green|Amachi|2009-04-29|2009-05-04|2011-12-21|Volunteer: Time constraint|Volunteer: Time constraint||31.6||2|2|1|1|M|Multi-Race (None of the above)||18|No|Mother|28211|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Black||35|28212||Single|Human Services: Non-Profit||2|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500003657|501639579|7|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501445222|501159806|500335346|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|515|Green|Amachi|2009-01-23|2009-03-12|2010-08-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||16.9||1|1|1|1|F|Black||18|No|Mother|28202|One Parent: Female|Unknown||||Yes||Relative|General Community|Amachi|Match Support|F|American Indian or Alaska Native||41|28277|Bachelors Degree|Single|Self-Employed, Entrepreneur||6|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501445507|31|0|2|6|0|2|10|2|500003586||4|1|500000294|-2||-2|0|3|||46|2|||1|500000294
501217004|501291789|500350906|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|599|Yellow||2009-03-19|2009-03-23|2010-11-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.7||1|1|1|1|M|Hispanic||18|No|Mother|28104|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||36|28277|Masters Degree|Single|Education: Teacher||0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501217280|3|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502114924|502019135|500457063|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|582|Green||2010-06-16|2010-06-24|2012-01-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.1||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||32|28207|Masters Degree|Single|Medical||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502115351|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|34|2|||7496|10|||1|
501375940|501857916|500410007|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|117|Green||2009-11-12|2009-12-10|2010-04-06|Volunteer: Moved|Volunteer: Moved||3.8||1|1|1|1|M|Black||18|No|Mother|28215|One Parent: Female|Unknown||||No||Service Organization|General Community||Match Support|M|White||33|28211|Bachelors Degree|Single|Business: Marketing|28213|2|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501376219|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|11|||7464|9|||1|
503052841|503122069|500660497|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1512|Green||2012-11-15|2013-01-24|NaT||||49.7||1|1|1|1|F|Hispanic||18|No|Mother|28277|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||24|28104|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503027860|3|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502875778|502885755|500597009|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|413|Red|Amachi|2012-02-08|2012-02-10|2013-03-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||13.6||1|1|1|1|F|Black||18|Yes|Mother|28213|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||44|28216|Associate Degree|Divorced|Finance: Banking||0|5|Charlotte Cares|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502877181|31|0|2|31|0|2|10|2|-2||4|3|500000294|-2||-2|0|10|||11246|6|||1|500000294
501868351|502163779|500463602|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|156|Green||2010-07-29|2010-08-16|2011-01-19|Volunteer: Time constraint|Volunteer: Time constraint||5.1||2|2|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|F|Black||34|28205|Masters Degree|Single|Finance: Accountant||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|501868724|31|0|2|31|0|2|7|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|
501868351|502438990|500515633|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|227|Green|2010-2012 OJJDP JJI|2011-02-04|2011-02-28|2011-10-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.5||2|2|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|F|Black||28|28227|Some College|Single|Student: College|28105|6|0|Big Champions|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|501868724|31|0|2|31|0|2|7|2|-2||4|1|500005291|-2||-2|0|10|||7461|12|||1|500005291
502549784|502558315|500541875|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|708|Green|2010-2012 OJJDP JJI|2011-06-17|2011-06-29|2013-06-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||23.3||1|1|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|$20,000 to $24,999||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||30|28227||Single|Transport: Driver||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502550237|31|0|1|31|0|1|10|2|-2||4|1|500005291|-2|500000294, 500004640|-2|0|10|||7496|10|||1|500005291
503268324|503253968|500676990|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|880|Yellow||2013-01-24|2013-01-26|2015-06-25|Child: Lost interest|Child: Lost interest||28.9||1|1|1|1|M|Black||18|Yes|Mother|28226|One Parent: Female|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Asian||29|28277|Bachelors Degree|Single|Real Estate: Realtor|28277|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503270085|31|0|1|4|0|1|10|2|-2||4|2|500000294|-2||-2|6854|8|||7464|9|||1|
502453042|502632959|500548075|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|726|Red|2010-2012 OJJDP JJI|2011-07-29|2011-08-03|2013-07-29|Volunteer: Time constraint|Volunteer: Time constraint||23.9||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||27|28213|Bachelors Degree|Single|Business: Marketing||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502453489|31|0|2|31|0|2|10|2|-2||4|3|500005291|-2||-2|0|10|||7464|9|||1|500005291
502308593|502262702|500492994|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1647|Red||2010-11-10|2010-11-23|2015-05-28|Child/Family: Moved|Child/Family: Moved||54.1||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||40|28278|Bachelors Degree|Married|Tech: Computer/Programmer||3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502309025|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||12183|14|1209|1|1|
500185812|500188912|500648551|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1305|Green||2012-10-19|2012-10-29|2016-05-26|Child: Graduated|Child: Graduated||42.9||2|3|2|3|F|Black||18|Yes|Mother|28210|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community|Amachi|Match Support|F|White||41|28214|Bachelors Degree|Single|Human Services: Non-Profit||3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|500187400|31|0|2|1|0|2|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|
500732858|500344509|500142645|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1613|Green||2006-11-22|2006-11-28|2011-04-29|Volunteer: Time constraint|Volunteer: Time constraint||53||1|1|1|1|M|Black||18|No|Mother|28203|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28212|Bachelors Degree|Single|Business: Marketing|28202|1|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500733125|31|0|1|1|0|1|5|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|
500948129|500213840|500248197|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|666|Green|Amachi|2008-02-26|2008-03-04|2009-12-30|Volunteer: Time constraint|Volunteer: Time constraint||21.9||2|2|4|4|F|Black||18|No|Mother|28217|One Parent: Female|$25,000 to $29,999|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||44|28078|Bachelors Degree|Single|Business: Mgt, Admin|28210|1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500948399|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
500948129|501891556|500438403|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2296|Green|Amachi|2010-03-01|2010-03-18|2016-06-30|Child: Graduated|Child: Graduated||75.4||2|2|1|1|F|Black||18|No|Mother|28217|One Parent: Female|$25,000 to $29,999|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||40|28203|Some College|Living w/ Significant Other|Finance: Banking|28281|1|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|500948399|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|34|2|||7464|9|||1|500000294
502185074|502490418|500533846|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1909|Green|2010-2012 OJJDP JJI|2011-04-28|2011-05-12|2016-08-02|Child: Graduated|Child: Graduated||62.7||2|2|1|1|F|Black||18|No|GrandMother|28208|Grandparents|Unknown||||Yes|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||68|28262|Bachelors Degree|Living w/ Significant Other|Business: Clerical||2|0|Relative|Relative|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500017732|502185503|31|0|2|31|0|2|10|2|-2||4|1|500005291|-2|500000294, 500004640|-2|5635|9|||17161|11|||1|500005291
502185074|502189418|500462607|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|217|Yellow||2010-07-26|2010-08-16|2011-03-21|Volunteer: Time constraint|Volunteer: Time constraint||7.1||2|2|1|1|F|Black||18|No|GrandMother|28208|Grandparents|Unknown||||Yes|Other|Faith Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28270|Bachelors Degree|Single|Medical: Nurse|28203|3|6|Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|502185503|31|0|2|31|0|2|10|2|-2||4|2|500005291|-2||-2|5635|9|||131|1|||1|
502053779|500189241|500677878|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|562|Red||2013-01-29|2013-02-13|2014-08-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||18.5||2|2|2|2|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||||No|Hampton Crest|Service Organization|General Community||Match Support|F|Black||49|28269|Bachelors Degree|Divorced|Finance|28282|0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|502054203|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|7295|11|||7496|10|||1|
502053779|501912080|500455628|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|813|Red||2010-06-04|2010-06-15|2012-09-05|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||26.7||2|2|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||||No|Hampton Crest|Service Organization|General Community||Match Support|F|Black||39|28216|||Education: College Professor||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502054203|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|7295|11|||7464|9|||1|
501724170|501681407|500370969|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|639|Green||2009-06-24|2009-07-06|2011-04-06|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||21||1|1|1|1|M|Black||18|No|Mother|28210|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|Asian||41|28210|Bachelors Degree|Married|Tech: Management|28255|8|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501724510|31|0|1|4|0|1|5|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
502358538|502078043|500481260|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|343|Green||2010-10-15|2010-11-17|2011-10-26|Child/Family: Moved|Child/Family: Moved||11.3||1|1|1|1|M|White||18|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||68|28107||Married|Retired||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501519460|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
502083495|502089653|500453681|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|512|Red|Amachi|2010-05-20|2010-05-26|2011-10-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.8||1|1|2|2|M|Black||18|Yes|Mother|28025|One Parent: Female|Unknown||||Yes||Service Organization|General Community|Amachi|Match Support|M|Black||52|28027||Married|Business: Human Resources|28273|0|0|Big Champions|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002335|502083919|31|0|1|31|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|11|||7461|12|||1|500000294
502083504|502089653|500454472|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|512|Red|Amachi|2010-05-26|2010-05-26|2011-10-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.8||1|1|2|2|M|Asian||18|Yes|Mother|28025|One Parent: Female|Unknown||||Yes||Service Organization|General Community|Amachi|Match Support|M|Black||52|28027||Married|Business: Human Resources|28273|0|0|Big Champions|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002335|502083919|4|0|1|31|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|11|||7461|12|||1|500000294
500237080|500220237|500057623|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2248|Green|Amachi|2005-11-16|2005-11-16|2012-01-12|Child: Severity of challenges|Child: Severity of challenges||73.9||1|1|2|2|M|Black||18|Yes|Mother|28206|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||40|28269||Married|Business: Marketing||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500237089|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500562813|500696796|500136350|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1209|Green||2006-11-01|2006-11-09|2010-03-02|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||39.7||1|1|1|1|M|Black||18|No|Mother|28217|One Parent: Female|Unknown||||No|AARTF|Neighbor/Friend|General Community||Enrollment|M|Black||38|28273||Single|Tech: Engineer||0|0|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500563065|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|6855|8|||6450|12|||1|
500565502|500805943|500172658|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1093|Green||2007-04-18|2007-04-30|2010-04-27|Volunteer: Moved|Volunteer: Moved||35.9||1|1|1|1|M|Black||18|No|Mother|28269|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||33|28269||Single|Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500565754|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
502230729|502483362|500518850|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|537|Yellow|2010-2012 OJJDP JJI|2011-02-21|2011-03-09|2012-08-27|Volunteer: Moved|Volunteer: Moved||17.6||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||36|28277|Bachelors Degree|Single|Student: College|28205|0|4|Recruitment Event|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|502231160|1|0|1|1|0|1|10|2|-2||4|2|500005291|-2|500000294, 500005291|-2|34|2|||7459|10|||1|500005291
500903162|500952574|500214404|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|988|Green|Amachi|2007-11-05|2007-11-12|2010-07-27|Volunteer: Moved|Volunteer: Moved||32.5||1|1|1|1|F|Black||18|Yes|Mother|28211|One Parent: Female|Less than $10,000|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Black||33|28269|Bachelors Degree|Single|Finance: Banking||1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500903432|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
500383923|500540549|500118470|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2192|Green||2006-08-18|2006-08-30|2012-08-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||72||1|1|2|2|M|Black||18||GrandMother|28205|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||66|28269||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|500384165|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
500186953|500189724|500037838|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2998|Red|Amachi|2004-05-25|2004-05-25|2012-08-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||98.5||1|1|2|2|M|Black||18|Yes|GrandMother|28214|Other Relative|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||45|28207||Single|Unknown|28209|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500188126|31|0|1|1|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
503216769|503344849|500698465|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1348|Red||2013-05-29|2013-06-21|2017-02-28|Child/Family: Moved|Child/Family: Moved||44.3||1|1|2|2|F|Black||18|No|Mother|28262|Two Parent|$75,000 to $99,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|Black||25|28269|Bachelors Degree|Single|Education: Teacher|28210|0|4|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503218550|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|34|2|||46|2|||1|
502570396|502545897|500539251|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1561|Green|2010-2012 OJJDP JJI|2011-06-01|2011-06-30|2015-10-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||51.3||1|1|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28215|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||35|28078|Bachelors Degree|Single|Tech: Computer/Programmer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|502570850|38|0|2|31|0|2|10|2|-2||4|1|500005291|-2||-2|34|2|||46|2|||1|500005291
501188642|501507244|500359356|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|822|Red||2009-04-24|2009-04-28|2011-07-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27||1|1|1|1|M|Black||18|No|Mother|28105|One Parent: Female|$45,000 to $49,999||||No||Neighbor/Friend|General Community||Match Support|M|White||56|28270|Bachelors Degree|Married|Real Estate: Realtor|28277|11|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501188916|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|8|||7496|10|||1|
500901271|501083173|500256530|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|796|Red||2008-04-03|2008-04-07|2010-06-12|Volunteer: Time constraint|Volunteer: Time constraint||26.2||2|2|1|1|M|Black||18|Yes|Mother|28216|One Parent: Female|$30,000 to $34,999||||No||Self|General Community|Amachi|RTBM|M|White||40|28269|Associate Degree|Single|Tech: Engineer||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500901541|31|0|1|1|0|1|7|2|||4|3|500000294|-2||-2|0|10|||46|2|||1|
500901271|502310515|500509461|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|230|Red|Amachi|2011-01-06|2011-01-12|2011-08-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.6||2|2|1|1|M|Black||18|Yes|Mother|28216|One Parent: Female|$30,000 to $34,999||||No||Self|General Community|Amachi|RTBM|M|Some Other Race||39|28216||Single|Retail: Sales||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|500901541|31|0|1|41|0|1|7|2|-2||4|3|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
502501319|502507619|500530032|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|179|Green|2010-2012 OJJDP JJI|2011-04-08|2011-04-29|2011-10-25|Volunteer: Time constraint|Volunteer: Time constraint||5.9||2|2|1|1|F|Black||18|No|Mother|28269|One Parent: Female|$45,000 to $49,999||||No||Relative|General Community|2010-2012 OJJDP JJI|Match Support|F|White||57|28269|Associate Degree|Single|Business: Sales|10580|14|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011184|502501768|31|0|2|1|0|2|10|2|-2||4|1|500005291|-2||-2|0|3|||7464|9|||1|500005291
502501319|502893544|500597799|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|182|Red||2012-02-13|2012-02-29|2012-08-29|Child: Lost interest|Child: Lost interest||6||2|2|1|1|F|Black||18|No|Mother|28269|One Parent: Female|$45,000 to $49,999||||No||Relative|General Community|2010-2012 OJJDP JJI|Match Support|F|White||50|28031|Some College|Married|Retired||0|0|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502501768|31|0|2|1|0|2|10|2|-2||4|3|500005291|-2||-2|0|3|||7438|1|||1|
502045258|502190790|500457916|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2257|Green||2010-06-23|2010-06-25|2016-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||74.2||1|1|1|1|F|Black||18|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||33|28262|Bachelors Degree|Single|Medical: Nurse|28262|4|9|AA Task Force|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502045664|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||6247|12|||1|
500186174|500189225|500038037|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|2652|Red||2005-09-06|2005-07-28|2012-10-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||87.1||2|2|2|2|F|Black||18||Mother|28208|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|F|Black||48|29715|Some College|Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011746|500187758|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502114704|502130736|500460157|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|508|Green||2010-07-07|2010-08-20|2012-01-10|Volunteer: Moved|Volunteer: Moved||16.7||1|1|1|1|F|Black||18|No|Mother|28270|One Parent: Female|Unknown||||Yes|Radio|Media|General Community||RTBM|F|White||32|28204|Masters Degree|Single|Business: Marketing||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502115131|31|0|2|1|0|2|7|2|-2||4|1||-2||-2|55|1|||7496|10|||1|
501614902|501745988|500370268|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|637|Green|Amachi|2009-06-22|2009-07-02|2011-03-31|Child/Family: Moved|Child/Family: Moved||20.9||1|1|1|1|M|Black||18|Yes|Mother|28105|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Black||39|28205|Bachelors Degree|Single|Business: Engineer||2|5|AA Task Force|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501615222|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||9226|6|||1|500000294
502510347|502677833|500557844|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1765|Green|2010-2012 OJJDP JJI|2011-09-26|2011-10-31|2016-08-30|Child: Graduated|Child: Graduated||58||1|1|1|1|F|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28262|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502510796|31|0|2|31|0|2|10|2|-2||4|1|500005291|-2||-2|0|5|||7464|9|||1|500005291
501285489|501185576|500274170|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|512|Green||2008-06-19|2008-06-19|2009-11-13|Child/Family: Moved|Child/Family: Moved||16.8||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|M|White||32|28203|Bachelors Degree|Married|Business: Marketing||0|2|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501285767|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|8|||46|2|||1|
500796255|501846438|500424314|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2612|Green||2010-01-04|2010-01-20|NaT||||85.8||3|3|1|1|M|White||18|No|Mother|28031|One Parent: Male|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||60|28269|||Medical: Admin|28207|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|500796529|1|0|1|1|0|1|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1|
500796255|501414689|500317055|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|303|Green||2008-11-18|2008-11-25|2009-09-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10||3|3|1|1|M|White||18|No|Mother|28031|One Parent: Male|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28269|Bachelors Degree|Married|Service: Restaurant||0|6|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500796529|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
500740295|500794907|500179696|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2586|Yellow||2007-06-11|2007-06-12|2014-07-11|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||85||1|1|1|1|M|Black||18||Mother|28216|One Parent: Female|$20,000 to $24,999||||No||Therapist/Counselor|General Community||Match Support|M|White||55|28216|Bachelors Degree|Divorced|Tech: Engineer||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500740560|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|5|||46|2|||1|
500185534|500189461|500093294|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2413|Red||2006-05-11|2006-05-13|2012-12-20|Child: Family structure changed|Child: Family structure changed||79.3||1|1|3|5|M|Black||18||Mother|28204|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||63|28206|Some College|Married|Self-Employed, Entrepreneur|28206|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500004169|500187159|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501176569|501457533|500327489|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1147|Green||2008-12-17|2009-01-08|2012-02-29|Child/Family: Moved|Child/Family: Moved||37.7||1|1|1|1|M|Multi-race (Black & White)||18||Mother|28031|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||32|28078|Bachelors Degree|Living w/ Significant Other|Education: Admin|28035|2|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501176843|36|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
501716075|501216868|500356008|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|309|Green||2009-04-07|2009-04-07|2010-02-10|Child: Lost interest|Child: Lost interest||10.2||1|1|3|3|M|Black||18|No|Mother|28025|Two Parent|Unknown||||No||School|General Community||Match Support|M|White||32|28078||Single|Education: Teacher||0|0|other|College Partner|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500002335|501716414|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|4|||7670|5|||1|
501938887|502014005|500447313|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|544|Red||2010-04-14|2010-04-30|2011-10-26|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.9||1|1|1|1|M|Black||18|No|Mother|28205|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|M|White||34|28205|||Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501939285|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|8|||7496|10|||1|
500252077|501365749|500317108|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2613|Red|Amachi|2008-11-18|2008-11-24|2016-01-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||85.8||3|3|1|1|M|Black||18|Yes|Mother|28215|One Parent: Female|Unknown||||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||32|28202|Bachelors Degree|Single|Tech: Computer/Programmer||0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501750989|31|0|1|1|0|1|10|2|500003586||4|3|500000294|-2||-2|7295|11|||46|2|||1|500000294
502370669|503472866|500700192|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1363|Green||2013-06-11|2013-06-22|NaT||||44.8||2|2|1|1|M|Black||18|No|Mother|28269|One Parent: Female|$40,000 to $44,999|||Y|Yes||Self|General Community||Match Support|M|White||57|28277|Some College|Married|Business: Sales||28|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502371107|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502370669|502731507|500573204|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|358|Red||2011-11-01|2011-12-07|2012-11-29|Volunteer: Moved|Volunteer: Moved||11.8||2|2|1|1|M|Black||18|No|Mother|28269|One Parent: Female|$40,000 to $44,999|||Y|Yes||Self|General Community||Match Support|M|Some Other Race||31|28205|Masters Degree|Single|Finance|28777|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502371107|31|0|1|41|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
501535016|501438980|500331054|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|982|Yellow||2009-01-07|2009-01-12|2011-09-21|Volunteer: Time constraint|Volunteer: Time constraint||32.3||1|1|1|1|F|Black||18|No|Mother|28273|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||36|28277|Masters Degree|Single|Finance: Banking||0|1|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|501535308|31|0|2|31|0|2|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1|
502034622|502127058|500456536|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|29|Green||2010-06-11|2010-06-23|2010-07-22|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||1||1|1|2|2|M|Black||18|No|Mother|28214|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|502035021|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||130|1|||1|
501781058|501429731|500367177|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|191|Green||2009-06-02|2009-06-02|2009-12-10|Volunteer: Time constraint|Volunteer: Time constraint||6.3||1|1|1|1|F|White||18|No|Mother|28075|Two Parent|Unknown||||No||Relative|General Community||Match Support|F|White||50|28078|High School Graduate|Married|Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501781413|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
502290482|501861156|500503975|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|311|Green||2010-12-09|2010-12-18|2011-10-25|Volunteer: Moved|Volunteer: Moved||10.2||2|2|1|1|F|Black||18|No|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||34|28202|Masters Degree||Finance: Banking||0|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011184|502290914|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294, 500004640|-2|0|10|||7464|9|||1|
502290482|503002021|500677084|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|387|Yellow||2013-01-24|2013-01-26|2014-02-17|Child/Family: Moved|Child/Family: Moved||12.7||2|2|1|1|F|Black||18|No|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||28|28209|Bachelors Degree|Single|Education: Teacher|29708|2|0|Local Print|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502290914|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7439|1|||1|
500402982|500467614|500103313|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1790|Green|Amachi|2006-06-29|2006-06-29|2011-05-24|Volunteer: Moved|Volunteer: Moved||58.8||1|1|1|1|M|White||18||Mother|28211|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||37|28212||Single|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500402926|1|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
500186215|501322823|500284070|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|245|Green|Amachi|2008-08-27|2008-10-20|2009-06-22|Vol: Lost Interest|Vol: Lost Interest||8||4|5|1|1|M|Multi-Race (None of the above)||18|Yes|GrandMother|28214|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||34|28214|Some College|Married|Business: Mgt, Admin|28217|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500187776|7|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||7462|13|||1|500000294
501729405|502361956|500501689|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|915|Green|Amachi, Project Big, Project Big AND Amachi|2010-12-02|2010-12-14|2013-06-16|Volunteer: Moved|Volunteer: Moved||30.1||2|2|1|1|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|RTBM|F|White||33|28204|Bachelors Degree|Single|Business: Sales|28210|0|7|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|501729745|31|0|2|1|0|2|7|2|500004772||4|1|500000294, 500004640, 500004901|-2|500000294|-2|0|4|||7464|9|||1|500000294, 500004640, 500004901
501729405|501443657|500379612|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|433|Yellow|Amachi, Project Big, Project Big AND Amachi|2009-08-18|2009-08-18|2010-10-25|Volunteer: Time constraint|Volunteer: Time constraint||14.2||2|2|1|1|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|RTBM|F|Black||30|28262|Bachelors Degree|Single|Finance: Banking|28288|0|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|501729745|31|0|2|31|0|2|7|2|500004772||4|2|500000294, 500004640, 500004901|-2||-2|0|4|||7464|9|||1|500000294, 500004640, 500004901
502698363|502641410|500557390|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|780|Red|Amachi|2011-09-23|2011-10-18|2013-12-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25.6||1|1|1|1|M|Black||18|Yes|GrandMother|28203|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Enrollment|M|Black||43|28208|Bachelors Degree|Single|Education|28217|0|0|Other|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502699208|31|0|1|31|0|1|5|2|500003586||4|3|500000294|-2||-2|0|10|||7452|6|||1|500000294
500853690|500846213|500173015|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1537|Yellow||2007-04-20|2007-05-07|2011-07-22|Child/Family: Moved|Child/Family: Moved||50.5||1|1|1|1|F|Multi-Race (None of the above)||18|No|Mother|28214|One Parent: Female|$15,000 to $19,999|||Y|No||BBBS Board/Staff|General Community||Match Support|F|White||38|28226||Living w/ Significant Other|Child/Day Care Worker||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500853959|7|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|13|||46|2|||1|
502868925|502885744|500607510|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Red||2012-04-02|2012-04-25|2014-09-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||35|28262|Bachelors Degree|Divorced|Finance: Banking||2|6|Charlotte Cares|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502870324|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||11246|6|||1|
501237971|501598429|500649363|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1202|Green||2012-10-23|2012-11-17|2016-03-03|Volunteer: Moved|Volunteer: Moved||39.5||2|2|3|3|F|Black||18|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||41|28269|||Business: Human Resources|28206|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503287812|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|
501237971|500839927|500257150|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|475|Green|Amachi|2008-04-07|2008-04-18|2009-08-06|Child/Family: Moved|Child/Family: Moved||15.6||2|2|2|2|F|Black||18|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||32|28075|Bachelors Degree||Child/Day Care Worker|28075|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|503287812|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||46|2|||1|500000294
501160894|501442606|500309909|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1020|Yellow||2008-11-04|2008-11-07|2011-08-24|Child/Family: Moved|Child/Family: Moved||33.5||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|$10,000 to $14,999||||Yes||Self|General Community||Match Support|M|White||33|28204||Single|Real Estate: Realtor|28204|2|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501161168|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503425736|503519747|500711543|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|973|Green||2013-09-17|2013-10-16|2016-06-15|Child: Graduated|Child: Graduated||32||1|1|1|1|F|Black||18|No|GrandMother|28213|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|White||29|28211|Juris Doctorate (JD)|Married|Law|28202|0|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503427601|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502317496|502860968|500602986|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|432|Red||2012-03-08|2012-04-12|2013-06-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.2||1|1|1|1|M|Black||18|Yes|Mother|28214|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, Project Big|Match Support|M|Black||42|28214|Some College|Married|Business|28217|17|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502317931|31|0|1|31|0|1|10|2|500004641||4|3|500000294, 500004640|-2||-2|0|4|||7462|13|||1|
502581751|502587677|500542041|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1046|Yellow||2011-06-20|2011-06-27|2014-05-08|Volunteer: Moved|Volunteer: Moved||34.4||1|1|1|1|M|Black||18|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||38|28206|Masters Degree|Single|Business: Human Resources|28255|4|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502582259|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501037140|501171628|500261234|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|512|Green||2008-04-16|2008-04-29|2009-09-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.8||1|1|1|1|M|Some Other Race||18|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|Hispanic||48|28277|High School Graduate|Domestic Partner|Business: Mgt, Admin|28217|1|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|501037413|41|0|1|3|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500791567|500578720|500155823|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2262|Yellow||2007-01-31|2007-01-31|2013-04-11|Volunteer: Time constraint|Volunteer: Time constraint||74.3||1|1|2|2|M|Multi-Race (None of the above)||18|No|Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||Match Support|M|Black||32|28215||Married|Finance: Banking||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500187654|7|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7447|3|||1|
501206897|501077272|500263885|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1141|Green||2008-04-30|2008-05-02|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||37.5||1|1|1|1|M|White||18|No|Mother|28215|One Parent: Female|$10,000 to $14,999||||Yes||Therapist/Counselor|General Community||Match Support|M|White||39|28204|Bachelors Degree|Married|Self-Employed, Entrepreneur|28208|8|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501207171|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|5|||7496|10|||1|
502421176|502419727|500517478|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|742|Red|2010-2012 OJJDP JJI|2011-02-14|2011-03-10|2013-03-21|Volunteer: Time constraint|Volunteer: Time constraint||24.4||2|2|1|1|F|Black||18|No|GrandMother|28214|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||33|28273|Bachelors Degree|Single|Insurance||0|0|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500004169|502421614|31|0|2|31|0|2|10|2|-2||4|3||-2|500000294, 500004640|-2|0|4|||46|2|||1|500005291
502421176|503497451|500710577|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1256|Green||2013-09-12|2013-09-30|2017-03-09|Volunteer: Time constraint|Volunteer: Time constraint||41.3||2|2|1|1|F|Black||18|No|GrandMother|28214|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||26|28078|Masters Degree|Single|Education: Teacher|28212|0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502421614|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502206676|502562455|500535587|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|147|Green|Amachi|2011-05-10|2011-05-31|2011-10-25|Child: Severity of challenges|Child: Severity of challenges||4.8||1|1|1|1|M|Black||18|Yes|Mother|28216|Other Relative|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|M|White||47|28269|Bachelors Degree|Married|Education: Teacher||7|0|Local Print|Media|Big|General Community|Amachi|RTBM|0|1|1|0|277|60|598|500000170|500011184|502207102|31|0|1|1|0|1|10|2|500003586||4|1|500000294, 500004640, 500004901|-2|500000294|-2|7016|11|||7439|1|||1|500000294
501340102|501316292|500287888|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1665|Red|Amachi|2008-09-12|2008-10-03|2013-04-25|Child/Family: Time constraints|Child/Family: Time constraints||54.7||1|1|1|1|M|Multi-race (Black & Hispanic)||18|Yes|Mother|28262|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||50|28269|Masters Degree|Married|Customer Service|28269|8|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501340381|38|0|1|1|0|1|10|2|500003586||4|3|500000294|-2||-2|0|10|||7464|9|||1|500000294
500341548|501503307|500348207|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|321|Green||2009-03-10|2009-03-11|2010-01-26|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||10.5||4|4|1|1|F|White||18|No|Father|28025|One Parent: Male|Unknown||||No||Relative|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||59|28027|Bachelors Degree|Divorced|Law: Police Officer|28075|7|1|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500002335|500341682|1|0|2|1|0|2|10|2|-2||4|1|500014681, 500016374|-2||-2|0|3|||7464|9|||1|
501250109|501790515|500381167|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1265|Red||2009-08-27|2009-09-11|2013-02-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||41.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28227|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501250385|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|6854|8|||7464|9|||1|
501730483|501721615|500368696|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|150|Green||2009-06-12|2009-07-17|2009-12-14|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||4.9||1|1|2|2|M|Black||18|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Hispanic||47|28215||Married|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501730818|31|0|1|3|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501730480|501588964|500365950|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|209|Green||2009-05-27|2009-05-28|2009-12-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||6.9||1|1|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||34|28210||Married|Business: Mgt, Admin|28255|0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501730818|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
501388847|501452657|500334726|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|971|Green||2009-01-21|2009-01-25|2011-09-23|Volunteer: Moved|Volunteer: Moved||31.9||1|1|1|1|M|Black||18|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||31|28202|Bachelors Degree|Single|Medical: Healthcare Worker|28207|1|5|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501389128|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7446|3|||1|
502805818|502704456|500585665|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|736|Green|Amachi|2011-12-09|2011-12-14|2013-12-19|Child/Family: Moved|Child/Family: Moved||24.2||1|1|1|1|F|Black||18|Yes|GrandMother|28205|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||45|28213|Some College|Single|Business: Mgt, Admin|28202|1|3|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500015820|502807093|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501621811|501621016|500344465|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2915|Yellow|Project Big|2009-02-24|2009-03-16|2017-03-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||95.8||1|1|1|1|F|Black||18|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||36|28269||Married|Self-Employed, Entrepreneur|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501622131|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|500004640
502227959|502198861|500462034|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|75|Red||2010-07-21|2010-07-23|2010-10-06|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||2.5||1|1|1|1|M|Black||18|No|GrandMother|28036|Grandparents|Unknown||||Yes||Relative|General Community||Match Support|M|White||56|28031|High School Graduate|Married|Consultant|28031|25|0|BFKS|Special Event|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|502228390|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|3|||7454|8|||1|
503026933|503758613|500761412|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|518|Yellow||2014-04-28|2014-05-30|2015-10-30|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17||2|2|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28216|Two Parent|$35,000 to $39,999|||Y|Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||37|28031|Masters Degree|Single|Business: Mgt, Admin|94103|1|1|BBBS National Site|Web Link|Big|General Community|VOL - Mentoring Hispanic Youth|Enrollment|0|1|0|1|277|60|598|500000170|500008321|503028507|38|0|2|1|0|2|10|2|-2||4|2|500011312|-2|500011312|-2|0|10|||46|2|||1|
503026933|503111607|500660471|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|216|Red||2012-11-15|2012-12-27|2013-07-31|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||7.1||2|2|1|1|F|Multi-race (Black & Hispanic)||18|No|Mother|28216|Two Parent|$35,000 to $39,999|||Y|Yes||Self|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|Black||33|28216|Bachelors Degree|Single|Finance: Banking|28269|6|10|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503028507|38|0|2|31|0|2|10|2|-2||4|3|500011312|-2||-2|0|10|||7496|10|||1|
500186645|500189545|500037636|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|4234|Green|Amachi|2004-06-03|2004-06-03|2016-01-06|Child: Graduated|Child: Graduated||139.1||1|1|1|1|M|Black||18|Yes|Mother|28208|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||51|28256|High School Graduate|Married|Unemployed||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|0|1|277|60|598|500000170|500018987|500188043|31|0|1|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502221904|502056302|500464397|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|909|Red|Amachi|2010-08-05|2010-08-06|2013-01-31|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||29.9||1|1|3|3|F|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||||Yes|Arby's|Workplace Partner/Business|General Community||Match Support|F|Black||36|28078|Masters Degree|Married|Business: Marketing|28273|1|1|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|0|1|1|0|277|60|598|500000170|500015820|502222335|31|0|2|31|0|2|10|2|500003586||4|3||-2|500014505, 500014506|-1|3394|14|||7671|13|||1|500000294
502183055|501035952|500463671|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|701|Red||2010-07-30|2010-07-30|2012-06-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||23||1|1|2|2|F|Black||18|No|Mother|28226|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||35|28270|Bachelors Degree|Single|Human Services: Social Worker||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502183484|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
500887862|500923430|500530980|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2164|Green|Cabarrus County|2011-04-13|2011-04-13|NaT||||71.1||2|2|2|2|F|Black||18|Yes|Mother|28025|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|F|Black||43|28027||Divorced|Finance: Banking||0|7|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|500888132|31|0|2|31|0|2|10|2|500016307||2|1|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|500016374
502839827|503311280|500677083|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1505|Green||2013-01-24|2013-01-31|NaT||||49.4||1|1|1|1|M|Black||18|No|Mother|28215|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|Black||41|28105|Bachelors Degree|Single|Tech: Management|28202|0|6|AA Task Force|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502841119|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||6247|12|||1|
501588819|501454413|500373948|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|680|Green||2009-07-14|2009-07-29|2011-06-09|Volunteer: Time constraint|Volunteer: Time constraint||22.3||2|2|1|1|F|Black||18||Mother|28208|Two Parent|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28273|Masters Degree|Single|Govt: Mgmt/Admin|28216|1|0|Newspaper|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501589139|31|0|2|31|0|2|10|2|-2||4|1|500004640, 500005291|-2||-2|0|10|||129|1|||1|
501588819|502643880|500552861|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|266|Green|Project Big, 2010-2012 OJJDP JJI|2011-08-31|2011-08-31|2012-05-23|Volunteer: Time constraint|Volunteer: Time constraint||8.7||2|2|1|1|F|Black||18||Mother|28208|Two Parent|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Hispanic||32|28273|Bachelors Degree|Single|Medical: Admin|28277|0|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501589139|31|0|2|3|0|2|10|2|-2||4|1|500004640, 500005291|-2||-2|0|10|||7464|9|||1|500004640, 500005291
500187011|501391987|500320719|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|596|Green|Amachi|2008-11-26|2008-12-08|2010-07-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.6||3|3|1|1|M|Multi-Race (None of the above)||18|No|Mother|28227|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Amachi|RTBM|M|White||34|28262|Bachelors Degree|Single|Finance: Banking||3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500188147|7|0|1|1|0|1|7|2|500003586||4|1|500000294|-2||-2|6854|8|||7464|9|||1|500000294
500859789|500856753|500169338|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2163|Red|Amachi|2007-03-29|2007-03-29|2013-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||71.1||1|1|1|1|F|Black||18|Yes|Mother|28208|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||65|28078|||Business: Mgt, Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008321|500860058|31|0|2|31|0|2|10|2|-2||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502482929|502489447|500531863|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|211|Red|2010-2012 OJJDP JJI|2011-04-19|2011-05-16|2011-12-13|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.9||1|1|1|1|M|Black||18|No|Mother|28078|One Parent: Female|Less than $10,000|||Y|Yes|Billboard|Media|General Community|2010-2012 OJJDP JJI|RTBM|M|Black||31|28227||Single|Retail: Mgt|28104|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502483376|31|0|1|31|0|1|7|2|-2||4|3|500005291|-2||-2|50|1|||7496|10|||1|500005291
501604443|501729878|500371104|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2806|Green||2009-06-25|2009-07-10|NaT||||92.2||1|1|1|1|M|Black||18|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||35|28209|Bachelors Degree|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501604760|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
500849042|501379402|500314655|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|767|Green||2008-11-13|2008-11-14|2010-12-21|Child/Family: Moved|Child/Family: Moved||25.2||2|3|1|1|F|Black||18|No|Mother|28206|One Parent: Female|Unknown||||No||Service Organization|General Community||Match Support|F|Black||33|28202|Bachelors Degree|Divorced|Finance: Accountant||0|4|Recruitment Event|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500849311|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|11|||7446|3|||1|
500767213|501175210|500263514|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|965|Green||2008-04-28|2008-04-30|2010-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.7||1|1|1|1|F|Black||18||Mother|28216|One Parent: Female|Unknown|||Y|No||Self|General Community|Project Big|Enrollment|F|White||44|28207||Married|Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500767473|31|0|2|1|0|2|5|2|-2||4|1|500004640|-2||-2|0|10|||7464|9|||1|
500826594|500920342|500185735|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3221|Green||2007-07-23|2007-08-21|2016-06-15|Child: Graduated|Child: Graduated||105.8||1|1|1|1|M|Black||18|No|Mother|28226|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|M|Some Other Race||36|28209|||Business: Sales||0|0|General|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500826861|31|0|1|41|0|1|10|2|-2||4|1||-2||-2|0|5|||6450|12|||1|
501378357|501174997|500339619|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2953|Green||2009-02-09|2009-02-13|NaT||||97||1|1|2|2|M|Multi-race (Black & White)||18|No|Mother|28213|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Mgt, Admin|28215|10|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501378636|36|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502162474|502536516|500533468|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|666|Red|2010-2012 OJJDP JJI|2011-04-26|2011-05-04|2013-02-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||21.9||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||35|28205|Associate Degree|Single|Student: College|28213|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502162903|31|0|1|1|0|1|5|2|-2||4|3|500005291|-2||-2|0|10|||7496|10|||1|500005291
502578459|502869485|500615803|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1697|Yellow|Cabarrus County|2012-05-22|2012-07-23|NaT||||55.8||1|1|1|1|M|Black||18|No|Mother|28025|One Parent: Female|$35,000 to $39,999|Yes: Active|No||Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||48|28269|Some College|Married|Tech: Management|28204|10|0|AA Task Force|BBBS Board/Staff|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502578962|31|0|1|31|0|1|10|2|500016307||2|2|500016374|-2|500016374|-2|6854|8|||9229|13|||1|500016374
501015962|501065096|500241396|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1570|Yellow|Amachi|2008-01-31|2008-02-12|2012-05-31|Volunteer: Time constraint|Volunteer: Time constraint||51.6||1|1|1|1|F|Black||18|Yes|GrandMother|28208|One Parent: Female|Less than $10,000||||Yes||Self|General Community|Amachi|Enrollment|F|White||33|28202|Bachelors Degree|Single|Education: Teacher|28025|1|4|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|501016235|31|0|2|1|0|2|5|2|500003586||4|2|500000294|-2||-2|0|10|||2238|7|||1|500000294
500186760|500189588|500037690|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2269|Green|Amachi|2004-08-09|2004-08-09|2010-10-26|Child: Family structure changed|Child: Family structure changed||74.5||1|1|1|1|M|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||||No|TV|Media|General Community|Amachi|Match Support|M|Black||43|28269|Bachelors Degree|Married|Finance: Banking||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188154|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|56|1|||2238|7|||1|500000294
501631059|501589359|500364875|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1203|Yellow||2009-05-21|2009-05-26|2012-09-10|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||39.5||1|1|1|1|F|Black||18|No|Mother|28202|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||29|28216|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501631382|31|0|2|31|0|2|10|2|-2||4|2||-2|500000294|-2|34|2|||7464|9|||1|
502980471|503258884|500678978|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|150|Red||2013-01-31|2013-02-16|2013-07-16|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||4.9||1|1|2|2|M|Black||18|No|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community|Project Big|Match Support|M|Asian|Indian|27|28277|Bachelors Degree|Single|Business|28277|0|2||Relative|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|502981923|31|0|1|4|18|1|10|2|-2||4|3|500004640|-2||-2|34|2|||0|11|||1|
500187059|500188568|500038123|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1377|Green|Amachi|2005-09-08|2005-09-08|2009-06-16|Child/Family: Lost contact with volunteer/agency Child: Lost interest|Child/Family: Lost contact with volunteer/agency|Child: Lost interest|45.2||1|1|1|1|M|Black||18|Yes|Mother|28212|One Parent: Female|Unknown|||Y|No||Neighbor/Friend|General Community|Amachi|Match Support|M|Black||45|28215|Bachelors Degree|Single|Human Services: Youth Worker||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500003657|500188021|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|8|||2238|7|||1|500000294
503039131|503483337|500703051|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|118|Red||2013-07-09|2013-07-26|2013-11-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.9||1|1|2|2|F|Black||18|No|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||45|28227|Bachelors Degree|Married|Customer Service|28262|18|0|Big For A Day|Special Event|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|503040727|31|0|2|31|0|2|5|2|-2||4|3||-2|500000294|-2|0|10|||16422|8|||1|
502177920|502387867|500509427|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|495|Red||2011-01-06|2011-01-14|2012-05-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.3||1|1|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||59|28212|Associate Degree|Divorced|Transport: Driver|28269|0|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500011746|502178349|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2||-2|34|2|||12183|14|||1|
502604900|502582742|500577855|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1276|Green||2011-11-14|2011-11-15|2015-05-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||41.9||1|1|1|1|M|White||18|No|Mother|28105|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||30|28211|Bachelors Degree|Single|Finance: Accountant|28204|0|5|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017777|502605417|1|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|6854|8|||7464|9|||1|
502974629|503188801|500682863|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1309|Red||2013-02-19|2013-02-25|2016-09-26|Child/Family: Moved|Child/Family: Moved||43||1|1|1|1|M|Black||18|No|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||33|28209|Bachelors Degree|Married|Business: Mgt, Admin|28202|6|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502976067|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500392860|501064465|500236600|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1288|Green||2008-01-10|2008-01-18|2011-07-29|Volunteer: Moved|Volunteer: Moved||42.3||2|2|2|2|M|Black||18||Aunt|28215|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community||Match Support|M|White||43|28227|High School Graduate|Married|Clergy||10|0|General|Other Big|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500008629|500393108|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|5|||6450|12|||1|
502472483|502453698|500518061|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1277|Red|Amachi|2011-02-16|2011-02-28|2014-08-28|Volunteer: Time constraint|Volunteer: Time constraint||42||1|1|1|1|F|Black||18|Yes|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||33|28202|Bachelors Degree|Single|Education|28208|4|10|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500013781|502472930|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2|500004640|-2|0|10|||7464|9|||1|500000294
500969481|501202092|500274109|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1178|Yellow|Project Big|2008-06-19|2008-07-22|2011-10-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38.7||1|1|2|2|F|Black||18|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|No||Therapist/Counselor|General Community||Match Support|F|Black||41|28209|Bachelors Degree|Single|Finance: Banking|28255|0|6|TV|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011639|500969749|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|5|||130|1|||1|500004640
501234599|501236882|500272343|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|552|Green||2008-06-12|2008-06-24|2009-12-28|Volunteer: Time constraint|Volunteer: Time constraint||18.1||3|3|1|1|M|Black||18|No|Mother|28215|Grandparents|Unknown||||No|TV|Media|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||47|28262|Some College|Divorced|Unknown|28204|10|0|Recruitment Event|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501234875|31|0|1|31|0|1|5|2|-2||4|1|500005291|-2||-2|56|1|||7458|9|||1|
501234599|501948189|500430307|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|64|Green||2010-01-27|2010-03-09|2010-05-12|Volunteer: Time constraint|Volunteer: Time constraint||2.1||3|3|1|1|M|Black||18|No|Mother|28215|Grandparents|Unknown||||No|TV|Media|General Community|2010-2012 OJJDP JJI|Enrollment|M|Multi-race (Hispanic & White)||40|28210|||Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501234875|31|0|1|35|0|1|5|2|-2||4|1|500005291|-2||-2|56|1|||7464|9|||1|
501234599|501974562|500462663|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|386|Green||2010-07-26|2010-08-09|2011-08-30|Volunteer: Time constraint|Volunteer: Time constraint||12.7||3|3|1|1|M|Black||18|No|Mother|28215|Grandparents|Unknown||||No|TV|Media|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||29|28215|||Retail: Sales||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501234875|31|0|1|1|0|1|5|2|-2||4|1|500005291|-2||-2|56|1|||7464|9|||1|
501072636|501637727|500368653|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1455|Red||2009-06-12|2009-06-25|2013-06-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||47.8||2|2|1|1|M|White||18||Mother|28134|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||50|28277|Bachelors Degree|Married|Tech: Management||10|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500004169|500965396|1|0|1|1|0|1|10|2|-2||4|3||-2|500000294|-2|0|10|||7462|13|||1|
501072636|500960208|500252733|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|326|Green||2008-03-17|2008-04-07|2009-02-27|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||10.7||2|2|1|1|M|White||18||Mother|28134|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||47|28277||Married|Service: Restaurant||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500965396|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501212047|501242250|500264889|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3235|Green||2008-05-06|2008-05-07|NaT||||106.3||1|1|1|1|F|White||18|No|Father|28207|One Parent: Male|Unknown||||No||Self|General Community||Match Support|F|White||33|28226||Single|Human Services: Non-Profit|28205|0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501212321|1|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503110827|503278385|500691045|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1424|Green||2013-04-02|2013-04-22|NaT||||46.8||1|1|1|1|M|Black||18|Yes|Mother|28262|One Parent: Female|$45,000 to $49,999|||Y|No||Self|General Community||Match Support|M|White||31|28203|Masters Degree|Single|Consultant||0|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503112489|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
500393731|501456966|500347189|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|421|Yellow||2009-03-05|2009-03-09|2010-05-04|Volunteer: Moved|Volunteer: Moved||13.8||1|1|1|1|M|Black||18||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||49|28269||Single|Finance: Accountant||7|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|500393981|31|0|1|31|0|1|10|2|-2||4|2||-2|500000294|-2|0|10|||7462|13|||1|
501194364|501143598|500265628|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1233|Yellow||2008-05-12|2008-05-27|2011-10-12|Volunteer: Moved|Volunteer: Moved||40.5||1|1|1|1|F|Multi-Race (None of the above)||18|No|Mother|28216|Two Parent|$15,000 to $19,999||||Yes||Self|General Community||Enrollment|F|Black||48|28214|Masters Degree|Single|Medical: Doctor, Provider|28207|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011639|501194638|7|0|2|31|0|2|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502861539|502683556|500589768|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|311|Red||2012-01-04|2012-01-10|2012-11-16|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||10.2||1|1|1|1|F|Black||18|No|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Asian||25|28105|Some College|Single|Business: Sales|28134|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502862935|31|0|2|4|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
500186955|500189726|500037840|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3561|Red|Amachi|2004-05-21|2004-05-21|2014-02-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||117||1|1|1|1|F|Black||18|No|Mother|28213|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||55|28226|||Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500188141|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501575246|501546450|500341366|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|915|Yellow||2009-02-16|2009-02-20|2011-08-24|Volunteer: Time constraint|Volunteer: Time constraint||30.1||1|1|1|1|M|Black||18|No|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||41|28212|Bachelors Degree|Married|Education: Teacher|28202|1|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501575542|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7671|13|||1|
502714414|502769005|500577485|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|265|Green||2011-11-11|2011-12-08|2012-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||8.7||1|1|1|1|M|Black||18|No|Mother|28206|One Parent: Female|Less than $10,000|||Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||26|28213|Some College|Single|Business||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502715293|31|0|1|31|0|1|10|2|-2||4|1|500005291|-2||-2|56|1|||7462|13|1208|5|1|
502114586|502081755|500462278|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|368|Green||2010-07-22|2010-08-27|2011-08-30|Volunteer: Time constraint|Volunteer: Time constraint||12.1||1|1|1|1|M|Black||18|No|Mother|28211|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||RTBM|M|White||40|28277|Bachelors Degree|Married|Construction||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502115013|31|0|1|1|0|1|7|2|-2||4|1||-2||-2|6854|8|||7464|9|||1|
502888277|502853546|500593701|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|211|Red|Amachi|2012-01-25|2012-01-31|2012-08-29|Child: Lost interest|Child: Lost interest||6.9||1|1|1|1|M|Black||18|Yes|Mother|28205|One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||63|28269|Bachelors Degree|Married|Business: Sales||9|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502889684|31|0|1|1|0|1|10|2|500003586||4|3|500000294|-2||-2|6854|8|||7464|9|||1|500000294
502588295|502601476|500553687|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|247|Red|Project Big, 2010-2012 OJJDP JJI|2011-09-08|2011-09-27|2012-05-31|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||8.1||1|1|1|1|F|Black||18|No|Mother|28208|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||38|28278|Bachelors Degree|Divorced|Business: Mgt, Admin|28269|1|0|Self|Self|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500011746|502588811|31|0|2|1|0|2|10|2|-2||4|3|500005291|-2||-2|0|10|||7464|9|||1|500004640, 500005291
502973981|503484061|500701296|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|206|Green||2013-06-19|2013-07-02|2014-01-24|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||6.8||1|1|1|1|F|Black||18|No|Mother|28217|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||55|28217|Masters Degree|Widowed|Education: Teacher|28208|0|6|BBBS National Site|Web Link|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500011349|502875571|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501253904|501227814|500336488|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|981|Green||2009-01-28|2009-02-17|2011-10-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||32.2|Y|1|1|1|1|M|White||18|No|Mother|28083|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||38|28115|High School Graduate|Married|Self-Employed, Entrepreneur||6|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501254180|1|0|1|1|0|1|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|
501526673|501361484|500332705|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1687|Yellow|Amachi|2009-01-14|2009-02-25|2013-10-09|Child: Lost interest|Child: Lost interest||55.4||1|1|1|1|F|White||18|Yes||28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||34|28213|Bachelors Degree|Single|Real Estate: Realtor|28215|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500012459|501526965|1|0|2|1|0|2|10|2|500003586||4|2||-2||-2|0|10|||7496|10|||1|500000294
501731841|501182066|500367022|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1547|Red|Amachi|2009-06-02|2009-06-05|2013-08-30|Child: Lost interest|Child: Lost interest||50.8||1|1|1|1|F|Black||18|Yes|Father|28210|One Parent: Male|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||49|28277|Bachelors Degree|Single|Business: Mgt, Admin||4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500008321|501732181|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||46|2|||1|500000294
501831576|502127296|500464171|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|290|Yellow|Amachi|2010-08-04|2010-08-16|2011-06-02|Volunteer: Time constraint|Volunteer: Time constraint||9.5||3|3|1|1|F|Black||18|Yes|Mother|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||37|28105||Single|Education: Teacher||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|501831944|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501831576|501427745|500387626|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|308|Yellow|Amachi|2009-09-24|2009-09-29|2010-08-03|Volunteer: Time constraint|Volunteer: Time constraint||10.1||3|3|1|1|F|Black||18|Yes|Mother|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||33|28211|Bachelors Degree|Single|Medical: Admin|28211|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|501831944|31|0|2|1|0|2|10|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
501831576|502697749|500556209|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|383|Yellow|Amachi|2011-09-20|2011-09-30|2012-10-17|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||12.6||3|3|1|1|F|Black||18|Yes|Mother|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||26|28262|Some College|Single|Retail: Sales||0|6|UNCC|College Partner|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|501831944|31|0|2|1|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||9221|5|1208|5|1|500000294
502102857|502240743|500463814|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|84|Red||2010-08-02|2010-08-05|2010-10-28|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||2.8|Y|2|2|1|1|M|Black||18|No|Mother|28278|One Parent: Female|Unknown||||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||63|28278|Some College|Married|Business: Engineer||25|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500009007|502103284|31|0|1|1|0|1|10|2|-2||4|3|500005291|-2|500000294|-2|0|4|||7464|9|||1|
502102857|502464465|500526162|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|816|Red|2010-2012 OJJDP JJI|2011-03-17|2011-03-25|2013-06-18|Volunteer: Moved|Volunteer: Moved||26.8||2|2|1|1|M|Black||18|No|Mother|28278|One Parent: Female|Unknown||||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||38|28273|Bachelors Degree|Married|Insurance|28202|2|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502103284|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2|500000294, 500004640|-2|0|4|||7446|3|||1|500005291
502499851|502690262|500562789|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1334|Red||2011-10-07|2011-11-11|2015-07-07|Agency: Concern with Volunteer re: child safety|Agency: Concern with Volunteer re: child safety||43.8||1|1|1|1|M|White||18|No|Mother|28210|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||39|28210|Masters Degree|Single|Finance|28106|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|502500300|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
501042226|501089377|500251470|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|434|Green|Amachi|2008-03-11|2008-03-11|2009-05-19|Volunteer: Health|Volunteer: Health||14.3||1|1|1|1|F|White||18|Yes|Mother|28213|One Parent: Female|$10,000 to $14,999||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||60|28227|Bachelors Degree|Married|Medical: Nurse|28269|1|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501042499|1|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||7464|9|||1|500000294
501386394|501818567|500388796|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|541|Yellow||2009-09-28|2009-09-30|2011-03-25|Volunteer: Time constraint|Volunteer: Time constraint||17.8||1|1|1|1|M|Black||18|No|Mother|28227|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||RTBM|M|Black||45|28215||Married|Tech: Research/Design||0|0|Mayfield Memorial|Faith Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501386675|31|0|1|31|0|1|7|2|-2||4|2||-2||-2|34|2|||9212|7|||1|
501309092|501322778|500300356|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1153|Green|Amachi|2008-10-16|2008-10-24|2011-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||37.9||1|1|1|1|M|Black||18|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Black||35|28269|Masters Degree|Single|Tech: Computer/Programmer|28110|3|0|Other|Service Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501309370|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7452|6|||1|500000294
502982301|503442370|500695892|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|806|Green||2013-05-07|2013-05-22|2015-08-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||26.5||1|1|2|2|M|Black||18|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||54|28262|Bachelors Degree|Married|Business||7|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|502983753|31|0|1|31|0|1|10|2|-2||4|1||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|
502319972|502911091|500607368|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1206|Yellow||2012-03-30|2012-04-30|2015-08-19|Volunteer: Moved|Volunteer: Moved||39.6||1|1|1|1|M|Black||18|No|Mother|28214|One Parent: Female|Less than $10,000||||Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||32|28214|Bachelors Degree|Married|Self-Employed, Entrepreneur|29715|0|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502320407|31|0|1|1|0|1|10|2|-2||4|2|500005291|-2||-2|6854|8|||7464|9|||1|
500814240|500981509|500248568|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3248|Green|Amachi|2008-02-27|2008-04-24|NaT||||106.7||1|1|1|1|M|Black||18|Yes|Mother|28212|One Parent: Female|Less than $10,000|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Black||46|28215|Bachelors Degree|Single|Business: Mgt, Admin|28226|0|8|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500814509|31|0|1|31|0|1|10|2|500003586||2|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
502708670|502756331|500584031|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|776|Red||2011-12-05|2011-12-23|2014-02-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||25.5||1|1|1|1|F|Black||18|No|Mother|28209|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||28|28215|Bachelors Degree|Single|Customer Service|28078|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502709557|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||7462|13|||1|
501345385|501375157|500324421|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|742|Green|Amachi|2008-12-09|2008-12-18|2010-12-30|Volunteer: Moved|Volunteer: Moved||24.4||1|1|1|1|M|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|M|White||31|28202|Bachelors Degree|Single|Finance: Banking|28207|0|1|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501345664|31|0|1|1|0|1|5|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||7464|9|||1|500000294
500876120|500830622|500176227|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1063|Red||2007-05-09|2007-05-16|2010-04-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||34.9||1|1|1|1|M|Black||17|No|Mother|28203|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|White||38|28207||Married|Finance: Banking||0|0|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500876387|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7447|3|||1|
501936316|501872326|500428557|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2405|Green||2010-01-21|2010-01-28|2016-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||79||1|1|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||54|28203|||Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017777|501936714|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
502241113|502460114|500538414|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|377|Red||2011-05-25|2011-06-17|2012-06-28|Child: Lost interest|Child: Lost interest||12.4||1|1|2|2|F|Black||17|No|GrandMother|28025|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||43|28027|Masters Degree||Education: Teacher|28027|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|502241544|31|0|2|31|0|2|10|2|-2||4|3||-2|500016374|-2|0|10|||7464|9|||1|
503026286|503259120|500674960|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1487|Red||2013-01-15|2013-01-31|2017-02-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||48.9||1|1|1|1|M|Hispanic||17|No|Mother|28277|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Asian||30|28277|Bachelors Degree|Single|Finance||1|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503027860|3|0|1|4|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502431042|502447496|500515174|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1044|Yellow|2010-2012 OJJDP JJI|2011-02-03|2011-02-10|2013-12-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.3||1|1|1|1|F|Black||17|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||34|28226|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502431483|31|0|2|1|0|2|10|2|-2||4|2|500005291|-2||-2|0|10|||7464|9|||1|500005291
501000843|503106526|500632934|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1072|Red||2012-09-07|2012-10-17|2015-09-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||35.2||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||26|28269|Bachelors Degree|Single|Business|28262|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501001116|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|34|2|||7496|10|||1|
503671116|503672609|500741347|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1140|Green||2014-01-06|2014-01-10|2017-02-23|Volunteer: Moved|Volunteer: Moved||37.5||1|1|1|1|M|White||17|No|GrandMother|28278|One Parent: Female|$20,000 to $24,999||||No||Self|General Community||Match Support|M|White||37|29708|Bachelors Degree|Single|Real Estate: Realtor|28273|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503673077|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501702616|501849169|500405205|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|336|Green||2009-11-03|2009-11-20|2010-10-22|Child/Family: Moved|Child/Family: Moved||11||1|1|1|1|M|Black||17|No|Mother|28134|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||58|29710|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501702954|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
503237270|503022525|500678178|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|237|Green||2013-01-29|2013-02-08|2013-10-03|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.8||1|1|1|1|M|Black||17|No|Mother|28278|One Parent: Female|Less than $10,000|Yes: Retired/Vet||Y|Yes||Self|General Community||RTBM|M|Some Other Race||34|28212|Bachelors Degree|Single|Customer Service|28212|0|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|503239061|31|0|1|41|0|1|7|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
502646551|502262622|500543369|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|369|Green|Project Big|2011-06-29|2011-06-30|2012-07-03|Child/Family: Moved|Child/Family: Moved||12.1||1|1|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|White||34|28210|High School Graduate|Single|Business: Sales|28269|0|8|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502598113|31|0|2|1|0|2|10|2|500004641||4|1|500004640|-2|500004640|-2|0|10|||7464|9|||1|500004640
503013779|501311929|500753159|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Yellow||2014-03-06|2014-03-28|2016-08-26|Volunteer: Time constraint|Volunteer: Time constraint||29||2|2|1|1|F|Multi-race (Black & White)||17|No|Mother|28134|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|Black||49|28269|Masters Degree|Single|Education: Admin|28213|13|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017777|503724588|36|0|2|31|0|2|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1|
503013779|502993965|500618402|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|400|Red||2012-06-07|2012-07-10|2013-08-14|Volunteer: Time constraint|Volunteer: Time constraint||13.1||2|2|1|1|F|Multi-race (Black & White)||17|No|Mother|28134|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|Asian||30|28270|Bachelors Degree|Married|Education|28211|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|503724588|36|0|2|4|0|2|10|2|-2||4|3||-2||-2|0|10|||7462|13|||1|
502874571|501375210|500617142|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|397|Red||2012-05-30|2012-06-27|2013-07-29|Volunteer: Moved|Volunteer: Moved||13||1|1|2|2|F|Hispanic||17|No|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|F|White||30|28202|Bachelors Degree|Single|Tech: Management|28202|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502875969|3|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|4|||7446|3|||1|
501919423|502034798|500442066|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2549|Green|Project Big|2010-03-18|2010-03-24|NaT||||83.7||1|1|1|1|M|Multi-race (Black & Hispanic)||17|No|Mother|28214|One Parent: Female|Unknown||||No|TV|Media|General Community|Project Big|Match Support|M|White||34|28164|Masters Degree||Finance|28210|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501919819|38|0|1|1|0|1|10|2|500004641||2|1|500004640|-2||-2|56|1|||7464|9|||1|500004640
502869635|503099564|500649374|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|646|Red||2012-10-23|2012-11-13|2014-08-21|Volunteer: Moved|Volunteer: Moved||21.2||1|1|1|1|F|Black||17|No|Mother|28206|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|F|Black||34|28210|Bachelors Degree|Single|Business: Marketing||1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502871029|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
502583109|502236275|500551832|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|316|Green|Amachi|2011-08-25|2011-10-26|2012-09-06|Child: Lost interest|Child: Lost interest||10.4||1|1|2|2|F|Black||17|Yes|Mother|28277|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community|Amachi|Match Support|F|White||39|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28217|1|7|Radio|Media|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500008629|502583617|31|0|2|1|0|2|10|2|-2||4|1|500000294|-2|500000294|-2|0|10|||131|1|||1|500000294
500361200|500368628|500085591|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|4013|Green|Cabarrus County|2006-03-21|2006-03-21|NaT||||131.8||2|2|1|1|F|White||17|No|Mother|28027|Two Parent|Unknown||||No||Relative|General Community|Cabarrus County|Match Support|F|White||32|28115|Bachelors Degree|Single|Human Services: Social Worker||0|0|other|College Partner|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|500361450|1|0|2|1|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|0|3|||7670|5|||1|500016374
500378354|501181060|500264206|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3241|Green||2008-05-01|2008-05-01|NaT||||106.5||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$40,000 to $44,999||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||36|28270|Juris Doctorate (JD)|Married|Law: Lawyer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500378596|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|6854|8|||46|2|||1|
501011735|502473442|500528270|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1424|Yellow|2010-2012 OJJDP JJI|2011-03-29|2011-04-11|2015-03-05|Child: Lost interest|Child: Lost interest||46.8||3|3|1|1|F|Black||17||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28215|High School Graduate|Married|Finance: Banking|28255|13|0|Recruitment Event|Workplace Partner|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500012459|500417756|31|0|2|31|0|2|10|2|-2||4|2|500005291|-2||-2|0|10|||7446|3|||1|500005291
501011735|502012852|500456661|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|250|Green||2010-06-14|2010-07-07|2011-03-14|Volunteer: Moved|Volunteer: Moved||8.2||3|3|1|1|F|Black||17||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||44|28204|Bachelors Degree|Divorced|Business: Marketing|28202|9|0|AA Task Force|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|500417756|31|0|2|1|0|2|10|2|-2||4|1|500005291|-2||-2|0|10|||6247|12|||1|
501011735|500728225|500239839|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|642|Green||2008-01-25|2008-01-25|2009-10-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.1||3|3|2|2|F|Black||17||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||33|28208||Single|Finance: Banking||0|3|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500001262|500417756|31|0|2|1|0|2|10|2|-2||4|1|500005291|-2|500000294|-2|0|10|||46|2|||1|
502173821|502264706|500491573|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1380|Red|Amachi|2010-11-05|2010-11-18|2014-08-29|Volunteer: Time constraint|Volunteer: Time constraint||45.3||2|2|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||32|28262|Masters Degree|Single|Finance: Banking|28262|3|11|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502174240|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2|500000294, 500004640|-2|7016|11|||7464|9|||1|500000294
502173821|502057248|500457033|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|131|Green|Amachi|2010-06-16|2010-06-16|2010-10-25|Volunteer: Time constraint|Volunteer: Time constraint||4.3||2|2|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||30|28205||Married|Child/Day Care Worker||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|502174240|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|7016|11|||7464|9|||1|500000294
502725777|502710032|500590950|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1315|Red|Amachi|2012-01-11|2012-01-23|2015-08-30|Volunteer: Moved|Volunteer: Moved||43.2||1|1|1|1|F|Black||17|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||31|28217||Single|Customer Service||0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502726673|31|0|2|31|0|2|10|2|-2||4|3|500000294|-2||-2|34|2|||7464|9|||1|500000294
501861660|501588905|500405168|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|90|Green||2009-11-03|2009-11-06|2010-02-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3||1|1|1|1|F|Hispanic||17||Mother|28273|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||35|28205|Bachelors Degree|Single|Business: Mgt, Admin|28255|4|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009242|501862033|3|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500871269|500798511|500177506|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1358|Green||2007-05-17|2007-05-23|2011-02-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||44.6||1|1|1|1|F|Black||17|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|F|Black||35|28227|Bachelors Degree|Single|Education: Teacher|28227|1|3|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500418342|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502253085|502087592|500467804|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|407|Green||2010-08-27|2010-09-13|2011-10-25|Volunteer: Moved|Volunteer: Moved||13.4||1|1|3|3|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||RTBM|M|Black||45|28262|Bachelors Degree|Married|Business|28202|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500011184|502253517|31|0|1|31|0|1|7|2|-2||4|1||-2|500014505, 500015184|-1|6854|8|||7462|13|||1|
502530688|502166996|500621632|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1425|Yellow||2012-06-25|2012-06-25|2016-05-20|Volunteer: Time constraint|Volunteer: Time constraint||46.8||2|2|3|3|M|Black||17||Mother|28210|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28277|Bachelors Degree|Married|Business||0|0|Michael Baisden|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502531141|31|0|1|31|0|1|10|2|-2||4|2|500005291|-2||-2|0|3|||11272|1|||1|
502530688|502166996|500571794|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|176|Red||2011-10-28|2011-11-16|2012-05-10|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||5.8||2|2|3|3|M|Black||17||Mother|28210|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28277|Bachelors Degree|Married|Business||0|0|Michael Baisden|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502531141|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2||-2|0|3|||11272|1|||1|
500931662|500894084|500193824|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3478|Green||2007-09-05|2007-09-07|NaT||||114.3||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$60,000 to $74,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||58|28270|Bachelors Degree|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|500931932|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1|
500912089|501173565|500262741|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|457|Yellow|Amachi|2008-04-24|2008-05-12|2009-08-12|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||15||1|1|1|1|M|Black||17|Yes|Mother|28208|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|Amachi|Match Support|M|Black||45|28214|Some College|Married|Business: Engineer||14|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500912359|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2||-2|0|10|||2238|7|||1|500000294
502492731|502677685|500557795|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|176|Yellow||2011-09-26|2011-10-05|2012-03-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.8||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||51|28213|Bachelors Degree|Married|Medical|28208|11|0|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502493180|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|6854|8|||7438|1|||1|
502057402|502196301|500461316|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|826|Red||2010-07-16|2010-07-28|2012-10-31|Volunteer: Time constraint|Volunteer: Time constraint||27.1||1|1|1|1|M|White||17|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|White||38|28078|Some College|Married|Military||14|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|502057826|1|0|1|1|0|1|5|2|-2||4|3||-2|500000294|-2|0|4|||7496|10|||1|
503662199|503639494|500741727|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|924|Yellow||2014-01-08|2014-01-17|2016-07-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||30.4||1|1|1|1|M|Black||17|No|Mother|28270|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||32|28226|Bachelors Degree|Married|Consultant|28202|4|4|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|503664159|31|0|1|1|0|1|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1|
502272172|502296220|500516654|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|491|Red|2010-2012 OJJDP JJI|2011-02-10|2011-02-23|2012-06-28|Volunteer: Moved|Volunteer: Moved||16.1||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||29|28277||Single|Student: College||0|0|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502272604|31|0|2|1|0|2|10|2|-2||4|3||-2|500004640|-2|6854|8|||7464|9|||1|500005291
502272172|502965088|500626278|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|741|Yellow||2012-07-26|2012-08-24|2014-09-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.3||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||27|28036|Bachelors Degree|Single|Business|28078|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502272604|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1|
500824205|500850058|500173690|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1099|Yellow||2007-04-24|2007-05-03|2010-05-06|Volunteer: Time constraint|Volunteer: Time constraint||36.1|Y|1|1|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Enrollment|F|White||36|28269|Juris Doctorate (JD)|Married|Law: Lawyer|28202|0|6||Relative|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500824474|31|0|1|1|0|2|5|2|-2||4|2||-2||-2|0|10|||0|11|||1|
503452382|503401641|500700156|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|76|Red||2013-06-11|2013-06-28|2013-09-12|Volunteer: Time constraint|Volunteer: Time constraint||2.5||1|1|1|1|F|Multi-race (Black & White)||17|No|Mother|28269|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||25|28262|Some College|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|503454248|36|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
502255150|502392989|500512287|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2222|Green|Amachi|2011-01-20|2011-02-14|NaT||||73||1|1|1|1|F|Black||17|Yes|Relative: Other|28227|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||34|28212|Masters Degree|Single|Education: Teacher|28216|6|3|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020752|502255582|31|0|2|1|0|2|10|2|500003586||2|1|500000294|-2|500000294, 500004640|-2|0|5|||7464|9|||1|500000294
503745830|503760503|500759184|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|145|Yellow||2014-04-10|2014-04-23|2014-09-15|Volunteer: Moved|Volunteer: Moved||4.8||1|1|1|1|M|Black||17|No|Mother|28206|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|Black||52|28212|Associate Degree|Divorced|Business: Mgt, Admin|60131|1|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018987|503747802|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501955308|501734595|500458840|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|533|Red||2010-06-28|2010-06-30|2011-12-15|Volunteer: Moved|Volunteer: Moved||17.5||1|1|1|1|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||||Yes||School|General Community||RTBM|F|Black||47|28227||Single|Laborer||9|0|New Beginnings Comm.|Faith Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501955706|31|0|2|31|0|2|7|2|-2||4|3||-2||-2|0|4|||9213|7|||1|
502673798|502860952|500590803|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|815|Yellow||2012-01-10|2012-01-30|2014-04-24|Volunteer: Time constraint|Volunteer: Time constraint||26.8||1|1|1|1|M|Black||17|No|Mother|28105|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|White||36|28173|Bachelors Degree|Separated|Business: Mgt, Admin|28110|15|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502674626|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501716763|502112513|500449029|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2380|Red||2010-04-26|2010-05-07|2016-11-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||78.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi, Cabarrus County|Match Support|F|Black||39|28269||Single|Self-Employed, Entrepreneur|28027|7|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500020753|501716992|31|0|2|31|0|2|10|2|-2||4|3|500000294, 500016374|-2|500016374|-2|6854|8|||7458|9|||1|
500186952|500189723|500037836|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|4627|Green|Amachi|2004-07-15|2004-07-15|NaT||||152||1|1|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||73|28203||Married|Self-Employed, Entrepreneur||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500018851|500188132|31|0|2|1|0|2|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502839019|502432390|500674451|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1099|Green||2013-01-11|2013-01-24|2016-01-28|Volunteer: Moved|Volunteer: Moved||36.1||1|1|1|1|M|Black||17|No|Mother|28210|One Parent: Female|$40,000 to $44,999|||Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||32|28203|Bachelors Degree|Single|Business: Mgt, Admin|28202|2|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502840311|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|6854|8|||7496|10|||1|
502076679|502003579|500446859|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|860|Red||2010-04-13|2010-04-30|2012-09-06|Volunteer: Time constraint|Volunteer: Time constraint||28.3||1|1|1|1|M|Black||17|No|Mother|28273|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|White||37|28278|||Finance: Banking||0|0|AA Task Force|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502077103|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|4|||9228|10|||1|
500892049|500765607|500176379|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|876|Green|Amachi|2007-05-10|2007-05-17|2009-10-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||28.8||1|1|1|1|F|Black||17|Yes|GrandMother|28208|One Parent: Female|Unknown||||No||Faith Organization|General Community|Amachi|Match Support|F|Black||62|28278||Married|Unemployed||0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500892316|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||2230|7|||1|500000294
500350138|500188874|500187149|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|904|Green||2007-08-06|2007-08-06|2010-01-26|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29.7||1|1|2|2|M|Black||17||Mother|28025|One Parent: Female|Unknown||||No||Relative|General Community||Match Support|M|Black||41|28027|Some College|Married|Law: Police Officer||5|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500350322|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
500636617|500756919|500151137|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2414|Red||2007-01-04|2007-01-10|2013-08-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||79.3||2|2|1|1|M|Black||17||Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|No|Big|Neighbor/Friend|General Community||Match Support|M|Black||33|28262||Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011746|500636863|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|6854|8|||7464|9|||1|
502555105|502598372|500570292|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|293|Yellow||2011-10-26|2011-11-11|2012-08-30|Child/Family: Moved|Child/Family: Moved||9.6||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|$25,000 to $29,999||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28205|Bachelors Degree|Married|Self-Employed, Entrepreneur|28205|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502555558|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|6854|8|||46|2|||1|
502566108|502562271|500535933|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1203|Green|2010-2012 OJJDP JJI|2011-05-11|2011-05-24|2014-09-08|Volunteer: Time constraint|Volunteer: Time constraint||39.5||1|1|1|1|F|Hispanic||17|No|Mother|28213|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||33|28209||Single|Student: College||0|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500017777|502566562|3|0|2|1|0|2|10|2|-2||4|1|500005291|-2|500005291|-2|0|4|||7464|9|||1|500005291
502702145|502204211|500582836|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1616|Red||2011-11-30|2011-12-21|2016-05-24|Child: Graduated|Child: Graduated||53.1||1|1|2|2|F|Black||17|No|Mother|28083|One Parent: Female|$60,000 to $74,999||||No|Big|Neighbor/Friend|General Community||Match Support|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500020753|502702991|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|6854|8|||7464|9|||1|
503360420|503831013|500765209|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|623|Yellow||2014-06-02|2014-06-20|2016-03-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.5||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|White||31|28262|Bachelors Degree|Single|Tech: Engineer|28262|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503362265|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
502443215|502348503|500510587|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|507|Red|2010-2012 OJJDP JJI|2011-01-12|2011-02-09|2012-06-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||16.7||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black|Other African|50|28215|Bachelors Degree|Divorced|Govt|28208|17|8|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500013709|502443662|31|0|2|31|31|2|10|2|-2||4|3|500005291|-2|500000294|-2|0|10|||7464|9|||1|500005291
502218269|502083213|500461413|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|273|Green|Amachi|2010-07-19|2010-07-30|2011-04-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||9||1|1|1|1|F|Black||17|Yes|Mother|28203|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Enrollment|F|White||27|28262||Single|Service: Restaurant||1|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502218700|31|0|2|1|0|2|5|2|-2||4|1|500000294|-2||-2|7016|11|||7496|10|||1|500000294
501356328|501371070|500315101|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1385|Green||2008-11-14|2008-11-21|2012-09-06|Volunteer: Time constraint|Volunteer: Time constraint||45.5||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||33|28269|Masters Degree|Single|Finance: Banking|28255|0|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501356607|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
502570183|502570153|500534090|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2126|Green|Amachi, Project Big, Project Big AND Amachi|2011-04-30|2011-04-30|2017-02-23|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||69.8||1|1|1|1|F|Black||17|Yes|Mother|28206|Other/Unknown|Unknown||||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||61|28134|Bachelors Degree|Married|Medical: Admin||33|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020910|502570637|31|0|2|31|0|2|10|2|500004772||4|1|500000294, 500004640, 500004901|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|500000294, 500004640, 500004901
502212598|502068243|500457783|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|371|Green|Amachi|2010-06-22|2010-07-22|2011-07-28|Volunteer: Moved|Volunteer: Moved||12.2||2|2|1|1|F|Black||17|Yes|Mother|28215|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||29|28205|Bachelors Degree|Single|Education: Teacher|28208|0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011184|502213028|31|0|2|1|0|2|10|2|-2||4|1|500000294|-2||-2|7016|11|||7464|9|||1|500000294
502212598|502715153|500558562|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|667|Red|Amachi|2011-09-27|2011-10-18|2013-08-15|Volunteer: Moved|Volunteer: Moved||21.9||2|2|1|1|F|Black||17|Yes|Mother|28215|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|White||28|28202|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502213028|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2||-2|7016|11|||7464|9|||1|500000294
501092957|500189785|500277573|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|692|Red||2008-07-14|2008-07-18|2010-06-10|Volunteer: Time constraint|Volunteer: Time constraint||22.7||2|2|2|2|M|Black||17|No|Mother|28027|One Parent: Female|$30,000 to $34,999||||No|Radio|Media|General Community||Match Support|M|Black||51|28269|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|501093231|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|55|1|||7496|10|||1|
501092957|502294662|500484597|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1283|Green||2010-10-22|2010-11-09|2014-05-15|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||42.2||2|2|1|1|M|Black||17|No|Mother|28027|One Parent: Female|$30,000 to $34,999||||No|Radio|Media|General Community||Match Support|M|White||44|28269||Married|Finance: Banking||5|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|501093231|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|55|1|||7459|10|||1|
501224288|500856618|500311410|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1129|Green|Amachi|2008-11-06|2008-11-17|2011-12-21|Volunteer: Moved|Volunteer: Moved||37.1|Y|1|1|2|2|M|Black||17|Yes|Mother|28270|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Enrollment|M|Black||49|28213|Bachelors Degree|Married|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501224558|31|0|1|31|0|1|5|2|500003586||4|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
500887773|500847506|500177121|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1315|Green|Amachi|2007-05-17|2007-05-25|2010-12-30|Volunteer: Time constraint|Volunteer: Time constraint||43.2||1|1|1|1|F|Black||17|Yes|Mother|28206|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Enrollment|F|Black||59|28205||Single|Business: Mgt, Admin|28277|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500888043|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500243491|502919490|500619145|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1710|Green||2012-06-13|2012-07-10|NaT||||56.2||4|4|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|F|Black||47|28269|Bachelors Degree|Single|Law: Paralegal|28202|0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|500188056|31|0|2|31|0|2|10|2|-2||2|1|500000294|-2||-2|0|4|||7464|9|||1|
500243491|500818069|500166029|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1323|Green|Amachi|2007-03-09|2007-03-13|2010-10-26|Volunteer: Moved|Volunteer: Moved||43.5||4|4|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|F|Black||37|28213|Bachelors Degree|Single|Medical: Nurse||2|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188056|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294
500243491|501689965|500505331|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|510|Red|Amachi|2010-12-13|2010-12-16|2012-05-09|Volunteer: Time constraint|Volunteer: Time constraint||16.8||4|4|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|F|Black||35|28270||Single|Business: Mgt, Admin||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500013781|500188056|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294, 500004640|-2|0|4|||7496|10|||1|500000294
501230541|501258738|500276331|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|337|Yellow|Amachi|2008-07-02|2008-07-09|2009-06-11|Volunteer: Lost contact with child/agency Vol: Other Reason|Volunteer: Lost contact with child/agency|Vol: Other Reason|11.1||1|1|1|1|M|Black||17|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|M|Black||35|28208|Bachelors Degree|Single|Business: Clerical|43220|3|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501230817|31|0|1|31|0|1|5|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
502539860|502498837|500529729|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1032|Green|Project Big, 2010-2012 OJJDP JJI|2011-04-06|2011-04-15|2014-02-10|Volunteer: Time constraint|Volunteer: Time constraint||33.9||1|1|1|1|M|Hispanic||17|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Hispanic||33|28270|Associate Degree|Married|Business: Sales||9|0|Other|BBBS Board/Staff|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500017777|502540313|3|0|1|3|0|1|10|2|500004641||4|1|500004640, 500005291|-2|500004640|-2|0|4|||7671|13|||1|500004640, 500005291
502172536|501279665|500475431|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2346|Green||2010-09-30|2010-10-13|NaT||||77.1||1|1|1|1|F|Black||17|No|Mother|28269|Two Parent|Unknown||||Yes||Relative|General Community||Match Support|F|Multi-race (Asian & White)||33|28205|Masters Degree|Married|Finance: Economist|28223|7|0|Newspaper|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502172965|31|0|2|37|0|2|10|2|-2||2|1||-2||-2|0|3|||129|1|||1|
502180719|502184470|500454904|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1385|Green|Amachi, Project Big, Project Big AND Amachi|2010-05-28|2010-06-04|2014-03-20|Volunteer: Moved|Volunteer: Moved||45.5||2|2|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|Black||42|28273|Masters Degree|Divorced|Business: Marketing||1|6|Michael Baisden|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|502181148|31|0|2|31|0|2|10|2|500004772||4|1|500000294|-2|500000294|-2|7016|11|||11146|1|||1|500000294, 500004640, 500004901
502180719|502391505|500755816|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1077|Green||2014-03-20|2014-04-04|NaT||||35.4||2|2|2|2|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|502181148|31|0|2|31|0|2|10|2|500003586||2|1|500000294|-2|500000294|-2|7016|11|||7438|1|||1|
500464540|500821840|500166915|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|671|Red||2007-03-14|2007-03-23|2009-01-22|Volunteer: Moved|Volunteer: Moved||22||1|1|1|1|F|Black||17||Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||32|28209|Bachelors Degree|Married|Unknown||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500187629|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501133304|501147729|500249703|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|562|Green|Amachi|2008-03-03|2008-03-26|2009-10-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||18.5||1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||37|28105|Bachelors Degree|Married|Construction|28273|3|5|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501115202|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502551092|502366844|500536172|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1623|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-05-12|2011-05-20|2015-10-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||53.3||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||42|28210||Single|Business: Human Resources||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502551545|31|0|2|1|0|2|10|2|-2||4|2|500004640, 500005291|-2||-2|0|4|||10326|3|460|3|1|500004640, 500005291
501809543|501333516|500375191|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|34|Green||2009-07-23|2009-08-07|2009-09-10|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||1.1||1|1|1|1|F|Multi-race (Black & White)||17|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Enrollment|F|White||52|28269|Associate Degree|Married|Business: Clerical|28075|0|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501809896|36|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186248|501470065|500340015|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|872|Yellow||2009-02-10|2009-03-09|2011-07-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.6||3|3|1|1|F|Black||17||Mother|28214|Other/Unknown|Unknown||||No||Self|General Community||Enrollment|F|Black||40|28216||Single|Finance: Banking||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|500187843|31|0|2|31|0|2|5|2|-2||4|2||-2||-2|0|10|||7462|13|||1|
502670076|501391123|500745456|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1102|Green|Cabarrus County|2014-01-28|2014-03-10|NaT||||36.2||2|2|3|3|F|Black||17|No|Mother|28083|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|Black||41|28027|PHD|Single|Medical: Doctor, Provider|28075|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502670904|31|0|2|31|0|2|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
502670076|502655392|500552412|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|603|Yellow||2011-08-30|2011-10-12|2013-06-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.8||2|2|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|Black||31|29223|||Human Services: Youth Worker||0|0|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502670904|31|0|2|31|0|2|10|2|-2||4|2|500000294, 500016374|-2||-2|0|10|||7459|10|||1|
503015906|503041890|500678458|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|93|Green||2013-01-30|2013-02-19|2013-05-23|Child: Lost interest|Child: Lost interest||3.1||1|1|2|2|M|White||17|No|Mother|28027|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|M|White||60|28027|Bachelors Degree|Separated|Insurance|28262|24|0|Local Radio|Media|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500015820|503017438|1|0|1|1|0|1|10|2|-2||4|1||-2|500016374|-2|0|10|||7437|1|||1|
502290600|502450688|500516671|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|437|Yellow|Amachi|2011-02-10|2011-02-18|2012-04-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.4||1|1|1|1|M|Black||17|Yes|Mother|28216|One Parent: Female|Unknown||||Yes|Radio|Media|General Community|Amachi|Enrollment|M|Some Other Race||52|28031|Some College|Married|Govt|28031|17|0|Other|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502291037|31|0|1|41|0|1|5|2|-2||4|2|500000294|-2||-2|55|1|||7452|6|||1|500000294
502828146|502860825|500607619|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|760|Red||2012-04-02|2012-04-30|2014-05-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25||1|1|1|1|M|Black||17|No|Father|28214|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|Black||37|28278|Bachelors Degree|Single|Unknown||0|0|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502829415|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||9229|13|||1|
501099857|500801514|500243554|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|764|Red||2008-02-07|2008-02-19|2010-03-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25.1||1|1|1|1|F|Black||17||Mother|28216|One Parent: Female|Unknown||||No||Service Organization|General Community||Match Support|F|Black||38|28216||Single|Finance: Banking||5|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501100131|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|11|||46|2|||1|
502745717|502712044|500583497|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|413|Red||2011-12-01|2012-01-12|2013-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||13.6||1|1|1|1|F|Multi-race (Black & White)||17|No|Mother|28278|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|F|Asian||34|28278|Bachelors Degree|Single|Govt|28226|0|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502746625|36|0|2|4|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500938154|501446421|500323753|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2985|Green||2008-12-08|2009-01-12|NaT||||98.1||2|2|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||32|28208|Associate Degree|Single|Service: Restaurant|28211|4|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|500938424|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502188863|502288935|500498784|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1035|Red|Project Big|2010-11-23|2010-12-31|2013-10-31|Volunteer: Moved|Volunteer: Moved||34||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|M|Some Other Race||30|28202|Some College|Single|Tech: Support, Writing|28210|0|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502189292|31|0|1|41|0|1|10|2|-2||4|3|500004640|-2|500004640|-2|0|10|||46|2|||1|500004640
502145270|500189131|500462648|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|453|Green||2010-07-26|2010-07-30|2011-10-26|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||14.9||1|1|2|2|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|F|Black||39|28262|Masters Degree|Single|Human Services: Psychologist||3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502145699|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|8|||7496|10|||1|
500336002|500801056|500490281|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|488|Red|Amachi|2010-11-03|2010-11-29|2012-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16||4|5|2|3|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||||No||School|General Community|Amachi|Match Support|F|White||33|28202||Single|Business: Marketing||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013709|500293247|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|0|4|||7464|9|||1|500000294
502961272|503009515|500614268|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|618|Yellow|Amachi|2012-05-11|2012-05-21|2014-01-29|Child/Family: Moved|Child/Family: Moved||20.3||1|1|1|1|F|White||17|Yes|Mother|28205|Grandparents|$25,000 to $29,999||||Yes||Self|General Community|Amachi|Match Support|F|White||62|28299|Some College|Divorced|Business: Sales||1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502962447|1|0|2|1|0|2|10|2|-2||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
500911385|501413944|500326312|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|662|Red||2008-12-12|2009-01-02|2010-10-26|Child/Family: Moved|Child/Family: Moved||21.7||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|$40,000 to $44,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||45|28262|Bachelors Degree||Finance: Banking|28078|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|500911655|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
501300013|500188952|500281427|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1356|Green|Amachi|2008-08-11|2008-08-14|2012-05-01|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||44.6||2|2|2|2|F|Black||17|Yes|GrandMother|28273|Grandparents|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|Black||40|28277|Associate Degree|Single|Unknown||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500561354|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2||-2|7294|13|||7464|9|||1|500000294
500970495|500965698|500285645|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3102|Yellow||2008-09-03|2008-09-10|2017-03-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||101.9||3|3|1|1|F|Black||17|No|Mother|28227|One Parent: Female|$35,000 to $39,999||||No|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black|Other African|44|28212||Single|Consultant||1|5|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500970766|31|0|2|31|31|2|10|2|-2||4|2||-2||-2|7294|13|||46|2|||1|
503664796|503674336|500744967|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|112|Green||2014-01-27|2014-01-31|2014-05-23|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.7||1|1|1|1|M|Black||17|No|Mother|28227|One Parent: Female|$45,000 to $49,999|||Y|Yes||Self|General Community||Match Support|M|White||51|28210|Bachelors Degree|Domestic Partner|Arts, Entertainment, Sports|28210|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002334|503666756|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500970264|502250629|500478922|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|964|Red|Amachi|2010-10-11|2010-10-27|2013-06-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.7||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|||Y|No|Other|Faith Organization|General Community|Amachi|Enrollment|M|Black||44|28269|Some High School|Single|Insurance||0|2|100 Men in 100 Days|Fraternity/Sorority|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|500970535|31|0|1|31|0|1|5|2|500003586||4|3|500000294|-2|500000294|-2|5635|9|||12183|14|1209|1|1|500000294
500970267|502084649|500468192|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2360|Green|Amachi|2010-08-31|2010-09-29|NaT||||77.5||1|1|1|1|F|Black||17|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||61|28204||Divorced|Self-Employed, Entrepreneur||0|0|Billboard|Media|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|500970535|31|0|2|1|0|2|10|2|500003586||2|1|500000294|-2|500000294|-2|5635|9|||125|1|||1|500000294
502571727|502769619|500586830|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1882|Green||2011-12-14|2012-01-13|2017-03-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||61.8||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|Black||45|28207|Masters Degree|Married|Tech: Management|28081|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502572181|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
500958307|500876132|500193868|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3466|Green|Amachi, Cabarrus County|2007-09-05|2007-09-19|NaT||||113.9|Y|1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$40,000 to $44,999|||Y|No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|Black||62|28213||Married|Finance: Economist||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|500958577|31|0|1|31|0|1|10|2|500003586||2|1|500000294, 500016374|-2|500000294, 500016374|-2|5635|9|||2238|7|||1|500000294, 500016374
501230772|501157134|500261012|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|833|Green|Amachi|2008-04-15|2008-04-22|2010-08-03|Volunteer: Moved|Volunteer: Moved||27.4||1|1|1|1|F|Black||17|Yes|Mother|28214|Two Parent|Unknown||||Yes||School|General Community||Match Support|F|White||34|28211|Associate Degree|Single|Business: Clerical||0|1|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501231048|31|0|2|1|0|2|10|2|500003586||4|1||-2||-2|0|4|||2238|7|||1|500000294
501257717|503426906|500700329|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|69|Red||2013-06-12|2013-06-22|2013-08-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||2.3||2|2|1|1|F|Black||17|No|GrandMother|28203|Grandparents|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|Black||37|28134|Masters Degree|Single|Business: Mgt, Admin|28202|0|2|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|501257994|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501257717|500839705|500271936|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1593|Green||2008-06-10|2008-06-20|2012-10-30|Volunteer: Time constraint|Volunteer: Time constraint||52.3||2|2|2|2|F|Black||17|No|GrandMother|28203|Grandparents|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|White||31|28204|Bachelors Degree|Single|Finance: Banking||0|3|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008321|501257994|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
503417576|503594017|500730510|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|751|Red||2013-11-13|2013-12-09|2015-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.7||1|1|1|1|F|White||17|No|Father|28269|Two Parent|$100,000 to $124,999|||Y|No||Relative|General Community||Match Support|F|White||29|28205|Some College|Single|Business: Mgt, Admin|29707|3|10|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|503419440|1|0|2|1|0|2|10|2|-2||4|3||-2|500000294|-2|0|3|||7464|9|||1|
503255669|500188812|500703771|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1034|Yellow||2013-07-16|2013-07-26|2016-05-25|Child: Lost interest|Child: Lost interest||34||1|1|2|3|M|Black||17|No|Mother|28216|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|Black||40|28202|Bachelors Degree|Single|Consultant|28281|4|5|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|0|1|0|1|277|60|598|500000170|500013781|503257474|31|0|1|31|0|1|10|2|-2||4|2||-2|500000294|-2|0|10|||2238|7|||1|
500938169|501370307|500320339|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|400|Green||2008-11-25|2008-12-08|2010-01-12|Volunteer: Time constraint|Volunteer: Time constraint||13.1||1|1|1|1|M|Multi-Race (None of the above)||17|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|No|BBBS National Site|Web Link|General Community||Enrollment|M|Asian||39|28207|Masters Degree|Single|Business: Sales|94085|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500981706|7|0|1|4|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
502666840|502872585|500594266|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|376|Red||2012-01-27|2012-02-17|2013-02-27|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.4||1|1|1|1|M|Black||17|No|Mother|28277|One Parent: Female|$20,000 to $24,999||||Yes|Arby's|Workplace Partner/Business|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||49|28173|Bachelors Degree|Single|Insurance|28210|21|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502667667|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2||-2|3394|14|||7496|10|||1|
500791785|500785783|500159822|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1309|Green|Amachi|2007-02-13|2007-02-13|2010-09-14|Volunteer: Moved|Volunteer: Moved||43||1|1|1|1|M|Multi-Race (None of the above)||17|Yes|Mother|28081|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|M|Black||42|28075||Married|Finance: Banking|28255|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500002335|500766037|7|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|3|||2238|7|||1|500000294
502674024|502660051|500581910|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1623|Green||2011-11-28|2011-12-07|2016-05-17|Child: Lost interest|Child: Lost interest||53.3||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Sales||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502674852|31|0|2|1|0|2|10|2|-2||4|1|500005291|-2||-2|0|10|||7496|10|||1|
502696388|502609046|500553973|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|178|Green|2010-2012 OJJDP JJI|2011-09-09|2011-09-27|2012-03-23|Volunteer: Moved|Volunteer: Moved||5.8||1|1|1|1|F|Black||17|No|Mother|28212|One Parent: Female|Unknown|||Y|Yes||Self|General Community||RTBM|F|White||28|28105|Masters Degree|Single|Medical: Healthcare Worker|28078|0|1|Recruitment Event|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502697233|31|0|2|1|0|2|7|2|-2||4|1||-2||-2|0|10|||7460|12|||1|500005291
501670169|501466072|500379969|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|917|Green||2009-08-19|2009-09-30|2012-04-04|Volunteer: Time constraint|Volunteer: Time constraint||30.1||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|F|Black||32|28269||Single|Consultant|28209|0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|501670507|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
501157075|502978065|500619009|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1300|Yellow||2012-06-12|2012-06-30|2016-01-21|Child: Lost interest|Child: Lost interest||42.7||3|4|1|1|F|Black||17||Relative: Other|28206|Grandparents|Unknown||||Yes||School|General Community|Amachi|Match Support|F|Black||37|28215|Masters Degree|Single|Human Services: Social Worker||2|0|Self|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500020752|501157349|31|0|2|31|0|2|10|2|-2||4|2|500000294|-2||-2|0|4|||7464|9|||1|
501157075|502261758|500467512|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|632|Red|Amachi|2010-08-26|2010-08-30|2012-05-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.8||3|4|2|2|F|Black||17||Relative: Other|28206|Grandparents|Unknown||||Yes||School|General Community|Amachi|Match Support|F|Black||34|28216|Masters Degree|Single|Business|28202|8|7|Self|Self|Big|General Site|mentor2.0, mentor2.0 2014|Match Support|0|1|1|0|277|60|598|500000170|500008629|501157349|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500014505, 500014506|-1|0|4|||7464|9|||1|500000294
503804225|503881040|500773105|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|501|Red||2014-08-21|2014-09-15|2016-01-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.5||1|1|1|1|F|Black||17|No|Mother|28208|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Multi-race (Black & Hispanic)||59|28216|Some College|Divorced|Law: Legal Secretary|28202|14|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503805695|31|0|2|38|0|2|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
501309634|501046221|500281317|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3107|Green|Amachi|2008-08-11|2008-09-12|NaT||||102.1||1|1|1|1|F|Black||17|Yes|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||46|27704|Associate Degree|Divorced|Medical: Admin||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500008321|501309912|31|0|2|31|0|2|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||7462|13|||1|500000294
503448711|503576769|500742906|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|631|Green||2014-01-15|2014-02-26|2015-11-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.7||1|1|1|1|M|Black||17|No|Mother|28226|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||34|28210|Masters Degree|Married|Real Estate: Realtor|28202|2|3|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|503450577|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
503331975|503796877|500769464|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|104|Red||2014-07-14|2014-07-25|2014-11-06|Child: Lost interest|Child: Lost interest||3.4||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||34|28269|Bachelors Degree|Married|Medical: Healthcare Worker|28209|0|4|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500012459|503333815|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500736177|502513250|500536659|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|555|Red|2010-2012 OJJDP JJI|2011-05-17|2011-05-25|2012-11-30|Volunteer: Time constraint|Volunteer: Time constraint||18.2||2|3|1|1|F|Black||17||Mother|28269|One Parent: Female|Unknown||||No||School|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||38|28206|Bachelors Degree|Single|Finance|28255|2|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|500710887|31|0|2|1|0|2|5|2|-2||4|3|500005291|-2||-2|0|4|||7464|9|||1|500005291
500843862|501098883|500272053|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|345|Green|Amachi|2008-06-11|2008-06-25|2009-06-05|Vol: Other Reason|Vol: Other Reason||11.3||2|2|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|No|TV|Media|General Community|Amachi|Enrollment|F|Multi-race (Black & Hispanic)||36|28202|Bachelors Degree|Single|Finance: Banking||0|10|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500844129|31|0|2|38|0|2|5|2|500003586||4|1|500000294|-2||-2|56|1|||46|2|||1|500000294
501582592|501783333|500373122|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|371|Red||2009-07-08|2009-08-20|2010-08-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.2||1|1|1|1|M|Multi-Race (None of the above)||17|No|Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Hispanic||34|28227|||Insurance||2|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501582912|7|0|1|3|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501796006|503531528|500705837|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|258|Yellow||2013-08-05|2013-08-23|2014-05-08|Child: Lost interest|Child: Lost interest||8.5||3|3|1|1|F|Black||17|No|Mother|28031|Two Parent|Unknown|||Y|Yes||School|General Community||Match Support|F|Black||48|28037|Some College|Married|Law: Paralegal|28036|6|0|Newspaper|Media|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500015820|501489205|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|4|||129|1|||1|
501796006|501621517|500396069|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|777|Green||2009-10-16|2009-11-03|2011-12-20|Volunteer: Time constraint|Volunteer: Time constraint||25.5||3|3|1|1|F|Black||17|No|Mother|28031|Two Parent|Unknown|||Y|Yes||School|General Community||Match Support|F|White||37|28078|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|501489205|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
501796006|502469185|500595418|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|398|Yellow||2012-02-01|2012-02-17|2013-03-21|Volunteer: Time constraint|Volunteer: Time constraint||13.1||3|3|1|1|F|Black||17|No|Mother|28031|Two Parent|Unknown|||Y|Yes||School|General Community||Match Support|F|White||37|28031|Masters Degree|Married|Finance: Banking|28202|7|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|501489205|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|4|||7462|13|||1|
502885468|502954219|500610806|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1781|Green||2012-04-19|2012-04-30|NaT||||58.5||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Black||47|28227|Bachelors Degree|Married|Tech: Engineer||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502886874|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
500383688|500358123|500085796|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1342|Green||2006-03-23|2006-03-23|2009-11-24|Volunteer: Time constraint|Volunteer: Time constraint||44.1||1|1|1|1|F|Black||17||Mother|28262|One Parent: Female|Unknown||||No||School|General Community||Enrollment|F|Native Hawaiian or Other Pacific Islander||44|28209|Bachelors Degree|Single|Business: Mgt, Admin|28202|10|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500383938|31|0|2|5|0|2|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502941572|502884011|500608269|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|371|Green|Amachi|2012-04-05|2012-04-16|2013-04-22|Child/Family: Moved|Child/Family: Moved||12.2||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||44|28269|PHD|Single|Medical|64506|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502942998|31|0|2|1|0|2|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
502371558|502528355|500568298|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1963|Green||2011-10-20|2011-10-31|NaT||||64.5||1|1|2|2|M|Black||17|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||30|28202|Bachelors Degree|Married|Business: Engineer|28202|1|9|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502371997|31|0|1|1|0|1|10|2|-2||2|1|500000294, 500005291|-2||-2|0|10|||132|8|||1|
502275241|502394690|500521625|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1669|Green|Amachi|2011-03-03|2011-03-21|2015-10-15|Child: Lost interest|Child: Lost interest||54.8||1|1|1|1|F|Black||17|No|Mother|28262|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||26|28031|Bachelors Degree|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|502275673|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7496|10|||1|500000294
502671420|502938924|500604987|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|356|Red||2012-03-19|2012-04-13|2013-04-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.7||1|1|1|1|M|Black||17|No|Mother|28210|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Multi-race (Black & White)||33|28277|Associate Degree|Married|Tech: Computer/Programmer||6|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502672248|31|0|1|36|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502129650|502598777|500646243|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1602|Green|Cabarrus County|2012-10-16|2012-10-26|NaT||||52.6||2|2|2|2|F|Black||17|No|GrandMother|28027|Grandparents|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|Black||42|28213|Bachelors Degree|Single|Finance: Banking|28202|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502130079|31|0|2|31|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
502129650|501733783|500502959|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|650|Yellow||2010-12-07|2010-12-17|2012-09-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.4||2|2|1|1|F|Black||17|No|GrandMother|28027|Grandparents|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|Black||29|28027|||Customer Service||0|0||High School Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502130079|31|0|2|31|0|2|10|2|-2||4|2|500016374|-2||-2|0|10|||0|4|||1|
502224918|502448424|500533984|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|155|Red|2010-2012 OJJDP JJI|2011-04-29|2011-05-10|2011-10-12|Volunteer: Time constraint|Volunteer: Time constraint||5.1||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|M|Asian||31|28202||Single|Law: Lawyer|28202|2|4|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014, Project Big|RTBM|0|1|1|0|277|60|598|500000170|500011639|502225349|31|0|1|4|0|1|7|2|-2||4|3|500005291|-2|500004640, 500014506|-1|0|10|||7671|13|||1|500005291
501386307|501294991|500307024|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|515|Yellow||2008-10-29|2008-11-17|2010-04-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.9||1|1|1|1|M|Black||17|No|Mother|28217|One Parent: Female|Unknown||||Yes||Relative|General Community||Enrollment|M|White||42|28277|Masters Degree|Married|Business: Sales|28277|0|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501386588|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|3|||7464|9|||1|
500948385|500885771|500187434|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1961|Yellow||2007-08-08|2007-08-28|2013-01-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||64.4||1|1|1|1|F|Black||17|No|Mother|28214|One Parent: Female|$30,000 to $34,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Asian|Chinese|32|28216|||Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|500948655|31|0|2|4|16|2|10|2|-2||4|2||-2||-2|34|2|||46|2|||1|
502139829|502178005|500462499|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1092|Red||2010-07-23|2010-08-12|2013-08-08|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.9||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||30|28226|Masters Degree|Single|Finance: Accountant||0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502140258|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501725162|501833178|500394157|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2542|Green||2009-10-13|2009-10-29|2016-10-14|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||83.5||1|1|1|1|M|Multi-race (Black & Asian)||17|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||32|28215|||Business: Engineer|28273|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|501724831|39|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502645484|502291769|500544311|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|502|Green|Project Big|2011-06-30|2011-06-30|2012-11-13|Child/Family: Moved|Child/Family: Moved||16.5||1|1|1|1|F|Black||17||Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||26|28223||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502508948|31|0|2|31|0|2|10|2|-2||4|1|500004640, 500005291|-2||-2|0|10|||7464|9|||1|500004640
501441404|501550442|500336614|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|302|Yellow||2009-01-28|2009-02-03|2009-12-02|Child/Family: Moved|Child/Family: Moved||9.9||1|1|1|1|F|Multi-race (Hispanic & White)||17|No|Mother|28120|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Multi-race (Hispanic & White)||34|28202|Juris Doctorate (JD)|Married|Law: Lawyer|28202|1|2|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501441689|35|0|2|35|0|2|10|2|-2||4|2||-2||-2|0|10|||7671|13|||1|
503124706|503609606|500755317|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|666|Green||2014-03-18|2014-03-31|2016-01-26|Volunteer: Moved|Volunteer: Moved||21.9||1|1|1|1|M|Black||17|No|Mother|28226|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|Multi-race (Black & White)||29|28215|Some College|Married|Student: College|28223|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503126373|31|0|1|36|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502526965|502881104|500606886|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1808|Green||2012-03-28|2012-04-03|NaT||||59.4||1|1|1|1|M|Black||17|No|Mother|28278|Two Mothers|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||32|28278|Bachelors Degree|Single|Medical|28208|3|5|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502527418|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||17161|11|||1|
500186901|500189670|500037782|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|2166|Green|Amachi|2005-01-24|2005-01-24|2010-12-30|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||71.2||1|1|1|1|F|Black||17||Mother|28216|One Parent: Female|Unknown|||Y|No|Brochure|Media|General Community|Amachi|Enrollment|F|Black||82|28215|Some High School|Widowed|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500187992|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|51|1|||2238|7|||1|500000294
502431187|503015009|500627361|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1238|Yellow||2012-08-03|2012-08-17|2016-01-07|Volunteer: Time constraint|Volunteer: Time constraint||40.7||2|2|1|1|F|Black||17|No|GrandMother|28208|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|RTBM|F|White||41|28105|Bachelors Degree|Divorced|Business|28112|1|3|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502431630|31|0|2|1|0|2|7|2|-2||4|2|500005291|-2||-2|0|5|||46|2|||1|
502431187|502616530|500545377|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|274|Red|2010-2012 OJJDP JJI|2011-07-13|2011-07-21|2012-04-20|Volunteer: Time constraint|Volunteer: Time constraint||9||2|2|1|1|F|Black||17|No|GrandMother|28208|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|RTBM|F|Black||27|28262|Some College|Single|Retail: Sales||0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502431630|31|0|2|31|0|2|7|2|-2||4|3|500005291|-2||-2|0|5|||7464|9|||1|500005291
503546374|503890372|500774577|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|178|Yellow|PERL 2014-2016|2014-09-04|2014-09-29|2015-03-26|Child: Severity of challenges|Child: Severity of challenges||5.8||1|1|2|2|M|Black||17|No|Mother|28216|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|M|Asian||33|28204|Bachelors Degree|Married|Business: Engineer|28007|3|9|Man Up Campaign|Media|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500015820|503548249|31|0|1|4|0|1|10|2|-2||4|2|500014681|-2|500000294, 500014681|-2|0|4|||17101|1|||1|500014681
500934906|500859806|500186448|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2023|Red|Amachi|2007-07-30|2007-07-31|2013-02-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||66.5||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Less than $10,000|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||52|28216|Bachelors Degree|Married|Tech: Engineer||13|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500011349|500935173|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|5635|9|||2238|7|||1|500000294
500787601|500189612|500153750|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1324|Yellow||2007-01-23|2007-01-24|2010-09-09|Volunteer: Moved|Volunteer: Moved||43.5||1|1|2|2|M|Black||17||Mother|28216|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|Black||47|28273||Married|Arts, Entertainment, Sports||0|6|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500010765|500787869|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7671|13|||1|
501379296|501296492|500297204|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1043|Green||2008-10-09|2008-10-15|2011-08-24|Child/Family: Moved|Child/Family: Moved||34.3||1|1|1|1|M|Black||17||Mother|28227|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||33|28211|Bachelors Degree|Single|Unemployed||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501161168|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500870948|501367743|500331371|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|95|Green|Amachi|2009-01-08|2009-01-12|2009-04-17|Vol: Changed School or Site|Vol: Changed School or Site||3.1||3|3|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||62|28105|Bachelors Degree|Married|Business: Mgt, Admin|28086|0|11|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501616314|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
500870948|501559777|500358785|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|678|Green|Amachi|2009-04-21|2009-05-22|2011-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||22.3||3|3|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|F|White||38|28204|Bachelors Degree|Single|Consultant|28036|0|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501616314|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
500271303|501291358|500354049|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2286|Green|Amachi|2009-04-01|2009-04-30|2015-08-03|Volunteer: Time constraint|Volunteer: Time constraint||75.1||2|2|1|1|F|Black||17|Yes|Mother|28227|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||31|28204|Bachelors Degree|Single|Business: Engineer|28269|0|2|TV|Media|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500011349|500271368|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||130|1|||1|500000294
501771253|501322818|500383563|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|569|Yellow||2009-09-09|2009-09-29|2011-04-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||18.7||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||34|28269|Bachelors Degree|Single|Medical: Nurse|28054|3|6|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500009007|501741899|31|0|2|31|0|2|5|2|500003586||4|2||-2|500000294|-2|0|10|||7462|13|||1|
502106926|503230500|500686913|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|555|Green||2013-03-08|2013-03-18|2014-09-24|Child/Family: Moved|Child/Family: Moved||18.2||2|2|1|1|M|Black||17|No|Mother|28031|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||53|28036|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0||Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502107353|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||0|11|||1|
502106926|502072628|500453665|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|765|Red||2010-05-20|2010-05-25|2012-06-28|Volunteer: Time constraint|Volunteer: Time constraint||25.1||2|2|1|1|M|Black||17|No|Mother|28031|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||32|28031||Single|Govt||0|0|AA Task Force|Special Event|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502107353|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||11098|8|||1|
500724632|500803551|500164708|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3662|Green||2007-03-02|2007-03-07|NaT||||120.3||1|1|1|1|F|Black||17||Mother|28213|One Parent: Female|Less than $10,000|||Y|No||School|General Community||Match Support|F|Black||32|28214|Bachelors Degree|Married|Architect|28270|0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|500724899|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|4|||46|2|||1|
500826596|501799403|500375650|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|607|Green||2009-07-27|2009-08-07|2011-04-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.9||3|3|1|1|M|Black||17|No|Mother|28226|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|M|Black||35|28226|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|500826861|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|5|||7464|9|||1|
500826596|502549323|500544976|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|872|Yellow|2010-2012 OJJDP JJI|2011-07-11|2011-07-28|2013-12-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.6||3|3|1|1|M|Black||17|No|Mother|28226|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|M|Black||29|28226|Some College|Single|Customer Service|28210|2|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011349|500826861|31|0|1|31|0|1|10|2|-2||4|2||-2|500000294|-2|0|5|||7464|9|||1|500005291
501292079|501519897|500323243|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1680|Green|Amachi|2008-12-05|2008-12-11|2013-07-18|Child: Lost interest|Child: Lost interest||55.2||1|1|1|1|F|Black||17|Yes|GrandMother|28214|Grandparents|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|F|White||31|28203|Bachelors Degree|Single|Consultant|28204|0|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|501292357|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|7294|13|||7464|9|||1|500000294
501312033|500881761|500280688|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|440|Yellow||2008-08-05|2008-08-12|2009-10-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.5||2|2|1|1|F|Black||17|No|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||38|28277|Bachelors Degree|Single|Business: Sales|60093|5|10|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501312311|31|0|2|1|0|2|10|2|-2||4|2|500000294|-2||-2|0|10|||7464|9|||1|
501312033|502053746|500452835|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|999|Red||2010-05-14|2010-06-04|2013-02-27|Child: Lost interest|Child: Lost interest||32.8||2|2|1|1|F|Black||17|No|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||35|28226|||Customer Service||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500015820|501312311|31|0|2|31|0|2|10|2|-2||4|3|500000294|-2||-2|0|10|||7464|9|||1|
501444237|502981694|500623203|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|188|Red||2012-07-09|2012-07-27|2013-01-31|Child: Lost interest|Child: Lost interest||6.2||3|3|1|1|M|Black||17||GrandMother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|Black||59|28213|Associate Degree|Single|Transport: Driver|28216|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500015820|501444522|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
501444237|502183206|500461448|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|441|Red||2010-07-19|2010-07-29|2011-10-13|Volunteer: Time constraint|Volunteer: Time constraint||14.5||3|3|1|1|M|Black||17||GrandMother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|Black||36|28213|Associate Degree|Single|Retail: Sales||3|6|Michael Baisden|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011639|501444522|31|0|1|31|0|1|10|2|-2||4|3||-2|500000294|-2|0|10|||11146|1|||1|
501444237|501358303|500326259|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|432|Green||2008-12-12|2008-12-14|2010-02-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.2||3|3|1|1|M|Black||17||GrandMother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||32|28262|High School Graduate|Single|Student: College||0|0|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500009242|501444522|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
502124485|501905673|500689671|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1452|Green||2013-03-25|2013-03-25|NaT||||47.7||2|2|2|2|F|Black||17|No|Mother|28217|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||34|28216||Single|Medical: Healthcare Worker||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502142970|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|4|||7496|10|||1|
502124485|502066586|500454581|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|459|Green||2010-05-26|2010-05-28|2011-08-30|Volunteer: Time constraint|Volunteer: Time constraint||15.1||2|2|1|1|F|Black||17|No|Mother|28217|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||32|28206||Single|Medical: Nurse||0|0|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502142970|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7438|1|||1|
502589869|501833131|500538612|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|102|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-05-26|2011-06-30|2011-10-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.4||2|2|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||43|28262||Married|Medical: Nurse|28208|0|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502590381|31|0|2|31|0|2|10|2|500004641||4|2|500004640, 500005291|-2|500004640|-2|0|4|459|3|10326|3|460|3|1|500004640, 500005291
502589869|502701252|500582617|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1429|Green|Project Big|2011-11-29|2011-11-30|2015-10-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||46.9||2|2|1|1|F|Black||17||Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28205|Bachelors Degree|Married|Business|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017777|502590381|31|0|2|1|0|2|10|2|500004641||4|1|500004640, 500005291|-2|500000294|-2|0|4|459|3|7496|10|||1|500004640
502907527|502996593|500624606|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|820|Yellow||2012-07-18|2012-08-23|2014-11-21|Volunteer: Moved|Volunteer: Moved||26.9||1|1|1|1|M|Black||17|Yes|Mother|28212|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||55|28202|Associate Degree|Married|Business||30|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502908938|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2||-2|0|10|||7464|9|||1|
502233625|502228626|500465112|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|160|Green||2010-08-10|2010-08-13|2011-01-20|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||5.3||3|3|1|1|F|Multi-race (Hispanic & White)||17|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||31|28269|Bachelors Degree|Single|Finance||3|0|Self|Self|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500011639|502234056|35|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502233625|503081963|500628685|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|424|Red||2012-08-15|2012-08-24|2013-10-22|Child/Family: Moved|Child/Family: Moved||13.9||3|3|1|1|F|Multi-race (Hispanic & White)||17|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||30|28209|Associate Degree|Single|Medical: Nurse|28210|2|6|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500011746|502234056|35|0|2|1|0|2|10|2|-2||4|3||-2|500000294|-2|0|10|||7464|9|||1|
502233625|502381327|500519189|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|485|Yellow|2010-2012 OJJDP JJI|2011-02-22|2011-03-02|2012-06-29|Volunteer: Moved|Volunteer: Moved||15.9||3|3|1|1|F|Multi-race (Hispanic & White)||17|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||29|28262|Bachelors Degree|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502234056|35|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|500005291
502591943|502757658|500593218|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|214|Red||2012-01-23|2012-01-29|2012-08-30|Child: Family structure changed|Child: Family structure changed||7||1|1|1|1|F|White||17|No|Mother|28278|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28209|Bachelors Degree|Single|Business: Mgt, Admin|28210|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502592460|1|0|2|1|0|2|10|2|||4|3|500005291|-2||-2|0|4|||7496|10|||1|
500234066|501840692|500387430|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|376|Red||2009-09-23|2009-10-15|2010-10-26|Child/Family: Moved|Child/Family: Moved||12.4||3|3|1|1|M|White||17||Mother|28226|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||31|28277|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|500234075|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502912141|502932948|500605880|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1534|Red||2012-03-23|2012-04-05|2016-06-17|Volunteer: Moved|Volunteer: Moved||50.4||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Business: Marketing|28203|0|8|Other Church Partner|Faith Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502913549|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|34|2|||7453|7|||1|
500477277|500491044|500134558|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1669|Green|Amachi|2006-10-29|2006-10-29|2011-05-25|Volunteer: Time constraint|Volunteer: Time constraint||54.8||1|1|1|1|F|Black||17||Mother|28213|One Parent: Female|Less than $10,000||||No||Service Organization|General Community||Match Support|F|Black||47|28027|Bachelors Degree|Single|Retail: Sales|28145|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500477524|31|0|2|31|0|2|10|2|500003586||4|1||-2||-2|0|11|||2238|7|||1|500000294
502197477|502422929|500515536|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2062|Green|2010-2012 OJJDP JJI|2011-02-04|2011-02-10|2016-10-03|Volunteer: Moved|Volunteer: Moved||67.7||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28202|Bachelors Degree|Single|Business: Sales|27560|1|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500017732|502197915|31|0|1|1|0|1|10|2|-2||4|1|500005291|-2|500000294, 500004640|-2|0|4|||7464|9|||1|500005291
502206673|502668179|500557233|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1349|Red|Amachi|2011-09-22|2011-10-13|2015-06-23|Child: Lost interest|Child: Lost interest||44.3||1|1|1|1|M|Black||17|Yes|GrandMother|28216|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||47|28216|Bachelors Degree|Married|Business: Engineer|28255|18|0|Self|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500013781|502207102|31|0|1|1|0|1|10|2|500003586||4|3|500000294|-2||-2|0|10|||7464|9|||1|500000294
502551116|500892262|500541956|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|763|Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|2011-06-17|2011-06-30|2013-08-01|Volunteer: Moved|Volunteer: Moved||25.1||1|1|2|2|F|Hispanic||17|Yes|GrandFather|28216|One Parent: Male|$15,000 to $19,999||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black|Other African|36|28105||Single|Consultant|28244|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502551569|3|0|2|31|31|2|10|2|500004772||4|2|500004640, 500005291|-2||-2|0|4|||46|2|||1|500000294, 500004640, 500004901, 500005291
501361902|501307192|500328424|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2974|Green|Amachi|2008-12-19|2009-01-23|NaT||||97.7||1|1|1|1|M|White||17|Yes|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||54|28227|Bachelors Degree|Divorced|Business: Sales|28273|9|5|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|501249611|1|0|1|1|0|1|10|2|500003586||2|1|500000294|-2||-2|0|10|||46|2|||1|500000294
501622502|502162227|500454573|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|606|Green||2010-05-26|2010-06-04|2012-01-31|Volunteer: Time constraint|Volunteer: Time constraint||19.9||2|2|1|1|M|Black||17|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||32|28210|Bachelors Degree|Single|Tech: Engineer||0|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501622822|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501622502|501307502|500356948|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|389|Yellow||2009-04-13|2009-04-24|2010-05-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.8||2|2|1|1|M|Black||17|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||32|28202|||Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501622822|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503476243|503334174|500710120|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|580|Red||2013-09-10|2013-09-20|2015-04-23|Child: Lost interest|Child: Lost interest||19.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||63|28210|Bachelors Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503478109|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7671|13|1561|2|1|
502700505|503029324|500619505|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1723|Green||2012-06-15|2012-06-27|NaT||||56.6||1|1|1|1|M|Black||17|No|Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Black||41|28210|Bachelors Degree|Separated|Arts, Entertainment, Sports|28202|2|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502701350|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
502839800|502847446|500627524|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|717|Green||2012-08-06|2012-08-25|2014-08-12|Volunteer: Moved|Volunteer: Moved||23.6||1|1|1|1|M|Black||17|No|Mother|28213|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||29|28213|Bachelors Degree||Tech: Sales, Mktg|28213|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503677894|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
500545328|501033808|500274449|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3012|Green||2008-06-23|2008-07-02|2016-09-30|Volunteer: Time constraint|Volunteer: Time constraint||99||3|3|1|1|F|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Match Support|F|Black||43|28208|Masters Degree|Single|Business: Sales|28078|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|500545578|7|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500545326|500697845|500134545|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3596|Red||2006-10-29|2006-10-29|2016-09-02|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||118.1|Y|1|1|1|1|M|Multi-Race (None of the above)||17||Mother|28215|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Match Support|M|Black||55|28214||Married|Clergy||12|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|500545578|7|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||2238|7|||1|
502469110|502564995|500535534|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1027|Green|2010-2012 OJJDP JJI|2011-05-09|2011-05-11|2014-03-03|Child/Family: Moved|Child/Family: Moved||33.7||1|1|1|1|M|Black||17|No|Mother|28216|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||35|28269|Associate Degree|Married|Arts, Entertainment, Sports|28262|3|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502469557|31|0|1|31|0|1|10|2|-2||4|1|500005291|-2||-2|0|10|||7496|10|||1|500005291
502997008|502908444|500613594|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|413|Yellow||2012-05-07|2012-05-30|2013-07-17|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||13.6||2|2|1|1|F|Black||17|No|Mother|28226|Two Parent|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||31|28273|Juris Doctorate (JD)|Single|Law: Lawyer||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502998473|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|34|2|||7464|9|||1|
502997008|503517750|500707415|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|427|Green||2013-08-20|2013-09-24|2014-11-25|Child: Lost interest|Child: Lost interest||14||2|2|1|1|F|Black||17|No|Mother|28226|Two Parent|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Education: Teacher Asst/Aid|28214|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|502998473|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|34|2|||7496|10|||1|
502083429|502653045|500590992|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1651|Red||2012-01-11|2012-02-11|2016-08-19|Volunteer: Moved|Volunteer: Moved||54.2||1|1|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Cabarrus County|Match Support|F|Black||29|28027|Bachelors Degree|Single|Education: Teacher||1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500020753|502083853|31|0|2|31|0|2|10|2|-2||4|3|500016374|-2|500016374|-2|7016|11|||7464|9|||1|
501726201|501734664|500371036|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2032|Red|Amachi|2009-06-24|2009-07-08|2015-01-30|Child/Family: Moved|Child/Family: Moved||66.8||1|1|1|1|F|Black||17|Yes|Mother|28212|One Parent: Female|Unknown||||Yes|YeaGod|Faith Organization|General Community|Amachi|Match Support|F|Black||51|28262|PHD|Married|Real Estate: Realtor||0|0|Weeping Willow|Faith Organization|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500008321|501726541|31|0|2|31|0|2|10|2|-2||4|3|500000294|-2||-2|5634|9|||9218|7|||1|500000294
502295599|502306663|500491842|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|421|Red||2010-11-08|2010-11-18|2012-01-13|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.8||1|1|1|1|F|Black||17|No|Mother|28211|One Parent: Female|Unknown||||No|AARTF|BBBS Board/Staff|General Community||Enrollment|F|White||28|28277||Single|Finance: Accountant||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502296031|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|7294|13|||7496|10|||1|
502846423|502877894|500609448|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|297|Yellow||2012-04-11|2012-05-07|2013-02-28|Volunteer: Time constraint|Volunteer: Time constraint||9.8||1|1|1|1|F|Black||17|No|Mother|28215|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Some Other Race||40|28205|Bachelors Degree|Married|Construction|28031|8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502847784|31|0|2|41|0|2|10|2|-2||4|2||-2||-2|0|4|||7496|10|||1|
502269033|502208867|500472485|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|181|Green|Amachi, Project Big, Project Big AND Amachi|2010-09-22|2010-09-29|2011-03-29|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||5.9||1|1|2|2|F|Multi-race (Black & White)||17|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Relative|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community|Project Big AND Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502265485|36|0|2|31|0|2|10|2|500004772||4|1|500004640, 500004901|-2|500004901|-2|0|3|||7464|9|||1|500000294, 500004640, 500004901
503833956|503635291|500761770|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|625|Green||2014-04-30|2014-05-12|2016-01-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.5||1|1|1|1|F|Black||17|No|Mother|28208|Two Parent|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||38|28262|Masters Degree|Single|Finance|28262|0|6|Agency Sponsored|Special Event|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|503835911|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|34|2|||16426|8|||1|
501786018|501559944|500380368|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|367|Green|Amachi|2009-08-21|2009-08-28|2010-08-30|Volunteer: Time constraint|Volunteer: Time constraint||12.1||4|4|1|1|M|Black||17|Yes|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||63|28078||Married|Business: Engineer|28288|0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500010355|501786373|31|0|1|1|0|1|10|2|500003586||4|1||-2||-2|0|10|||7464|9|||1|500000294
501786018|500757564|500468420|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|131|Green|Amachi|2010-09-01|2010-09-22|2011-01-31|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||4.3||4|4|3|3|M|Black||17|Yes|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||51|28216||Married|Craftsman||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|501786373|31|0|1|31|0|1|10|2|500003586||4|1||-2|500000294|-2|0|10|||2238|7|||1|500000294
501786018|503914867|500776457|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|892|Green||2014-09-17|2014-10-06|NaT||||29.3||4|4|1|1|M|Black||17|Yes|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||39|28269|Bachelors Degree|Married|Arts, Entertainment, Sports|28202|15|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|501786373|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501786018|502800403|500589712|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|522|Red|Amachi|2012-01-04|2012-01-23|2013-06-28|Volunteer: Moved|Volunteer: Moved||17.1||4|4|1|1|M|Black||17|Yes|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Asian||28|28203||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501786373|31|0|1|4|0|1|10|2|500003586||4|3||-2||-2|0|10|||7496|10|||1|500000294
501376745|500725077|500350905|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2476|Green||2009-03-19|2009-04-01|2016-01-11|Volunteer: Time constraint|Volunteer: Time constraint||81.3||1|1|3|4|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||34|28269|||Business: Marketing||1|4|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|501377024|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|6854|8|||46|2|||1|
502419933|502442556|500523858|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|211|Green|2010-2012 OJJDP JJI|2011-03-08|2011-03-28|2011-10-25|Volunteer: Time constraint|Volunteer: Time constraint||6.9||2|2|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$40,000 to $44,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||59|28204|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011184|502371107|31|0|1|1|0|1|5|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|500005291
502419933|502669194|500571419|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1002|Yellow||2011-10-27|2011-12-07|2014-09-04|Volunteer: Time constraint|Volunteer: Time constraint||32.9||2|2|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$40,000 to $44,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||58|28031|Bachelors Degree|Living w/ Significant Other|Business: Mgt, Admin||22|0|Big Day|Special Event|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502371107|31|0|1|1|0|1|5|2|-2||4|2|500005291|-2||-2|0|10|||7456|8|||1|
503533026|502485670|500717656|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1244|Green||2013-10-09|2013-10-19|NaT||||40.9||1|1|2|2|F|Black||17|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503534897|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7462|13|1204|3|1|
502067798|502062408|500459576|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2442|Green||2010-06-30|2010-07-09|NaT||||80.2||1|1|1|1|M|Black||17|No|Mother|29732|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||52|28270|Bachelors Degree|Married|Business: Mgt, Admin||4|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502074089|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|
501529921|502554719|500581908|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1169|Green||2011-11-28|2012-01-23|2015-04-06|Volunteer: Time constraint|Volunteer: Time constraint||38.4||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||48|28031|Some College|Divorced|Medical|28031|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501530213|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501529921|501571404|500337752|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|902|Yellow||2009-02-02|2009-02-06|2011-07-28|Volunteer: Time constraint|Volunteer: Time constraint||29.6||2|2|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||39|28209|Masters Degree|Married|Finance: Banking|28202|1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501530213|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501766666|501541222|500386249|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|305|Green|Amachi|2009-09-21|2009-10-02|2010-08-03|Child/Family: Moved|Child/Family: Moved||10||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||31|28211|Bachelors Degree|Single|Unknown|28209|0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500003657|501765484|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
500385150|502330464|500513934|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|318|Yellow|2010-2012 OJJDP JJI|2011-01-27|2011-02-28|2012-01-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.4||3|4|1|1|F|Black||17||Mother|28206|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|RTBM|F|Black||37|28269||Single|Unknown||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500003657|500385400|31|0|2|31|0|2|7|2|-2||4|2|500005291|-2|500000294, 500004640|-2|0|10|||7496|10|||1|500005291
501428903|501441245|500331206|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2226|Green||2009-01-08|2009-01-21|2015-02-25|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||73.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|White||53|15001|Masters Degree|Single|Consultant|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501429188|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502365086|502426330|500509521|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|285|Yellow|Amachi|2011-01-06|2011-01-13|2011-10-25|Child: Lost interest|Child: Lost interest||9.4||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||||Yes|TV|Media|General Community|Amachi|Match Support|M|Black||34|28269|Masters Degree|Married|Tech: Research/Design|19355|1|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502365524|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|56|1|||7446|3|||1|500000294
500947259|501418481|500330761|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|595|Yellow||2009-01-06|2009-01-09|2010-08-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.5||2|2|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$20,000 to $24,999||||No||Self|General Community||RTBM|M|White||52|28205|Masters Degree|Single|Tech: Production Line||0|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|500947529|31|0|1|1|0|1|7|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503209438|503464333|500707202|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|242|Red||2013-08-19|2013-08-31|2014-04-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||8||1|1|1|1|F|Black||17||Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|F|White||29|28205|Masters Degree|Single|Finance: Accountant|28277|1|10|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503211213|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
503014417|503518076|500706096|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1087|Green||2013-08-07|2013-08-26|2016-08-17|Child: Lost interest|Child: Lost interest||35.7||1|1|1|1|F|Black||17|No|Mother|28203|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||29|28110|Masters Degree|Single|Education: Teacher||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503015947|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500293140|500191399|500062178|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1892|Green||2005-12-05|2005-12-05|2011-02-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||62.2||2|2|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||35|28205|Some College|Single|Business: Clerical||0|10|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500191330|31|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|0|10|||46|2|||1|
500293140|503529360|500708612|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|373|Yellow||2013-08-29|2013-09-16|2014-09-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.3||2|2|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||30|28212|Masters Degree|Single|Finance: Accountant|28111|0|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|500191330|31|0|1|1|0|1|10|2|-2||4|2|500005291|-2||-2|0|10|||7464|9|||1|
500914579|501345550|500323102|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2179|Yellow||2008-12-04|2008-12-16|2014-12-04|Child: Severity of challenges|Child: Severity of challenges||71.6||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||Match Support|M|White||32|28277|Bachelors Degree|Single|Tech: Engineer|28117|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500015820|500914849|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502312413|502410938|500509858|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|716|Green|Amachi|2011-01-07|2011-01-18|2013-01-03|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||23.5||1|1|1|1|M|Black||17|Yes|Mother|28211|One Parent: Female|Unknown||||No|Hampton Crest|Service Organization|General Community|Amachi|Match Support|M|White||33|28209|Bachelors Degree|Single|Finance: Economist|60602|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502312845|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|7295|11|||7496|10|||1|500000294
502307585|501519450|500521250|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2187|Green|Amachi, Project Big, Project Big AND Amachi|2011-03-02|2011-03-21|NaT||||71.9||1|1|1|1|F|Black||17|Yes|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||53|28031||Divorced|Medical: Admin|28207|3|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502308017|31|0|2|1|0|2|10|2|500004772||2|1|500000294, 500004640, 500004901|-2||-2|0|4|||7446|3|||1|500000294, 500004640, 500004901
502490193|502547160|500536146|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|596|Red|2010-2012 OJJDP JJI|2011-05-12|2011-05-24|2013-01-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.6||1|1|1|1|M|Black||17|No|Mother|28211|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||40|28277|Masters Degree|Single|Medical: Pharmacist||0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500004169|502490640|31|0|1|1|0|1|5|2|-2||4|3|500005291|-2||-2|6854|8|||7496|10|||1|500005291
501877080|501811850|500440340|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|155|Green||2010-03-10|2010-03-31|2010-09-02|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||5.1||1|1|3|3|M|Black||17|No|Mother|28215|One Parent: Female|Unknown||||Yes|Radio|Media|General Community||Enrollment|M|White||36|28202|||Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|501877453|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|55|1|||7464|9|||1|
502920861|503097126|500639233|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1271|Yellow||2012-09-27|2012-10-29|2016-04-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||41.8||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||34|28203|Juris Doctorate (JD)|Single|Law: Lawyer||2|11|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|502922278|31|0|1|1|0|1|10|2|-2||4|2||-2|500000294|-2|0|10|||7464|9|||1|
502173588|502678947|500677086|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|103|Yellow||2013-01-24|2013-01-31|2013-05-14|Volunteer: Moved|Volunteer: Moved||3.4||2|2|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||||No|A Child's Place|Service Organization|General Community|Amachi|Enrollment|F|White||47|28216|Bachelors Degree|Divorced|Medical: Healthcare Worker|28202|0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502174017|31|0|2|1|0|2|5|2|-2||4|2|500000294|-2||-2|7016|11|||7464|9|||1|
502173588|502085998|500463449|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|734|Yellow|Amachi|2010-07-28|2010-08-27|2012-08-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.1||2|2|1|1|F|Black||17|Yes|Mother|28217|One Parent: Female|Unknown||||No|A Child's Place|Service Organization|General Community|Amachi|Enrollment|F|White||29|28217|Bachelors Degree|Single|Customer Service||5|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502174017|31|0|2|1|0|2|5|2|500003586||4|2|500000294|-2||-2|7016|11|||7496|10|||1|500000294
502570188|502366830|500533448|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2126|Green|Project Big, 2010-2012 OJJDP JJI|2011-04-26|2011-04-30|2017-02-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||69.8||1|1|1|1|F|Black||17|No|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||56|28226|Masters Degree|Married|Medical: Nurse|28217|34|0|Healthy Kids Club|Workplace Partner|Big|General Community|Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020910|502570642|31|0|2|1|0|2|10|2|500004641||4|1|500004640, 500005291|-2|500004640|-2|0|4|||10326|3|||1|500004640, 500005291
502117432|500189709|500438904|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|383|Green||2010-03-03|2010-03-03|2011-03-21|Child/Family: Moved|Child/Family: Moved||12.6||1|1|4|4|F|Black||17|No|Father|28027|One Parent: Male|Unknown||||Yes||BBBS Board/Staff|General Community||Match Support|F|Black||48|28075|Bachelors Degree|Single|Human Services: Non-Profit|28205|0|0|Friendship Missionar|Faith Organization|Big|General Community|Amachi, Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500011639|502117859|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294, 500016374|-2|0|13|||2230|7|||1|
502976039|503150561|500658198|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|104|Red||2012-11-09|2012-11-16|2013-02-28|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||3.4||1|1|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||29|28205|Some College|Single|Medical||2|0|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502977487|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7438|1|||1|
502926909|502880005|500600626|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|503|Red||2012-02-27|2012-03-30|2013-08-15|Volunteer: Moved|Volunteer: Moved||16.5||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community||Match Support|M|White||42|28205|PHD|Divorced|Education: Teacher||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502928325|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|7294|13|||7464|9|||1|
501219652|501216187|500269828|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|646|Green||2008-06-04|2008-06-16|2010-03-24|Volunteer: Time constraint|Volunteer: Time constraint||21.2||1|1|1|1|F|Multi-Race (None of the above)||17|No|Mother|28216|Two Parent|$35,000 to $39,999|||Y|Yes||Therapist/Counselor|General Community||Enrollment|F|White||39|28202|Masters Degree|Married|Business: Marketing|28203|0|1|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|501219928|7|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|5|||46|2|||1|
501015965|500189376|500447721|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1259|Yellow|Amachi|2010-04-16|2010-04-29|2013-10-09|Child: Lost interest|Child: Lost interest||41.4||2|2|2|2|F|Black||17|Yes|Mother|28208|One Parent: Female|Less than $10,000||||Yes||Self|General Community|Amachi|Match Support|F|Black||60|28269|Bachelors Degree|Married|Human Services: Non-Profit||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|501016235|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
501015965|501012047|500238959|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|462|Green|Amachi|2008-01-22|2008-02-12|2009-05-19|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||15.2||2|2|1|1|F|Black||17|Yes|Mother|28208|One Parent: Female|Less than $10,000||||Yes||Self|General Community|Amachi|Match Support|F|White||36|28270|Masters Degree|Married|Finance: Auditor||4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501016235|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||46|2|||1|500000294
501318837|501357948|500304715|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|595|Green||2008-10-24|2008-11-04|2010-06-22|Volunteer: Moved|Volunteer: Moved||19.5||2|2|1|1|M|Black||17|No|Mother|28205|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||39|28202|Juris Doctorate (JD)|Single|Law: Lawyer|10017|0|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501319115|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|6854|8|||7464|9|||1|
501318837|502170420|500459741|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|938|Red||2010-07-01|2010-08-04|2013-02-27|Volunteer: Time constraint|Volunteer: Time constraint||30.8||2|2|1|1|M|Black||17|No|Mother|28205|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Retail: Sales||0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|501319115|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|6854|8|||7496|10|||1|
501528770|501801101|500378639|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|355|Yellow||2009-08-13|2009-08-21|2010-08-11|Volunteer: Time constraint|Volunteer: Time constraint||11.7||1|1|1|1|M|Black||17|Yes|Mother|28214|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|White||34|28209|||Business: Sales|32246|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|501529062|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
500418050|500417272|500093386|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2392|Green|Amachi|2006-05-12|2006-05-12|2012-11-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||78.6||1|1|1|1|M|Black||17|Yes|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||34|28273|High School Graduate|Single|Transport: Driver|28216|0|10|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500188055|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
502015842|502160380|500461467|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|462|Green|Amachi|2010-07-19|2010-07-21|2011-10-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||15.2||1|1|1|1|M|Black||17|Yes|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|RTBM|M|White||35|28211|Bachelors Degree|Single|Finance||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|502016241|31|0|1|1|0|1|7|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501340097|501353925|500284012|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|468|Green|Amachi|2008-08-27|2008-09-18|2009-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||15.4||2|2|1|1|M|Multi-race (Black & Hispanic)||17|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||39|28205|Bachelors Degree|Single|Tech: Engineer|28205|0|8|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501340376|38|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||46|2|||1|500000294
501340097|501934966|500440292|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2372|Red|Amachi|2010-03-10|2010-03-23|2016-09-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||77.9||2|2|1|1|M|Multi-race (Black & Hispanic)||17|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Hispanic||28|28277|Some College|Single|Student: College|28223|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|501340376|38|0|1|3|0|1|10|2|500003586||4|3|500000294|-2||-2|0|10|||7464|9|||1|500000294
502710796|502926804|500608316|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1798|Green|Project Big|2012-04-05|2012-04-13|NaT||||59.1||1|1|1|1|M|Black||17|No|GrandMother|28208|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community|Project Big|Match Support|M|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502711683|31|0|1|1|0|1|10|2|500004641||2|1|500004640|-2||-2|6854|8|||7464|9|||1|500004640
500764138|500696779|500154924|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2206|Green|Amachi|2007-01-26|2007-02-07|2013-02-21|Volunteer: Time constraint|Volunteer: Time constraint||72.5||2|2|1|1|M|Black||17|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community|Amachi|Match Support|M|Black||33|28214||Single|Tech: Research/Design||1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500764404|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500764138|503707921|500758491|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|662|Red||2014-04-07|2014-05-31|2016-03-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.7||2|2|1|1|M|Black||17|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community|Amachi|Match Support|M|White||29|28210|Bachelors Degree|Single|Finance||2|4|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|500764404|31|0|1|1|0|1|10|2|-2||4|3|500000294|-2|500000294|-2|0|10|||7464|9|||1|
502137968|502417993|500521032|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|672|Red|2010-2012 OJJDP JJI|2011-03-01|2011-03-08|2013-01-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||22.1||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||41|28078|Bachelors Degree|Married|Govt|28262|7|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502138397|31|0|1|1|0|1|10|2|-2||4|3|500005291|-2|500000294, 500004640|-2|34|2|||7464|9|||1|500005291
502732602|502766077|500588408|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|510|Yellow||2011-12-21|2012-01-25|2013-06-18|Volunteer: Moved|Volunteer: Moved||16.8||1|1|1|1|F|Black||17|No|Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|White||29|28203|Masters Degree|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502733499|31|0|2|1|0|2|10|2|-2||4|2|500005291|-2||-2|0|5|||7464|9|||1|
500426096|500433762|500101957|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1444|Red||2006-06-21|2006-06-26|2010-06-09|Volunteer: Time constraint|Volunteer: Time constraint||47.4||1|1|1|1|M|Black||17||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||35|28262|Bachelors Degree|Single|Tech: Support, Writing|28211|0|8|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500426342|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502259046|502502361|500537239|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|845|Yellow||2011-05-20|2011-05-25|2013-09-16|Volunteer: Time constraint|Volunteer: Time constraint||27.8||1|1|1|1|F|White||17|No|Mother|28025|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Enrollment|F|White||64|28083|High School Graduate|Married|Finance: Banking||0|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502259478|1|0|2|1|0|2|5|2|||4|2||-2||-2|6854|8|||7464|9|||1|
502097843|502643791|500550390|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1809|Green|2010-2012 OJJDP JJI|2011-08-16|2011-08-29|2016-08-11|Child: Lost interest|Child: Lost interest||59.4||1|1|2|2|M|Black||17|No|Mother|28078|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Hispanic||35|28078|Bachelors Degree|Single|Business: Mgt, Admin|28031|13|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|502098263|31|0|1|3|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|500005291
502494753|502481799|500529173|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|922|Yellow|Amachi, Project Big, Project Big AND Amachi|2011-04-04|2011-04-14|2013-10-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||30.3||1|1|1|1|F|Black||17|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28212|Masters Degree|Single|Business|28105|5|8|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502495202|31|0|2|31|0|2|10|2|500004772||4|2|500000294, 500004640, 500004901|-2||-2|0|4|||7438|1|||1|500000294, 500004640, 500004901
502802219|503060158|500623104|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|577|Green||2012-07-06|2012-07-30|2014-02-27|Volunteer: Time constraint|Volunteer: Time constraint||19||1|1|1|1|M|White||17|No|Mother|28209|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|White||35|28212|Some College|Single|Tech: Computer/Programmer|28212|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502803493|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500340183|500785600|500163811|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|973|Green||2007-02-27|2007-03-13|2009-11-10|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||32||3|3|1|1|M|Black||17|No|Relative: Other|28208|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||39|28209|Associate Degree|Married|Business: Sales|28079|2|9|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500340317|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500340183|501933993|500419988|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1351|Yellow||2009-12-09|2009-12-18|2013-08-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||44.4||3|3|1|1|M|Black||17|No|Relative: Other|28208|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction||0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|500340317|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
500340183|503868914|500766977|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|996|Green||2014-06-18|2014-06-24|NaT||||32.7||3|3|1|1|M|Black||17|No|Relative: Other|28208|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||29|28205||Single|Consultant|2210|2|10|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|500340317|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1|
503443162|500234684|500705816|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|540|Yellow||2013-08-05|2013-08-20|2015-02-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.7||1|1|2|2|M|Black||17|No|Mother|28262|One Parent: Female|$25,000 to $29,999||||Yes||Relative|General Community||Match Support|M|Black||34|28213|Bachelors Degree|Single|Finance: Banking|28202|0|2|Recruitment Event|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503445028|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|3|||7458|9|||1|
502828131|502881454|500607446|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1065|Red||2012-04-01|2012-04-30|2015-03-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||35||1|1|1|1|F|Multi-Race (None of the above)||17|No|Father|28214|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|White||33|28216|Bachelors Degree|Single|Business: Sales|28270|2|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502829415|7|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500829028|501978180|500498594|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2298|Green||2010-11-22|2010-11-30|NaT||||75.5||3|3|2|2|F|Black||17|No|Mother|28209|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|F|White||39|28210|Masters Degree|Single|Education|28212|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020910|502254499|31|0|2|1|0|2|10|2|-2||2|1||-2|500000294, 500004640|-2|0|10|||7464|9|||1|
500829028|502192090|500467543|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|60|Green||2010-08-26|2010-09-03|2010-11-02|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||2||3|3|2|2|F|Black||17|No|Mother|28209|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|F|White||32|28134|Bachelors Degree|Single|Finance: Banking|28288|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|502254499|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502868969|503574667|500736904|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1184|Green||2013-12-05|2013-12-18|NaT||||38.9||1|1|1|1|F|Black||17|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||26|11237||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020753|502870370|31|0|2|1|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||46|2|||1|
502469903|502868874|500594396|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1849|Green||2012-01-27|2012-02-22|NaT||||60.7||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|$15,000 to $19,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||34|28269|Bachelors Degree|Single|Business: Human Resources|28025|2|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502470350|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|5|||4748|14|1360|3|1|
503580303|503487684|500715761|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|246|Green||2013-10-03|2013-10-15|2014-06-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.1||1|1|1|1|M|Black||17|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|M|White||42|28212|Bachelors Degree|Single|Business: Engineer||0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|503582180|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500781019|500713642|500167249|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1317|Red||2007-03-16|2007-03-23|2010-10-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||43.3||1|1|1|1|M|Black||17|No|Mother|28105|One Parent: Female|$30,000 to $34,999|||Y|No|BBBS National Site|Web Link|General Community||Enrollment|M|White||40|28270||Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500781287|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
503813942|503873603|500773055|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|913|Green||2014-08-21|2014-08-30|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||30||1|1|1|1|M|Black||17|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|M|Black||38|28269||Single|Unemployed||0|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503815919|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|3|||17101|1|||1|
500433644|501882367|500430294|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|664|Red||2010-01-27|2010-02-04|2011-11-30|Volunteer: Time constraint|Volunteer: Time constraint||21.8||2|2|1|1|M|Black||17||Mother|28269|One Parent: Female|Unknown||||No||Relative|General Community||Enrollment|M|Black||60|28078|Bachelors Degree|Married|Tech: Computer/Programmer|28202|25|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|500433894|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|0|3|||7464|9|||1|
502602958|502578040|500552390|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1992|Green|Project Big, 2010-2012 OJJDP JJI|2011-08-29|2011-09-11|2017-02-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||65.4||1|1|1|1|M|Black||17|No|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||52|28207|Masters Degree|Married|Business|28202|0|7|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|501480402|31|0|1|1|0|1|10|2|500004641||4|1|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291
501195410|501277677|500278978|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3135|Green||2008-07-23|2008-08-15|NaT||||103||1|1|1|1|M|Black||17|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Asian||35|28210|Bachelors Degree|Married|Business: Sales|28217|5|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501195684|31|0|1|4|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503873575|504004351|500796129|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|332|Green||2014-11-17|2014-11-24|2015-10-22|Child/Family: Moved|Child/Family: Moved||10.9||1|1|1|1|F|Black||17|No|Mother|28269|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||39|28078|Bachelors Degree|Single|Business: Sales|28117|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503875571|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
503923102|503996589|500781196|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|885|Green||2014-10-07|2014-10-13|NaT||||29.1||1|1|1|1|M|Black||17|No|Mother|28213|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|Black||48|28262||Single|Retired||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503925109|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1|
503796616|503828896|500772098|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|421|Green||2014-08-12|2014-08-25|2015-10-20|Volunteer: Time constraint|Volunteer: Time constraint||13.8||1|1|1|1|F|Black||17|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||30|28273|Bachelors Degree|Single|Business: Human Resources|28203|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503798593|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
502761850|503632186|500738602|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1146|Green|Cabarrus County|2013-12-12|2014-01-25|NaT||||37.7||2|2|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||41|28027|Bachelors Degree|Married|Human Services|28025|0|9|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502762654|31|0|2|31|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
502761850|502925181|500623917|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|369|Yellow||2012-07-12|2012-07-18|2013-07-22|Volunteer: Moved|Volunteer: Moved||12.1||2|2|1|1|F|Black||17|No|Mother|28083|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||26|28212|Some College|Single|Military||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500012459|502762654|31|0|2|31|0|2|10|2|-2||4|2|500016374|-2||-2|0|10|||7496|10|||1|
501330620|501236896|500290146|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|899|Green||2008-09-22|2008-09-29|2011-03-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29.5||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||43|28078|Masters Degree|Married|Self-Employed, Entrepreneur||1|6|Self|Self|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500011184|501330898|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503587930|500942257|500742670|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|374|Yellow||2014-01-14|2014-01-27|2015-02-05|Volunteer: Time constraint|Volunteer: Time constraint||12.3||1|1|3|3|M|Black||16|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||26|28203|Bachelors Degree|Single|Finance: Banking|28213|0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503589807|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501735420|500956022|500428818|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2025|Green||2010-01-21|2010-01-26|2015-08-13|Child: Lost interest|Child: Lost interest||66.5||2|2|2|2|F|Black||16||GrandMother|28215|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||41|28277|Bachelors Degree|Single|Business: Mgt, Admin||9|0|General|Other Big|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500017732|501735760|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|6854|8|||6450|12|||1|
501735420|501596594|500374040|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|92|Yellow||2009-07-15|2009-08-13|2009-11-13|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3||2|2|1|1|F|Black||16||GrandMother|28215|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||37|28227|||Retail: Sales|28213|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501735760|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1|
500713817|501834795|500396466|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2694|Green||2009-10-19|2009-10-30|NaT||||88.5||2|2|1|1|M|Black||16||Mother|28216|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28078|||Medical: Pharmacist|28210|10|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|500714084|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1|
501234606|501233675|500287478|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3103|Green||2008-09-11|2008-09-16|NaT||||101.9||1|1|1|1|F|Black||16|No|Mother|28216|Grandparents|Unknown||||No|TV|Media|General Community||Match Support|F|Black||42|28212|Bachelors Degree|Single|Unknown|28202|8|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501234882|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|56|1|||7464|9|||1|
500872671|501202985|500262133|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|392|Green|Amachi|2008-04-22|2008-04-22|2009-05-19|Volunteer: Moved|Volunteer: Moved||12.9||1|1|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community|Amachi|Match Support|M|White||33|28202|Bachelors Degree|Single|Construction|28217|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500872940|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||46|2|||1|500000294
502221847|502103416|500459547|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|407|Green|Amachi|2010-06-30|2010-07-12|2011-08-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.4||2|2|1|1|F|Black||16|Yes|GrandMother|28213|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28212|Bachelors Degree|Single|Law|29715|2|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502222278|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7496|10|||1|500000294
502221847|502654877|500556560|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1997|Green|Amachi|2011-09-21|2011-09-27|NaT||||65.6||2|2|1|1|F|Black||16|Yes|GrandMother|28213|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||24|28027|Some College|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502222278|31|0|2|31|0|2|10|2|500003586||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
500896024|500865849|500341304|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|468|Green|Amachi|2009-02-16|2009-02-20|2010-06-03|Volunteer: Time constraint|Volunteer: Time constraint||15.4||1|1|2|2|M|Black||16|Yes|Mother|28027|One Parent: Female|Unknown||||No||Faith Organization|General Community|Amachi|Match Support|M|Black||55|28083||Single|Govt: Mgmt/Admin||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002335|500896288|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
502294498|502639594|500546657|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|735|Red|2010-2012 OJJDP JJI|2011-07-19|2011-08-11|2013-08-15|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.1||1|1|1|1|M|Some Other Race||16|No|Mother|28105|One Parent: Female|Unknown||||No||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Enrollment|M|Black||47|28227|Some College|Single|Finance: Banking|28262|22|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502294930|41|0|1|31|0|1|5|2|-2||4|3|500005291|-2||-2|0|5|||7464|9|||1|500005291
501588821|501359582|500429105|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|833|Green||2010-01-22|2010-02-10|2012-05-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27.4||1|1|2|2|F|Black||16||Mother|28208|Two Mothers|Unknown||||Yes||Self|General Community||Match Support|F|Black||34|28273|Masters Degree|Living w/ Significant Other|Consultant|28273|1|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501589141|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
502551045|502864071|500597976|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|743|Yellow||2012-02-13|2012-02-22|2014-03-06|Volunteer: Health|Volunteer: Health||24.4||2|2|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||54|28031|Bachelors Degree|Married|Business: Mgt, Admin|28262|8|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502551498|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|4|||7464|9|||1|
502551045|503859553|500772207|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|244|Red||2014-08-13|2014-08-29|2015-04-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||8||2|2|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||34|28269|Masters Degree|Single|Medical|28025|1|7|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|502551498|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||17159|12|||1|
500185624|500923420|500182113|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2070|Yellow|Amachi|2007-06-25|2007-06-28|2013-02-26|Child/Family: Moved|Child/Family: Moved||68||1|1|1|1|M|Black||16|Yes|Mother|28213|Other/Unknown|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||61|28205||Married|Tech: Management||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500012459|500187258|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|5635|9|||2238|7|||1|500000294
501955313|500915390|500427542|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|564|Green||2010-01-19|2010-01-29|2011-08-16|Volunteer: Moved|Volunteer: Moved||18.5||2|2|1|1|F|Black||16||Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28270||Single|Business: Clerical||10|0|TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|501955711|31|0|2|1|0|2|10|2|-2||4|1|500005291|-2||-2|0|10|||130|1|||1|
501955313|502609427|500558508|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|402|Red|2010-2012 OJJDP JJI|2011-09-27|2011-10-31|2012-12-06|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||13.2||2|2|1|1|F|Black||16||Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||26|28262|Some College|Single|Business: Clerical||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500015820|501955711|31|0|2|31|0|2|10|2|-2||4|3|500005291|-2|500004640|-2|0|10|||7496|10|||1|500005291
500870686|501101027|500248098|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1207|Red||2008-02-26|2008-02-26|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||39.7||1|1|1|1|M|Black||16|No|Mother|28078|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|White||38|28031|Bachelors Degree|Single|Business: Mgt, Admin||0|7|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500870955|31|0|1|1|0|1|10|2|||4|3||-2||-2|0|10|||46|2|||1|
501831955|501972975|500418296|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|320|Green||2009-12-04|2009-12-11|2010-10-27|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||10.5||1|1|1|1|M|White||16||Mother|28027|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||37|28025|High School Graduate|Divorced|Unknown||1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501832323|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502211307|502371462|500512414|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1176|Yellow|Amachi|2011-01-21|2011-02-03|2014-04-24|Volunteer: Time constraint|Volunteer: Time constraint||38.6||1|1|1|1|M|Black||16|Yes|Mother|28278|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||51|28214|Bachelors Degree|Single|Business: Sales|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|502211737|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2|500000294|-2|7016|11|||7496|10|||1|500000294
502540400|502540283|500533007|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|276|Red|Project Big, 2010-2012 OJJDP JJI|2011-04-23|2011-04-25|2012-01-26|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||9.1||1|1|1|1|M|Black||16|No|GrandMother|28208|Grandparents|Unknown|||Y|Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||68|28025||Widowed|Education|28212|5|0|A Child's Place|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502540853|31|0|1|1|0|1|10|2|500004641||4|3|500004640, 500005291|-2||-2|7016|11|||11610|6|1210|1|1|500004640, 500005291
500900251|501174923|500269471|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|216|Green|Amachi|2008-06-02|2008-06-10|2009-01-12|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.1||1|1|2|2|M|Black||16|Yes|Mother|28078|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|M|Black||70|28078|Bachelors Degree|Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500900521|31|0|1|31|0|1|5|2|500003586||4|1|500000294|-2||-2|0|10|||46|2|||1|500000294
501833031|502427342|500518294|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1710|Red|2010-2012 OJJDP JJI|2011-02-17|2011-02-28|2015-11-04|Volunteer: Moved|Volunteer: Moved||56.2||1|1|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28205|Masters Degree|Single|Medical: Doctor, Provider|28277|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|501833394|31|0|2|1|0|2|10|2|-2||4|3|500005291|-2||-2|0|10|||7464|9|||1|500005291
502580335|502677590|500571804|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1933|Green||2011-10-28|2011-11-30|NaT||||63.5||1|1|1|1|F|Black||16||GrandMother|28269|Grandparents|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28269|Masters Degree|Single|Finance: Banking|28255|15|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502580838|31|0|2|31|0|2|10|2|-2||2|1|500005291|-2||-2|0|10|||7464|9|||1|
501347793|500928548|500289533|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|711|Green||2008-09-19|2008-11-10|2010-10-22|Volunteer: Time constraint|Volunteer: Time constraint||23.4||1|1|1|1|M|Black||16|No|Mother|28202|One Parent: Female|Unknown||||Yes||Neighbor/Friend|General Community||Match Support|M|White||33|28211|Bachelors Degree|Single|Business: Marketing|28202|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501348072|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|8|||46|2|||1|
502615628|502635965|500551985|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|110|Green||2011-08-25|2011-09-09|2011-12-28|Volunteer: Time constraint|Volunteer: Time constraint||3.6||1|1|2|2|M|Black||16|No|Mother|28215|One Parent: Female|$10,000 to $14,999||||Yes||Therapist/Counselor|General Community||RTBM|M|Black||27|28262|Associate Degree|Divorced|Medical: Nurse|28203|1|0|Self|Self|Big|General Site||Match Support|0|1|1|0|277|60|598|500000170|500001281|502616240|31|0|1|31|0|1|7|2|-2||4|1||-2||-1|0|5|||7464|9|||1|
503524036|503913408|500774440|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|893|Green|PERL 2014-2016|2014-09-04|2014-09-19|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||29.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Black||39|28262|Bachelors Degree|Single|Finance|28262|3|2|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|503525911|31|0|1|31|0|1|10|2|-2||4|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681
502290880|502261364|500471473|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1258|Green|Project Big|2010-09-20|2010-10-20|2014-03-31|Child/Family: Time constraints|Child/Family: Time constraints||41.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|M|White||35|28202|Bachelors Degree|Single|Real Estate: Realtor|28208|2|10|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502291312|31|0|1|1|0|1|10|2|500004641||4|1|500004640|-2||-2|0|4|||7496|10|||1|500004640
503767186|503788125|500766047|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|997|Green||2014-06-10|2014-06-23|NaT||||32.8||1|1|1|1|F|Black||16|No|Mother|28227|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||30|28205|Bachelors Degree|Single|Business|28262|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503769162|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
504085882|503977000|500794719|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|830|Red|PERL 2014-2016|2014-11-12|2014-11-21|2017-02-28|Child/Family: Time constraints|Child/Family: Time constraints||27.3||1|1|1|1|F|Black||16|No|GrandMother|28269|One Parent: Female|Unknown|||Y|Yes||Foster Home|General Community|PERL 2014-2016|Match Support|F|Black||24|28217|Bachelors Degree|Single|Finance||0|2|AA Task Force|BBBS Board/Staff|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503144847|31|0|2|31|0|2|10|2|-2||4|3|500014681|-2|500014681|-2|0|7|||9229|13|||1|500014681
502256918|502143354|500501039|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|870|Red||2010-12-01|2010-12-07|2013-04-25|Child/Family: Moved|Child/Family: Moved||28.6||1|1|1|1|M|Hispanic||16|No|Mother|28212|One Parent: Female|Unknown||||No|Spanish Print|Media|General Community||Match Support|M|White||38|28209|Juris Doctorate (JD)|Single|Law||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502257350|3|0|1|1|0|1|10|2|-2||4|3||-2||-2|7063|1|||7464|9|||1|
501628854|503374490|500682899|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|605|Yellow||2013-02-19|2013-03-05|2014-10-31|Volunteer: Moved|Volunteer: Moved||19.9||3|3|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||42|28205|Associate Degree|Single|Transport: Flight Attendant||8|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500015820|501629177|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1|
501628854|501595632|500368527|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|534|Green|Amachi|2009-06-11|2009-06-15|2010-12-01|Volunteer: Time constraint|Volunteer: Time constraint||17.5||3|3|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||34|28217|||Business: Engineer|28134|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|501629177|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501628854|502091655|500521158|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|609|Green||2011-03-02|2011-03-31|2012-11-29|Volunteer: Moved|Volunteer: Moved||20||3|3|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||33|28277|Bachelors Degree|Married|Finance|28209|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501629177|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7496|10|||1|
501096791|503803014|500768008|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|974|Green||2014-06-27|2014-07-16|NaT||||32||3|3|1|1|F|Black||16|Yes|Mother|28206|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|Black||28|28223|Masters Degree|Single|Student: College|28223|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|501097065|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|4|||46|2|||1|
502307352|502217265|500485187|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|248|Green|Amachi, Project Big, Project Big AND Amachi|2010-10-25|2010-11-22|2011-07-28|Volunteer: Moved|Volunteer: Moved||8.1||2|2|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community|Project Big AND Amachi|Match Support|F|Black||34|28208|PHD|Single|Medical: Doctor, Provider||1|0|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011184|502307784|31|0|2|31|0|2|10|2|500004772||4|1|500004901|-2|500004640|-2|0|4|||7464|9|||1|500000294, 500004640, 500004901
502307352|502636073|500552236|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|547|Red|Amachi, Project Big AND Amachi|2011-08-29|2011-08-31|2013-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18||2|2|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community|Project Big AND Amachi|Match Support|F|Black||33|28217|PHD|Single|Medical: Doctor, Provider||0|0|Recruitment Event|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502307784|31|0|2|31|0|2|10|2|500004772||4|3|500004901|-2||-2|0|4|||7460|12|||1|500000294, 500004901
502787524|502272989|500587325|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|947|Red||2011-12-15|2012-01-25|2014-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||31.1||1|1|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Asian||29|28202||Single|Tech: Computer/Programmer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502788707|38|0|2|4|0|2|10|2|-2||4|3||-2|500004640|-2|0|10|||7496|10|||1|
502555551|503207140|500674218|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1296|Green||2013-01-10|2013-01-30|2016-08-18|Child/Family: Moved|Child/Family: Moved||42.6||2|2|1|1|M|Black||16|No|Aunt|28213|One Parent: Female|$40,000 to $44,999||||Yes||School|General Community|Project Big|Match Support|M|White||33|28209|Associate Degree|Married|Business: Mgt, Admin||0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|502556004|31|0|1|1|0|1|10|2|-2||4|1|500004640|-2||-2|0|4|||7464|9|||1|
502555551|502629285|500546255|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|371|Red|Project Big|2011-07-14|2011-07-21|2012-07-26|Volunteer: Moved|Volunteer: Moved||12.2||2|2|1|1|M|Black||16|No|Aunt|28213|One Parent: Female|$40,000 to $44,999||||Yes||School|General Community|Project Big|Match Support|M|White||27|28205|Associate Degree|Single|Service: Restaurant||0|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502556004|31|0|1|1|0|1|10|2|-2||4|3|500004640|-2||-2|0|4|||7464|9|||1|500004640
502268597|502097001|500466598|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|419|Green||2010-08-23|2010-09-01|2011-10-25|Child/Family: Moved|Child/Family: Moved||13.8||1|1|1|1|F|Black||16|No|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||37|28211|Bachelors Degree|Single|Arts, Entertainment, Sports||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502269029|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500824037|500789337|500165956|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3654|Green||2007-03-08|2007-03-15|NaT||||120||1|1|1|1|F|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||Match Support|F|White||34|28210|Bachelors Degree|Single|Education: Teacher|28226|0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|500824306|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502568883|502501016|500533467|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|384|Red|Project Big, 2010-2012 OJJDP JJI|2011-04-26|2011-05-13|2012-05-31|Volunteer: Time constraint|Volunteer: Time constraint||12.6||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|$15,000 to $19,999||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||30|28262|Masters Degree|Single|Customer Service|28262|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502569337|31|0|2|31|0|2|5|2|500004641||4|3|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291
502581328|503144090|500681651|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|879|Yellow||2013-02-13|2013-02-28|2015-07-27|Child: Lost interest|Child: Lost interest||28.9||1|1|1|1|F|Black||16|No|GrandMother|28212|One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||46|28262|PHD|Single|Education: College Professor|28223|5|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|502581832|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1|
502063945|502295138|500478943|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2115|Yellow||2010-10-11|2010-10-21|2016-08-05|Volunteer: Time constraint|Volunteer: Time constraint||69.5||1|1|1|1|M|White||16|No|Mother|28213|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community||Match Support|M|White||37|28205||Married|Real Estate: Realtor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502064367|1|0|1|1|0|1|10|2|500004641||4|2||-2||-2|0|5|||7496|10|||1|
501750507|501582859|500374145|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|560|Green||2009-07-15|2009-07-29|2011-02-09|Volunteer: Time constraint|Volunteer: Time constraint||18.4||2|2|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||42|28262||Single|Finance: Banking|28255|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501750847|31|0|2|1|0|2|5|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|
501750507|502275127|500557811|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|622|Red||2011-09-26|2011-09-30|2013-06-13|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||20.4||2|2|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|Black||35|28212|Masters Degree|Single|Human Services: Social Worker|28204|2|5|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500015820|501750847|31|0|2|31|0|2|5|2|-2||4|3|500005291|-2|500004640|-2|0|10|||7464|9|||1|
502596391|502485670|500540403|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|800|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-06-08|2011-06-12|2013-08-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||26.3||1|1|2|2|F|Black||16|No|Mother|28208|Two Mothers|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28217|Bachelors Degree|Single|Finance||0|1|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502596909|31|0|2|31|0|2|10|2|500004641||4|2|500004640, 500005291|-2||-2|0|4|||7462|13|1204|3|1|500004640, 500005291
502338222|502255795|500483087|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|700|Red|Project Big|2010-10-20|2010-10-27|2012-09-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||23||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Enrollment|F|Black||43|28105|Some College|Single|Business: Mgt, Admin|28226|11|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502338658|31|0|2|31|0|2|5|2|500004641||4|3|500004640|-2|500004640|-2|0|4|||7496|10|||1|500004640
502338225|502312449|500483095|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2038|Yellow|Project Big|2010-10-20|2010-10-27|2016-05-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||67||1|1|1|1|F|Black||16||Mother|28212|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|F|White||33|28227|Bachelors Degree|Single|Unknown||9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|0|1|277|60|598|500000170|500008321|502338658|31|0|2|1|0|2|10|2|500004641||4|2|500004640|-2|500004640|-2|0|4|||7496|10|||1|500004640
500930012|501207610|500269442|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|250|Red||2008-06-02|2008-06-06|2009-02-11|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||8.2||1|1|1|1|F|Black||16|No|Aunt|28208|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community||Match Support|F|White||40|28205|Bachelors Degree|Single|Business: Mgt, Admin|28202|0|10|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|500930282|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
502307478|502035292|500503967|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|486|Red|Project Big|2010-12-09|2010-12-31|2012-04-30|Volunteer: Moved|Volunteer: Moved||16||1|1|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Enrollment|M|Black||40|28215|Some College|Married|Transport: Driver||3|0|Michael Baisden|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013709|502307910|31|0|1|31|0|1|5|2|||4|3|500004640|-2||-2|0|4|||11146|1|||1|500004640
500186245|502989318|500614903|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1757|Green|Amachi|2012-05-15|2012-05-24|NaT||||57.7||2|3|1|1|M|Black||16|Yes|Mother|28216|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Match Support|M|White||34|28203|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|500187840|31|0|1|1|0|1|10|2|500003586||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501524313|501508941|500381084|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|213|Green||2009-08-26|2009-09-22|2010-04-23|Child/Family: Moved|Child/Family: Moved||7||2|2|2|2|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||36|28278|Bachelors Degree|Single|Retail: Sales|30071|5|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500009242|501524605|31|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|
501524313|502615076|500547406|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|993|Green|2010-2012 OJJDP JJI|2011-07-25|2011-08-02|2014-04-21|Volunteer: Moved|Volunteer: Moved||32.6||2|2|1|1|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28208|Bachelors Degree|Single|Finance: Economist|28202|5|6|Recruitment Event|BBBS Board/Staff|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500017777|501524605|31|0|1|1|0|1|10|2|-2||4|1|500005291|-2|500005291|-2|0|10|||7462|13|||1|500005291
500583932|500713684|500149413|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|707|Green||2006-12-19|2007-01-31|2009-01-07|Volunteer: Moved Vol: Other Reason|Volunteer: Moved|Vol: Other Reason|23.2||1|1|1|1|M|Black||16||Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|M|White||41|28217||Single|Finance: Economist||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500584184|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502505252|503429848|500699545|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|148|Red||2013-06-05|2013-06-26|2013-11-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||4.9||2|2|1|1|F|Black||16|No|Mother|28209|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||56|28217|Some College|Single|Finance||9|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502505701|31|0|2|31|0|2|10|2|-2||4|3|500005291|-2||-2|0|10|||7464|9|||1|
502505252|502350629|500525884|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|556|Yellow|2010-2012 OJJDP JJI|2011-03-16|2011-03-21|2012-09-27|Volunteer: Moved|Volunteer: Moved||18.3||2|2|1|1|F|Black||16|No|Mother|28209|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||30|28202|Bachelors Degree|Single|Finance: Accountant|28203|2|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500011746|502505701|31|0|2|1|0|2|10|2|-2||4|2|500005291|-2|500005291|-2|0|10|||7464|9|||1|500005291
502168082|502240884|500505682|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|386|Red|2010-2012 OJJDP JJI|2010-12-14|2011-01-05|2012-01-26|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.7||1|1|1|1|F|Black||16|No|GrandMother|28208|Grandparents|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|F|White||43|28210|Bachelors Degree|Single|Business: Sales|6830|3|0|Self|Self|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500013709|502168511|31|0|2|1|0|2|10|2|-2||4|3|500005291|-2||-2|34|2|||7464|9|||1|500005291
502307545|502782829|500582593|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|638|Green|Project Big|2011-11-29|2011-11-30|2013-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||21||2|2|1|1|F|Hispanic||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|F|Hispanic||38|28209|Bachelors Degree||Business||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502307977|3|0|2|3|0|2|10|2|500004641||4|1|500004640|-2||-2|0|4|||7464|9|||1|500004640
502307545|502172480|500483395|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|363|Yellow|Project Big|2010-10-20|2010-10-27|2011-10-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.9||2|2|1|1|F|Hispanic||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|F|Hispanic||33|28216|Some College|Widowed|Retail: Mgt||5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011184|502307977|3|0|2|3|0|2|10|2|500004641||4|2|500004640|-2|500004640|-2|0|4|||7496|10|||1|500004640
501227649|503316978|500677437|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1491|Green|Cabarrus County|2013-01-25|2013-02-14|NaT||||49||2|2|1|1|M|White||16|Yes|GrandMother|28083|Grandparents|Unknown|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||51|28117|Masters Degree|Divorced|Consultant|28117|12|11|Local Print|Media|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|501227925|1|0|1|1|0|1|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|10|||7439|1|||1|500016374
501227649|501485340|500340341|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|999|Green|Amachi|2009-02-11|2009-02-12|2011-11-08|Volunteer: Time constraint|Volunteer: Time constraint||32.8||2|2|1|1|M|White||16|Yes|GrandMother|28083|Grandparents|Unknown|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||37|28083|Masters Degree|Single|Business: Sales||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501227925|1|0|1|1|0|1|10|2|500003586||4|1|500000294, 500016374|-2||-2|0|10|||7464|9|||1|500000294
500761491|502189613|500465204|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|938|Green||2010-08-10|2010-08-27|2013-03-22|Volunteer: Time constraint|Volunteer: Time constraint||30.8||3|3|1|1|F|Black||16||Aunt|28213|One Parent: Female|$40,000 to $44,999|||Y|No||Self|General Community||Enrollment|F|Black||61|28269|Bachelors Degree|Divorced|Education: Teacher|28215|1|1|LPL Financial|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|500761759|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||11247|3|||1|
500761491|500188903|500268793|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|713|Green||2008-05-28|2008-06-04|2010-05-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||23.4||3|3|2|2|F|Black||16||Aunt|28213|One Parent: Female|$40,000 to $44,999|||Y|No||Self|General Community||Enrollment|F|Black||34|28215|Bachelors Degree|Single|Finance: Banking||0|1|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500761759|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500783100|500777047|500174449|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3409|Yellow||2007-04-30|2007-04-30|2016-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||112||1|1|1|1|M|Black||16||Mother|28206|Two Parent|Less than $10,000|||Y|No||Self|General Community||Match Support|M|White||36|28203|||Retail: Sales|28226|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017777|500783368|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
501867805|501645507|500388447|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|298|Green|Amachi|2009-09-27|2009-09-27|2010-07-22|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||9.8||1|1|2|2|M|Black||16|Yes|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|Black||52|28107|Some College|Divorced|Tech: Engineer|28262|3|0|Local Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501868178|31|0|1|31|0|1|5|2|500003586||4|1||-2||-2|0|10|||7437|1|||1|500000294
503296945|503381327|500687021|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|754|Green||2013-03-11|2013-03-13|2015-04-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.8||1|1|1|1|M|Black||16|Yes|Mother|28273|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||43|29707|Bachelors Degree|Separated|Govt||10|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503298770|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502725760|502687867|500589763|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|975|Yellow|Amachi|2012-01-04|2012-01-23|2014-09-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||32||1|1|1|1|M|Black||16|Yes|Mother|28273|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community|Amachi|Match Support|M|Black||28|28226|Bachelors Degree|Single|Business: Sales|28217|0|2|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502726656|31|0|1|31|0|1|10|2|-2||4|2|500000294|-2||-2|0|10|||4748|14|633|1|1|500000294
500191104|501610596|500427661|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|264|Green||2010-01-19|2010-01-29|2010-10-20|Child/Family: Moved|Child/Family: Moved||8.7||3|3|2|2|M|Black||16|No|Mother|28025|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||42|28027|Bachelors Degree|Single|Finance|28262|0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500002335|500191107|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||7464|9|||1|
500191104|501579814|500358644|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|217|Green||2009-04-21|2009-05-01|2009-12-04|Volunteer: Time constraint|Volunteer: Time constraint||7.1||3|3|1|1|M|Black||16|No|Mother|28025|One Parent: Female|Unknown||||No||Neighbor/Friend|General Community||Match Support|M|Black||35|28027|Bachelors Degree|Single|Finance: Banking||0|6|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|500191107|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|8|||7446|3|||1|
502760967|502666332|500579826|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1925|Green||2011-11-18|2011-12-08|NaT||||63.2||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|$25,000 to $29,999|||Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||29|28120|Bachelors Degree|Single|Govt: Clerical||0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|502761879|31|0|2|31|0|2|10|2|-2||2|1|500005291|-2||-2|2203|12|||7464|9|||1|
502177629|502247130|500495930|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|329|Yellow||2010-11-17|2010-11-30|2011-10-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.8||1|1|1|1|M|Black||16|No|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community||RTBM|M|White||59|28277|Associate Degree|Divorced|Unknown||0|0|CIAA Tournament|Special Event|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011184|502178058|31|0|1|1|0|1|7|2|-2||4|2||-2|500000294, 500004640|-2|0|10|||11248|8|||1|
501631140|501628976|500367187|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2451|Green||2009-06-02|2009-06-17|2016-03-03|Volunteer: Moved|Volunteer: Moved||80.5||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||37|28209|Bachelors Degree|Single|Service: Hotel|28202|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501631463|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503149009|503199095|500696674|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|775|Red||2013-05-13|2013-06-13|2015-07-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||25.5||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|$15,000 to $19,999|Yes: Active|Yes|Y|Yes|AARTF|Neighbor/Friend|General Community||Match Support|F|Black||37|28269|Masters Degree|Single|Business: Human Resources|28262|1|3|Recruitment Event|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503150686|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|6855|8|||7460|12|||1|
500740296|500928282|500181834|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1549|Yellow||2007-06-21|2007-06-25|2011-09-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||50.9||2|2|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community||Match Support|F|Black||33|28269|Bachelors Degree|Single|Human Services: Non-Profit||0|6|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500740560|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|5|||7671|13|||1|
500740296|502893901|500611525|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1777|Yellow||2012-04-24|2012-05-04|NaT||||58.4||2|2|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community||Match Support|F|Asian||32|28216|Bachelors Degree|Single|Business: Mgt, Admin|28208|0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|500740560|31|0|2|4|0|2|10|2|-2||2|2||-2||-2|0|5|||7464|9|||1|
501904094|501342148|500420809|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1251|Red||2009-12-11|2010-01-15|2013-06-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||41.1||1|1|1|1|F|Black||16|No|Mother|28214|One Parent: Female|Unknown|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||56|28208|Some College|Single|Finance: Accountant|28203|19|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500004169|501904482|31|0|2|31|0|2|10|2|-2||4|3||-2|500000294|-2|34|2|||7446|3|||1|
502234504|502129464|500463451|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2423|Yellow|Project Big|2010-07-28|2010-07-28|NaT||||79.6||1|1|2|2|F|Black||16|No|GrandMother|28208|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community|Project Big|Match Support|F|Black||37|28216|Bachelors Degree|Single|Customer Service||8|0|LPL Financial|Workplace Partner|Big|General Site||Match Support|0|1|0|1|277|60|598|500000170|500008321|502234935|31|0|2|31|0|2|10|2|500004641||2|2|500004640|-2||-1|0|4|||11247|3|1204|3|1|500004640
502652785|502619698|500548958|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|252|Yellow|2010-2012 OJJDP JJI|2011-08-08|2011-08-19|2012-04-27|Volunteer: Time constraint|Volunteer: Time constraint||8.3||1|1|1|1|M|Multi-race (Black & Hispanic)||16|No|Mother|28270|One Parent: Female|$40,000 to $44,999||||No|Arby's|Workplace Partner/Business|General Community|2010-2012 OJJDP JJI|RTBM|M|Some Other Race||43|28210|Associate Degree|Married|Finance: Banking|28204|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500001281|502653521|38|0|1|41|0|1|7|2|-2||4|2|500005291|-2||-1|3394|14|||7462|13|||1|500005291
502262725|502231024|500467811|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|234|Yellow||2010-08-27|2010-08-30|2011-04-21|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.7||1|1|2|2|F|Black||16|No|Mother|28217|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||29|28277|Bachelors Degree|Single|Consultant|28204|0|11|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011639|502263157|31|0|2|1|0|2|5|2|-2||4|2||-2|500000294|-2|6854|8|||46|2|||1|
500960992|500904815|500193937|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|743|Green||2007-09-06|2007-09-20|2009-10-02|Volunteer: Time constraint|Volunteer: Time constraint||24.4||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|F|White||40|28205|Masters Degree|Single|Business: Sales|17405|0|6|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500961262|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7459|10|||1|
501225346|501412131|500325871|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|531|Green||2008-12-11|2009-01-15|2010-06-30|Child/Family: Moved|Child/Family: Moved||17.4||1|1|1|1|M|Multi-race (Black & Hispanic)||16|No|Mother|27401|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||34|29640|Juris Doctorate (JD)|Single|Law: Lawyer|28226|1|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501225622|38|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502171910|502141964|500460627|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1852|Red|Amachi|2010-07-12|2010-07-30|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||60.8||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Black||42|28214|Some College|Married|Medical||3|6|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500015820|502172339|31|0|1|31|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|5|||7464|9|||1|500000294
502866475|502961396|500614954|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1758|Green||2012-05-15|2012-05-23|NaT||||57.8||1|1|1|1|M|Black||16|No|Mother|28270|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|White||29|28203|Bachelors Degree||Finance: Accountant||1|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502867876|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
500544921|502079132|500523387|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Red|Amachi, Project Big, Project Big AND Amachi|2011-03-07|2011-03-31|2013-08-29|Child: Lost interest|Child: Lost interest||29||2|2|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$15,000 to $19,999|||Y|No|TV|Media|General Community|Project Big AND Amachi|Match Support|M|White||31|28211|Bachelors Degree|Married|Finance: Banking|28202|0|2|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011746|500545173|31|0|1|1|0|1|10|2|500004772||4|3|500004901|-2||-2|56|1|||7464|9|||1|500000294, 500004640, 500004901
500540847|500866129|500181618|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1422|Green|Amachi|2007-06-20|2007-07-02|2011-05-24|Volunteer: Moved|Volunteer: Moved||46.7||2|2|1|1|F|Black||16|Yes|Mother|28208|One Parent: Female|$20,000 to $24,999|||Y|No||Service Organization|General Community|Amachi|Match Support|F|Black||41|28216|||Finance: Accountant||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500541089|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|11|||2238|7|||1|500000294
502088477|502013648|500451408|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|92|Green||2010-05-05|2010-05-24|2010-08-24|Child/Family: Moved|Child/Family: Moved||3||1|1|1|1|M|Black||16|Yes|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Black||35|28210|||Personal Trainer/Coach||0|0|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500010355|502070907|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|
502630686|502630052|500552346|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1069|Yellow|Amachi, Project Big AND Amachi|2011-08-29|2011-09-02|2014-08-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.1||1|1|1|1|M|Black||16|Yes|Mother|28216|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|Amachi|Match Support|M|Multi-race (Black & Hispanic)||39|28208|Bachelors Degree|Single|Business: Marketing||1|6|Recruitment Event|BBBS Board/Staff|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500015820|502631341|31|0|1|38|0|1|10|2|500003586||4|2|500000294|-2|500005291|-2|0|5|||7462|13|||1|500000294, 500004901
502681369|502726053|500568638|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|673|Green|2010-2012 OJJDP JJI|2011-10-21|2011-10-26|2013-08-29|Child: Lost interest|Child: Lost interest||22.1||1|1|1|1|F|White||16|No|Mother|28262|One Parent: Female|$25,000 to $29,999||||No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||36|28205|Bachelors Degree|Single|Business: Human Resources|28202|4|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502682197|1|0|2|1|0|2|10|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|500005291
503983132|503995895|500791249|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|850|Green|PERL 2014-2016|2014-11-03|2014-11-17|NaT||||27.9||1|1|1|1|M|Black||16|Yes|GrandMother|28270|One Parent: Female|$15,000 to $19,999|||Y|No||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||49|28226|Juris Doctorate (JD)|Married|Law: Lawyer|28202|4|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|503985143|31|0|1|1|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|0|5|||46|2|||1|500014681
502590651|502589724|500542166|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|784|Red|Project Big, 2010-2012 OJJDP JJI|2011-06-20|2011-06-30|2013-08-22|Volunteer: Time constraint|Volunteer: Time constraint||25.8||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||36|28205|Bachelors Degree|Single|Business: Marketing|28117|7|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011746|502591168|31|0|2|1|0|2|10|2|500004641||4|3|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291
502538068|502672354|500554099|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|126|Green||2011-09-12|2011-09-27|2012-01-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||4.1||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||28|28215||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502538521|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
503597088|503642924|500731612|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|879|Green||2013-11-15|2013-12-06|2016-05-03|Volunteer: Moved|Volunteer: Moved||28.9||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Retail: Sales|28217|0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503598965|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500363212|500797130|500176231|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2014|Green|Amachi|2007-05-09|2007-05-24|2012-11-27|Volunteer: Moved|Volunteer: Moved||66.2||2|2|1|1|F|Multi-Race (None of the above)||16||Mother|28025|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||34|28211|Associate Degree|Living w/ Significant Other|Business: Clerical|28211|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500013781|500188099|7|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
500363209|500371073|500099752|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1681|Green|Amachi|2006-05-24|2006-05-24|2010-12-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||55.2||1|1|1|1|F|Multi-Race (None of the above)||16|Yes|Mother|28025|Other/Unknown|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||57|28262||Married|Finance: Banking||0|9|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188099|7|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500918264|501074231|500236477|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1476|Yellow||2008-01-09|2008-02-13|2012-02-28|Child: Severity of challenges|Child: Severity of challenges||48.5||1|1|1|1|M|Multi-Race (None of the above)||16|No|Mother|28227|Two Mothers|$45,000 to $49,999||||No||Self|General Community||Match Support|M|Black||33|28269|Some College|Single|Business: Clerical||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500918534|7|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
502210299|501993351|500456811|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|411|Green||2010-06-15|2010-06-16|2011-08-01|Volunteer: Moved|Volunteer: Moved||13.5||1|1|1|1|M|Hispanic||16|No|Mother|28213|Two Parent: Not Married|Unknown|||Y|Yes||School|General Community||RTBM|M|White||39|28209|||Transport: Pilot||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|502210728|3|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502478428|502555822|500533009|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2149|Green|2010-2012 OJJDP JJI|2011-04-23|2011-04-28|NaT||||70.6||1|1|1|1|M|White||16|No|Mother|28277|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||54|28205|Some College|Separated|Self-Employed, Entrepreneur|28214|29|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502478875|1|0|1|1|0|1|10|2|-2||2|1|500005291|-2||-2|0|10|||7464|9|||1|500005291
501919692|502219683|500465111|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|595|Red||2010-08-10|2010-08-13|2012-03-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.5||1|1|1|1|M|White||16|No|Mother|28270|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|White||35|28270|Associate Degree|Married|Firefighter||1|6|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013709|501920088|1|0|1|1|0|1|5|2|-2||4|3||-2|500000294|-2|0|10|||7464|9|||1|
503496889|503490051|500708903|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|611|Green||2013-09-03|2013-09-25|2015-05-29|Volunteer: Moved|Volunteer: Moved||20.1||1|1|1|1|M|Black||16|No|Mother|28273|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||28|28207|Bachelors Degree|Single|Education: Teacher||1|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503498757|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502939293|502855925|500632744|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|423|Red||2012-09-06|2012-09-24|2013-11-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||13.9||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|F|White||48|28269|Bachelors Degree|Single|Finance: Banking||18|0|Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502940718|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|4|||131|1|||1|
501597228|501397328|500379964|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2750|Green|Amachi|2009-08-19|2009-09-04|NaT||||90.3||1|1|1|1|F|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||40|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28204|0|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501597548|31|0|2|31|0|2|10|2|500003586||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
502319984|502290677|500607367|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1058|Red||2012-03-30|2012-04-30|2015-03-24|Volunteer: Time constraint|Volunteer: Time constraint||34.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|28203|Bachelors Degree|Single|Finance|28216|3|0|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502320419|31|0|1|1|0|1|10|2|-2||4|3|500005291|-2||-2|6854|8|||17161|11|||1|
502138562|502380370|500502780|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|905|Green||2010-12-07|2010-12-14|2013-06-06|Child: Lost interest|Child: Lost interest||29.7||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||38|28216|Masters Degree|Single|Finance: Auditor|28217|3|0|100 Men in 100 Days|Fraternity/Sorority|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502138991|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||12183|14|||1|
503556265|503498990|500715926|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|286|Green||2013-10-04|2013-10-18|2014-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||9.4||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Enrollment|F|Black||42|28216|Bachelors Degree|Single|Business: Mgt, Admin|28210|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503558140|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502537469|502227984|500534571|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|485|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-05-02|2011-05-04|2012-08-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||15.9||3|3|1|1|F|Black||16|No|Mother|28208|One Parent: Female|$15,000 to $19,999||||No||School|General Site||Match Support|F|White||38|28205|Bachelors Degree|Divorced|Customer Service||1|3|TV|Media|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500001281|502537922|31|0|2|1|0|2|10|2|500004641||4|2||-1|500004640|-2|0|4|||130|1|1204|3|1|500004640, 500005291
502537469|503323641|500702088|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|751|Green||2013-06-26|2013-07-17|2015-08-07|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||24.7||3|3|2|2|F|Black||16|No|Mother|28208|One Parent: Female|$15,000 to $19,999||||No||School|General Site||Match Support|F|White||34|28078|Masters Degree|Single|Medical: Doctor, Provider|28001|0|2|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|502537922|31|0|2|1|0|2|10|2|-2||4|1||-1|500007920, 500011315, 500011316|-2|0|4|||46|2|||1|
502240203|502110142|500460976|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|370|Green|Amachi|2010-07-14|2010-07-23|2011-07-28|Volunteer: Moved|Volunteer: Moved||12.2||2|2|1|1|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||||Yes||Self|General Community|Amachi|RTBM|F|Black||38|28262|Bachelors Degree|Single|Finance: Banking||5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502240634|31|0|2|31|0|2|7|2|||4|1|500000294|-2|500000294|-2|0|10|||7496|10|||1|500000294
502240203|502668316|500556356|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|182|Yellow||2011-09-20|2011-09-29|2012-03-29|Volunteer: Time constraint|Volunteer: Time constraint||6||2|2|1|1|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||||Yes||Self|General Community|Amachi|RTBM|F|Black||31|28216||Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502240634|31|0|2|31|0|2|7|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|
502240205|502657850|500553471|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|993|Green|Amachi|2011-09-07|2011-09-22|2014-06-11|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||32.6||3|3|2|2|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||48|28203|Bachelors Degree|Married|Business: Mgt, Admin|28202|1|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002334|502240634|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
502240205|502203053|500460610|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|57|Yellow||2010-07-12|2010-07-15|2010-09-10|Volunteer: Time constraint|Volunteer: Time constraint||1.9||3|3|1|1|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||35|28202|Bachelors Degree|Single|Retail: Sales||0|8|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|502240634|31|0|2|1|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1|
502240205|502249748|500472560|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|297|Green|Amachi|2010-09-22|2010-10-04|2011-07-28|Volunteer: Moved|Volunteer: Moved||9.8||3|3|1|1|F|Black||16|Yes|GrandMother|28216|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||31|28209|Bachelors Degree|Single|Business: Sales|28092|0|3|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502240634|31|0|2|1|0|2|10|2|||4|1|500000294|-2|500000294|-2|0|10|||46|2|||1|500000294
501143674|502958999|500612879|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1550|Yellow||2012-05-01|2012-05-08|2016-08-05|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||50.9||3|3|1|1|F|Black||16||Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||28|28211|Bachelors Degree|Single|Human Services||2|0|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501143948|31|0|2|1|0|2|10|2|500004641||4|2||-2||-2|0|10|||132|8|||1|
500826100|502605848|500549342|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|307|Green|2010-2012 OJJDP JJI|2011-08-10|2011-08-26|2012-06-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||10.1||4|4|1|1|F|Black||16|No|Mother|28213|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||RTBM|F|White||41|28204|Bachelors Degree|Divorced|Retail: Mgt|28027|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|500801835|31|0|2|1|0|2|7|2|-2||4|1||-2||-2|0|10|||7496|10|||1|500005291
500826100|500648169|500167025|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1325|Green||2007-03-15|2007-03-21|2010-11-05|Volunteer: Moved|Volunteer: Moved||43.5||4|4|1|1|F|Black||16|No|Mother|28213|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||RTBM|F|Black||37|28262|Masters Degree|Single|Finance: Accountant||0|0|General|Other Big|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500801835|31|0|2|31|0|2|7|2|-2||4|1||-2||-2|0|10|||6450|12|||1|
500826100|503877762|500774526|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|201|Green||2014-09-04|2014-09-19|2015-04-08|Volunteer: Moved|Volunteer: Moved||6.6||4|4|1|1|F|Black||16|No|Mother|28213|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||RTBM|F|Black||30|28269|Masters Degree|Single|Medical||0|11|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500011349|500801835|31|0|2|31|0|2|7|2|-2||4|1||-2|500000294|-2|0|10|||46|2|||1|
500826100|502225881|500501827|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|140|Green||2010-12-03|2010-12-10|2011-04-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.6||4|4|1|1|F|Black||16|No|Mother|28213|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||RTBM|F|Black||26|28269||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|500801835|31|0|2|31|0|2|7|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502185085|502335257|500482493|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|184|Yellow||2010-10-19|2010-10-30|2011-05-02|Child: Lost interest|Child: Lost interest||6||1|1|2|2|M|White||16|No|Mother|28031|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||53|28117|Bachelors Degree|Married|Real Estate: Realtor|28031|0|0|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|502185514|1|0|1|1|0|1|10|2|-2||4|2||-2|500000294, 500004901|-2|6854|8|||7464|9|||1|
500910037|500856100|500368834|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2824|Green||2009-06-15|2009-06-22|NaT||||92.8||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Match Support|M|White||46|28277||Married|Business: Mgt, Admin||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|500910307|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
500843863|501078655|500241388|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3039|Green|Amachi|2008-01-31|2008-02-21|2016-06-17|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||99.8||2|2|1|1|F|Black||16|Yes|Mother|28217|One Parent: Female|$15,000 to $19,999|||Y|No|TV|Media|General Community|Amachi|Match Support|F|Black||32|28269|Bachelors Degree|Single|Business: Marketing|28273|0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500844129|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|56|1|||2238|7|||1|500000294
502567548|502564910|500534824|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|523|Red|Amachi, Project Big AND Amachi|2011-05-03|2011-05-27|2012-10-31|Child/Family: Moved|Child/Family: Moved||17.2||1|1|2|2|F|Hispanic||16|Yes|Mother|28227|One Parent: Female|Unknown||||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||45|28262|Masters Degree|Married|Education|28206|1|0|Relative|Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502568002|3|0|2|31|0|2|10|2|500003586||4|3|500004640, 500004901|-2||-2|0|4|||17161|11|||1|500000294, 500004901
501068953|500874318|500380111|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|907|Green||2009-08-20|2009-10-06|2012-03-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||29.8||2|2|2|2|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||40|28262|Bachelors Degree|Married|Law: Paralegal|28280|4|5|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501060469|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
501068953|501004437|500223479|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|487|Green||2007-11-27|2007-11-27|2009-03-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||16||2|2|2|2|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Black||39|28105|Masters Degree|Single|Business: Mgt, Admin|28204|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|501060469|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
501288021|501249338|500281778|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2714|Green||2008-08-13|2008-08-27|2016-02-01|Volunteer: Moved|Volunteer: Moved||89.2||1|1|1|1|F|Black||16|No|Mother|28211|Two Parent|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||37|28027|PHD|Single|Education: College Professor|27411|1|8|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500018851|501288299|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
500936718|501027885|500224574|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3101|Green||2007-11-29|2007-12-20|2016-06-16|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||101.9||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28210|Bachelors Degree|Married|Business: Sales||0|4|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|1|0|0|1|277|60|598|500000170|500017732|500915629|31|0|1|1|0|1|10|2|-2||4|1||-2|500014505, 500015184|-1|34|2|||46|2|||1|
501825910|501196986|500380446|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2587|Yellow|Amachi|2009-08-24|2009-08-24|2016-09-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||85||1|1|1|1|M|Black||16|Yes|Mother|28213|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||51|28214|Masters Degree|Married|Business: Sales|94108|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|500188141|31|0|1|1|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7496|10|||1|500000294
502610186|502913393|500601697|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1816|Green||2012-03-01|2012-03-26|NaT||||59.7||1|1|1|1|F|Black||16|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Asian||35|28210|Masters Degree|Married|Arts, Entertainment, Sports|28202|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502610737|31|0|2|4|0|2|10|2|-2||2|1||-2||-2|6854|8|||7671|13|||1|
502896701|502888938|500610476|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|364|Yellow||2012-04-18|2012-04-30|2013-04-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12||1|1|1|1|M|Black||16|No|Mother|28214|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|White||64|28216|Juris Doctorate (JD)|Divorced|Law: Lawyer||3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502898109|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503187841|503789478|500762532|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|767|Green||2014-05-07|2014-05-15|2016-06-20|Child/Family: Moved|Child/Family: Moved||25.2||1|1|1|1|M|White||16||Mother|28277|One Parent: Female|$40,000 to $44,999|||Y|No||Self|General Community||Match Support|M|White||60|28105|Bachelors Degree|Married|Tech: Research/Design|28277|4|0|Recruitment Event|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503189585|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7460|12|||1|
501604887|501743226|500373295|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|366|Red||2009-07-09|2009-07-27|2010-07-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12||2|2|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Site|Amachi|Match Support|M|White||26|28270|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501605207|31|0|1|1|0|1|10|2|-2||4|3|500000294|-1|500000294|-2|0|10|||46|2|||1|
503262762|503114924|500678106|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|340|Red||2013-01-29|2013-01-31|2014-01-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.2||1|1|1|1|F|Black||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||29|28203|Bachelors Degree|Single|Education: Teacher|28031|1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503264570|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
500465506|500496966|500118121|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3860|Yellow|Amachi|2006-08-15|2006-08-21|NaT||||126.8||1|1|1|1|M|Black||16|Yes|Mother|28262|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community|Amachi|Match Support|M|White||54|28226|Bachelors Degree|Married|Arts, Entertainment, Sports||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500465757|31|0|1|1|0|1|10|2|500003586||2|2|500000294|-2|500000294|-2|0|4|||2238|7|||1|500000294
501990745|502098002|500447817|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|838|Red||2010-04-19|2010-05-14|2012-08-29|Child: Severity of challenges|Child: Severity of challenges||27.5||1|1|1|1|M|Black||16||Mother|28269|One Parent: Female|Unknown||||Yes||BBBS Board/Staff|General Community||Match Support|M|Black||35|28213||Married|Human Services: Youth Worker||0|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501991144|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|13|||4748|14|||1|
502666718|500932879|500548835|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|706|Red|2010-2012 OJJDP JJI|2011-08-05|2011-08-19|2013-07-25|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||23.2||1|1|2|2|F|Black||16|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||38|28202|Masters Degree||Business: Clerical||7|0|Recruitment Event|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502667545|31|0|2|31|0|2|10|2|-2||4|3|500005291|-2||-2|0|10|||7458|9|||1|500005291
501353940|501587399|500360226|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|712|Yellow|Amachi|2009-04-29|2009-05-29|2011-05-11|Volunteer: Time constraint|Volunteer: Time constraint||23.4||3|3|1|1|M|Black||16|No|Relative: Other|28205|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||35|28211||Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|501354219|31|0|1|1|0|1|10|2|500003586||4|2|500000294, 500005291|-2||-2|34|2|||7464|9|||1|500000294
501353940|502710990|500574615|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1933|Green|Amachi|2011-11-04|2011-11-30|NaT||||63.5||3|3|1|1|M|Black||16|No|Relative: Other|28205|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||33|28226|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|10|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501354219|31|0|1|1|0|1|10|2|500003586||2|1|500000294, 500005291|-2||-2|34|2|||17161|11|||1|500000294
501353940|501317674|500287832|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|120|Green|Amachi|2008-09-12|2008-09-23|2009-01-21|Volunteer: Moved|Volunteer: Moved||3.9||3|3|1|1|M|Black||16|No|Relative: Other|28205|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI, Amachi|Match Support|M|White||31|28211|Bachelors Degree|Single|Business: Clerical|28210|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501354219|31|0|1|1|0|1|10|2|500003586||4|1|500000294, 500005291|-2||-2|34|2|||7496|10|||1|500000294
502064627|500773055|500462574|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2400|Green||2010-07-26|2010-08-20|NaT||||78.9||1|1|2|2|M|Black||16|No|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Hispanic|Other Central American|37|28204||Single|Construction||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502065051|31|0|1|3|14|1|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
502997211|502926434|500614826|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|461|Yellow||2012-05-15|2012-06-01|2013-09-05|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||15.1||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|F|White||27|28105|Some College||Student: College||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011349|502998689|31|0|2|1|0|2|7|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502482642|502601273|500541388|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|405|Red|Project Big, 2010-2012 OJJDP JJI|2011-06-15|2011-06-22|2012-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.3||2|2|1|1|F|Black||16|No|Mother|28052|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||30|28204|Masters Degree|Single|Finance: Auditor|28202|2|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502391834|31|0|2|1|0|2|10|2|-2||4|3|500004640, 500005291|-2|500004640|-2|0|10|||7496|10|||1|500004640, 500005291
502482642|503118336|500679560|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|858|Yellow||2013-02-04|2013-02-11|2015-06-19|Child/Family: Moved|Child/Family: Moved||28.2||2|2|1|1|F|Black||16|No|Mother|28052|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||29|28277|Bachelors Degree|Single|Business|28217|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|502391834|31|0|2|1|0|2|10|2|-2||4|2|500004640, 500005291|-2||-2|0|10|||7464|9|||1|
502264006|502274748|500470897|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2349|Red||2010-09-16|2010-09-22|2017-02-26|Child: Lost interest|Child: Lost interest||77.2||1|1|1|1|F|Hispanic||16|No|Mother|28211|One Parent: Female|Unknown||||Yes|Spanish Print|Media|General Community||Match Support|F|Hispanic||38|28202|Bachelors Degree|Single|Tech: Engineer|28202|12|0|Big Day|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502264438|3|0|2|3|0|2|10|2|-2||4|3||-2||-2|7063|1|||7456|8|||1|
501525308|501536144|500335230|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2313|Green||2009-01-23|2009-02-16|2015-06-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||76||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|White||40|28205|Some College|Married|Retail: Sales|28206|1|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|501525600|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|6854|8|||7464|9|||1|
502198485|500188656|500508298|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|644|Red|Amachi|2010-12-28|2011-01-12|2012-10-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||21.2||1|1|2|2|M|Black||16|Yes|Mother|28262|One Parent: Female|Unknown||||Yes||School|General Community|Amachi|Match Support|M|Black||53|28262|Some College|Married|Business: Clerical||0|0|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500012459|502198914|31|0|1|31|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|4|||7464|9|||1|500000294
501074345|501158523|500250038|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3272|Green|Amachi, Cabarrus County|2008-03-04|2008-03-31|NaT||||107.5||1|1|1|1|M|White||16|Yes|GrandMother|28025|Grandparents|Unknown||||No|Other|Faith Organization|General Community|Amachi, Cabarrus County|Match Support|M|White||46|28027|Bachelors Degree|Divorced|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|501074618|1|0|1|1|0|1|10|2|500003586||2|1|500000294, 500016374|-2|500016374|-2|5635|9|||46|2|||1|500000294, 500016374
501249953|501292229|500278068|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|568|Red||2008-07-16|2008-08-14|2010-03-05|Child: Lost interest|Child: Lost interest||18.7||1|1|1|1|M|Multi-race (Black & White)||16|No|Mother|28226|One Parent: Female|Unknown||||No|TV|Media|General Community||Match Support|M|White||33|28277|Bachelors Degree|Living w/ Significant Other|Finance: Economist|28277|2|0|Coworker|Workplace Partner|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500009007|501250229|36|0|1|1|0|1|10|2|-2||4|3||-2||-2|56|1|||7447|3|||1|
502753870|502785389|500574313|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1065|Yellow||2011-11-03|2011-11-30|2014-10-30|Volunteer: Time constraint|Volunteer: Time constraint||35||2|2|1|1|F|Hispanic||16|No|Mother|28262|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|F|White||31|28210|Masters Degree|Single|Medical: Doctor, Provider||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502751081|3|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
502753870|503869569|500794392|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|598|Red||2014-11-11|2014-12-08|2016-07-28|Child: Lost interest|Child: Lost interest||19.6||2|2|2|2|F|Hispanic||16|No|Mother|28262|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|F|White||26|28210|Bachelors Degree|Single|Medical: Admin|28209|1|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500013781|502751081|3|0|2|1|0|2|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|
502549829|502594393|500541795|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2086|Green|Amachi, Project Big, Project Big AND Amachi|2011-06-16|2011-06-30|NaT||||68.5||1|1|1|1|M|Black||16|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|Amachi, PERL 2014-2016, Project Big, Project Big AND Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Business: Engineer|30357|6|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502550279|31|0|1|31|0|1|10|2|500004772||2|1|500000294, 500004640, 500004901, 500014681|-1||-2|0|4|||7464|9|||1|500000294, 500004640, 500004901
501957505|501718938|500432245|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|765|Green|Amachi|2010-02-03|2010-02-25|2012-03-31|Volunteer: Moved|Volunteer: Moved||25.1||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||55|28078|||Business: Marketing|28070|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501957903|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|500000294
501165117|503119136|500690258|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|217|Red||2013-03-27|2013-03-28|2013-10-31|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.1||2|3|1|1|F|Black||16||Mother|28205|Other/Unknown|Unknown||||Yes||Self|General Community||Enrollment|F|White||33|28209|Bachelors Degree|Single|Human Services: Non-Profit||6|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|501165391|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500934908|500856560|500218659|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|533|Green|Amachi|2007-11-15|2007-12-03|2009-05-19|Volunteer: Moved|Volunteer: Moved||17.5||2|2|1|1|M|Black||16|Yes|Aunt|28216|One Parent: Female|Less than $10,000|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||50|28262||Married|Business: Sales||1|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500935173|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|5635|9|||2238|7|||1|500000294
500934908|502107314|500456443|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2463|Green|Amachi|2010-06-11|2010-06-18|NaT||||80.9||2|2|1|1|M|Black||16|Yes|Aunt|28216|One Parent: Female|Less than $10,000|||Y|No|Other|Faith Organization|General Community|Amachi|Match Support|M|White||34|20175|Bachelors Degree|Single|Business: Sales|28211|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|500935173|31|0|1|1|0|1|10|2|500003586||2|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
502248736|502266779|500472618|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|120|Green||2010-09-22|2010-10-11|2011-02-08|Volunteer: Health|Volunteer: Health||3.9||1|1|1|1|M|Black||16|No|Mother|28027|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|Black||61|28027||Single|Business: Marketing||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|502249167|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502393980|502928199|500613992|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1756|Green|Amachi|2012-05-09|2012-05-25|NaT||||57.7||2|2|1|1|F|Multi-race (Black & White)||16|Yes|Aunt|28269|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||54|28078|Associate Degree|Married|Tech: Support, Writing|28210|2|6|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502394418|36|0|2|31|0|2|10|2|500003586||2|1|500005291|-2||-2|0|5|||7462|13|||1|500000294
502393980|502454075|500554127|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|213|Green|Amachi|2011-09-12|2011-09-30|2012-04-30|Volunteer: Time constraint|Volunteer: Time constraint||7||2|2|1|1|F|Multi-race (Black & White)||16|Yes|Aunt|28269|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||31|28078|Some College|Married|Medical: Healthcare Worker|28262|0|6|Big Champions|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502394418|36|0|2|31|0|2|10|2|-2||4|1|500005291|-2||-2|0|5|||7461|12|||1|500000294
502931305|502500246|500608719|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|95|Green||2012-04-09|2012-04-27|2012-07-31|Child: Family structure changed|Child: Family structure changed||3.1||1|1|2|2|M|Black||16|No|Mother|28214|One Parent: Female|$100,000 to $124,999||||No||Self|General Community||Match Support|M|White||31|28269|Masters Degree|Single|Insurance|28262|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502932726|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
502670071|502685522|500557057|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|876|Yellow|Amachi, 2010-2012 OJJDP JJI|2011-09-22|2011-10-26|2014-03-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.8||1|1|1|1|F|Black||16|Yes|Mother|28083|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|F|Black||36|28269|Masters Degree|Single|Human Services: Youth Worker|28027|2|2|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502670906|31|0|2|31|0|2|5|2|500003586||4|2|500005291|-2||-2|0|10|||9229|13|||1|500000294, 500005291
502380578|502138981|500579112|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|905|Yellow||2011-11-17|2011-11-22|2014-05-15|Child/Family: Moved|Child/Family: Moved||29.7||2|2|3|3|F|Black||16||Mother|28213|Other/Unknown|Unknown||||Yes||School|General Community||Match Support|F|Black||29|28262|Bachelors Degree|Single|Student: College||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502381016|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|4|||7496|10|||1|
500280148|500865221|500179364|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|849|Green|Amachi|2007-06-07|2007-06-13|2009-10-09|Volunteer: Time constraint|Volunteer: Time constraint||27.9||3|3|1|1|F|Black||16|Yes|Mother|28205|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|F|Black||37|28216|Some College|Single|Business: Clerical||3|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500003657|500188151|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|3|||2238|7|||1|500000294
500280148|502118494|500460767|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2438|Yellow|Amachi|2010-07-13|2010-07-13|NaT||||80.1||3|3|1|1|F|Black||16|Yes|Mother|28205|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|F|Black||30|28216|Bachelors Degree|Single|Human Services: Non-Profit|28216|0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|500188151|31|0|2|31|0|2|10|2|500003586||2|2|500000294|-2||-2|0|3|||7464|9|||1|500000294
502530223|502501248|500533054|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|753|Red|2010-2012 OJJDP JJI|2011-04-25|2011-04-29|2013-05-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||24.7||1|1|1|1|M|Hispanic||16||Mother|28213|One Parent: Female|Unknown||||No||School|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||44|28078|Masters Degree|Married|Business|28036|8|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502530676|3|0|1|3|0|1|10|2|-2||4|3|500005291|-2||-2|0|4|||7464|9|||1|500005291
502495214|502346954|500519656|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|395|Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|2011-02-23|2011-02-28|2012-03-29|Volunteer: Time constraint|Volunteer: Time constraint||13||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||61|28056||Married|Medical: Pharmacist||0|0|Healthy Kids Club|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502495663|31|0|2|31|0|2|10|2|500004772||4|2|500004640, 500005291|-2||-2|0|4|459|3|10326|3|||1|500000294, 500004640, 500004901, 500005291
502593613|502601730|500547881|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2020|Yellow||2011-07-28|2011-08-19|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||66.4||1|1|1|1|F|Black||16|No|Mother|28208|Two Parent|$35,000 to $39,999|||Y|Yes||Relative|General Community||Match Support|F|Hispanic||26|28217|Bachelors Degree|Single|Service: Restaurant||3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502594130|31|0|2|3|0|2|10|2|-2||4|2||-2||-2|0|3|||7464|9|||1|
503225805|503317460|500680855|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1173|Red||2013-02-08|2013-03-08|2016-05-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38.5||1|1|1|1|F|White||16|No|Mother|28082|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|F|White||33|28138|Associate Degree|Divorced|Insurance||2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503227593|1|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
501305368|501174923|500339693|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|522|Green||2009-02-09|2009-03-09|2010-08-13|Volunteer: Time constraint|Volunteer: Time constraint||17.1||2|2|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|Black||70|28078|Bachelors Degree|Married|Retired||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501305646|31|0|1|31|0|1|7|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501305368|502665365|500552025|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|649|Green||2011-08-26|2011-09-09|2013-06-19|Volunteer: Moved|Volunteer: Moved||21.3||2|2|1|1|M|Black||16|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||29|28202|Bachelors Degree|Single|Finance: Banking|28202|0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|501305646|31|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
503459852|503208612|500703588|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|418|Green||2013-07-15|2013-07-31|2014-09-22|Volunteer: Time constraint|Volunteer: Time constraint||13.7||1|1|1|1|F|Hispanic||16|No|Mother|28078|One Parent: Female|Less than $10,000||||Yes|BBBS National Site|Web Link|General Community||RTBM|F|Hispanic||28|28031|Bachelors Degree||Business|28202|0|2|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503461718|3|0|2|3|0|2|7|2|-2||4|1||-2||-2|34|2|||46|2|||1|
502304267|503343217|500682425|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1282|Yellow||2013-02-15|2013-02-27|2016-09-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||42.1||2|2|1|1|M|White||16|No|Mother|28277|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||47|28277|Bachelors Degree|Married|Business|28217|20|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502304699|1|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7671|13|||1|
502304267|502301421|500483429|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|713|Red||2010-10-20|2010-10-28|2012-10-10|Volunteer: Moved|Volunteer: Moved||23.4||2|2|1|1|M|White||16|No|Mother|28277|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||32|28270|Masters Degree|Living w/ Significant Other|Unemployed||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502304699|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
500267459|500464544|500121193|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2353|Red||2006-09-07|2006-09-19|2013-02-27|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||77.3||1|1|1|1|M|Black||16||Mother|28203|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||39|28202|Bachelors Degree|Single|Finance: Accountant||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011746|500187395|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
500727291|500857838|500176403|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3361|Green||2007-05-10|2007-05-17|2016-07-29|Child: Graduated|Child: Graduated||110.4||1|1|1|1|M|Black||16|No|Mother|28216|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|Black||46|28269|||Human Services: Non-Profit||0|0|BBBS National Site|Web Link|Big|General Community|VOL - Adjudicated, VOL - Cultural Comp, VOL - PreMatch|Match Support|1|0|0|1|277|60|598|500000170|500008321|500727558|31|0|1|31|0|1|10|2|-2||4|1||-2|500007913, 500007920, 500011311|-2|0|10|||46|2|||1|
501614040|501864748|500404360|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1205|Red||2009-11-02|2009-11-11|2013-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||39.6||1|1|1|1|M|Hispanic||16|No|Mother|28273|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||29|28273|||Facilities/Maintenance||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|501614360|3|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502179379|502161458|500461681|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1832|Red|Project Big|2010-07-20|2010-07-25|2015-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||60.2||1|1|1|1|F|Black||16|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|Black||34|28269||Single|Student: College||0|0|UNCC|College Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502179808|31|0|2|31|0|2|10|2|-2||4|3|500004640|-2||-2|0|10|||9221|5|||1|500004640
500417281|500349297|500112798|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2376|Green|Amachi|2006-07-31|2006-07-31|2013-01-31|Volunteer: Time constraint|Volunteer: Time constraint||78.1|Y|1|1|1|1|F|White||16||Mother|28211|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||48|28211|Masters Degree|Married|Finance: Banking|28202|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|500402926|1|0|2|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||2238|7|||1|500000294
503379566|503407492|500697331|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1393|Green|Cabarrus County|2013-05-17|2013-05-23|NaT||||45.8||1|1|1|1|M|Black||16||Mother|28027|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||51|28269|Bachelors Degree|Married|Business: Sales||6|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|503381423|31|0|1|1|0|1|10|2|500016307||2|1|500016374|-2|500016374|-2|34|2|||46|2|||1|500016374
500382177|500188566|500122093|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3263|Yellow||2006-09-14|2006-09-18|2015-08-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||107.2||1|1|2|2|M|Black||16||Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||43|28215|Bachelors Degree|Single|Finance: Banking|28262|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500012459|500382427|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
503472839|503503841|500702872|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|672|Green||2013-07-08|2013-07-26|2015-05-29|Child/Family: Moved|Child/Family: Moved||22.1||1|1|1|1|F|Black||16|Yes|Mother|28214|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||25|28223|Some College|Single|Student: College|28223|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503474705|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501663624|501440384|500349001|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|120|Green||2009-03-11|2009-03-17|2009-07-15|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.9||1|1|1|1|F|White||16|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|F|White||30|28027|Some College|Single|Student: College||0|0|Recruitment Event|College Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001262|501663922|1|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7448|5|||1|
503395663|503735537|500744097|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|594|Green||2014-01-22|2014-02-21|2015-10-08|Volunteer: Moved|Volunteer: Moved||19.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28204|Masters Degree|Single|Finance: Accountant|28202|4|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503397520|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
502495123|502473441|500524205|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|649|Red|Project Big, 2010-2012 OJJDP JJI|2011-03-09|2011-03-31|2013-01-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||21.3||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||34|28207|Bachelors Degree|Single|Finance: Economist|28255|5|0||Relative|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502495572|31|0|2|1|0|2|10|2|500004641||4|3|500004640, 500005291|-2|500004640|-2|0|4|||0|11|||1|500004640, 500005291
502589865|502625828|500544108|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1582|Red|Project Big, 2010-2012 OJJDP JJI|2011-06-30|2011-06-30|2015-10-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||52||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Black||40|28037|Bachelors Degree|Married|Medical: Doctor, Provider||2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502590381|31|0|1|31|0|1|10|2|500004641||4|3|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291
502083450|500863980|500605881|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|559|Yellow||2012-03-23|2012-04-05|2013-10-16|Volunteer: Time constraint|Volunteer: Time constraint||18.4||2|2|3|3|M|Black||16|No|Mother|28027|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||49|28027|Bachelors Degree|Married|Transport: Driver|28208|6|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|0|1|1|0|277|60|598|500000170|500002335|502083874|31|0|1|31|0|1|10|2|-2||4|2|500005291|-2|500014505, 500014506|-1|7016|11|||7671|13|||1|
502083450|502104415|500453680|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|463|Green|Amachi|2010-05-20|2010-05-20|2011-08-26|Volunteer: Time constraint|Volunteer: Time constraint||15.2||2|2|1|1|M|Black||16|No|Mother|28027|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||44|28262||Divorced|Service: Restaurant|28027|0|10|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|502083874|31|0|1|31|0|1|10|2|500003586||4|1|500005291|-2||-2|7016|11|||7464|9|12|3|1|500000294
501428294|501517334|500317955|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1064|Green||2008-11-19|2008-11-25|2011-10-25|Volunteer: Time constraint|Volunteer: Time constraint||35||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|M|Black||40|28209|Associate Degree|Married|Unknown|28208|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501428579|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|6854|8|||7671|13|||1|
502083456|502542333|500548042|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|719|Green||2011-07-29|2011-08-03|2013-07-22|Child/Family: Moved|Child/Family: Moved||23.6||1|1|1|1|F|Black||16|No|Mother|28025|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||29|28262|Masters Degree|Single|Finance: Banking|28208|4|0|Other|BBBS Board/Staff|Big|General Site|mentor2.0 2014|Enrollment|0|1|1|0|277|60|598|500000170|500012459|502083880|31|0|2|31|0|2|10|2|-2||4|1||-2|500014506|-1|0|10|||7671|13|||1|
502310004|502331000|500483762|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1283|Yellow|Amachi, Project Big, Project Big AND Amachi|2010-10-21|2010-10-26|2014-05-01|Volunteer: Moved|Volunteer: Moved||42.2||1|1|1|1|F|Black||16|Yes|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Enrollment|F|White||37|28078||Single|Business||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500015820|502310436|31|0|2|1|0|2|5|2|500003586||4|2|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7496|10|||1|500000294, 500004640, 500004901
503830048|503559585|500757050|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|149|Red||2014-03-27|2014-04-08|2014-09-04|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||4.9||1|1|1|1|F|Hispanic||16|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||47|28205|Associate Degree|Single|Medical: Nurse||1|0|BBBS National Site|Web Link|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500017777|503832027|3|0|2|1|0|2|10|2|-2||4|3||-2||-2|34|2|||46|2|||1|
502260656|502249984|500475564|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|883|Red||2010-09-30|2010-10-18|2013-03-19|Volunteer: Moved|Volunteer: Moved||29||2|2|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28078|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||33|28078|Associate Degree|Married|Education: Teacher Asst/Aid||3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502261088|38|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502260656|502031924|500466370|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|23|Green||2010-08-19|2010-08-30|2010-09-22|Volunteer: Moved|Volunteer: Moved||0.8||2|2|1|1|F|Multi-race (Black & Hispanic)||16|No|Mother|28078|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||32|28025|Bachelors Degree|Single|Customer Service||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|502261088|38|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502545735|502388739|500542256|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|346|Red||2011-06-21|2011-07-12|2012-06-22|Volunteer: Health|Volunteer: Health||11.4||1|1|1|1|M|Multi-race (Hispanic & White)||16|No|Mother|28227|One Parent: Female|$25,000 to $29,999||||No|Big|Neighbor/Friend|General Community||RTBM|M|White||41|28205|Bachelors Degree|Married|Finance|28255|9|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502546188|35|0|1|1|0|1|7|2|-2||4|3||-2||-2|6854|8|||7464|9|||1|
503934189|503918487|500796401|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|842|Green||2014-11-17|2014-11-25|NaT||||27.7||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|White||35|28211|Masters Degree|Single|Finance: Accountant|28202|2|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503936197|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|4|||17101|1|||1|
503556065|501284751|500741332|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|637|Yellow||2014-01-06|2014-01-10|2015-10-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||20.9||1|1|3|3|M|Black||16|No|Mother|28269|One Parent: Female|$50,000 to $59,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||50|28031|Masters Degree|Married|Self-Employed, Entrepreneur||0|0|Bowl For Kids Sake|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017777|503557940|31|0|1|31|0|1|10|2|-2||4|2||-2|500007920, 500011315, 500011316|-2|34|2|||132|8|||1|
502233621|502255664|500465113|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|985|Green||2010-08-10|2010-08-14|2013-04-25|Child/Family: Moved|Child/Family: Moved||32.4||1|1|2|2|M|Multi-race (Hispanic & White)||16|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Construction|28208|1|1|Igniting Breakfast|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500011746|502234052|35|0|1|1|0|1|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|10|||17266|8|||1|
502193174|502187342|500465373|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|497|Green||2010-08-11|2010-08-18|2011-12-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16.3||2|2|1|1|M|Black||16||Mother|28273|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|Black||49|28277|Associate Degree|Married|Tech: Engineer||0|9|Recruitment Event|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|502193603|31|0|1|31|0|1|5|2|-2||4|1||-2|500000294|-2|0|4|||7443|2|||1|
502193174|503100143|500677433|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|910|Green||2013-01-25|2013-01-31|2015-07-30|Volunteer: Moved|Volunteer: Moved||29.9||2|2|1|1|M|Black||16||Mother|28273|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|White||32|28273|Bachelors Degree|Single|Business: Mgt, Admin|28217|3|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|502193603|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
500566159|500966678|500230690|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1510|Yellow||2007-12-13|2008-01-23|2012-03-12|Volunteer: Time constraint|Volunteer: Time constraint||49.6||2|2|1|1|F|Black||16||Mother|28269|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Enrollment|F|White||35|28207|||Business: Clerical||3|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500012459|500565754|31|0|2|1|0|2|5|2|-2||4|2||-2||-2|34|2|||46|2|||1|
502876870|502818822|500599930|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|331|Yellow||2012-02-23|2012-03-06|2013-01-31|Volunteer: Time constraint|Volunteer: Time constraint||10.9||2|2|1|1|F|Black||16|No|GrandMother|28206|Grandparents|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|White||30|28205|Associate Degree|Single|Business: Mgt, Admin|28204|0|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502878273|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502876870|503104166|500684838|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1241|Red||2013-02-27|2013-03-05|2016-07-28|Volunteer: Changed workplace/school partnership|Volunteer: Changed workplace/school partnership||40.8||2|2|1|1|F|Black||16|No|GrandMother|28206|Grandparents|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Multi-race (Asian & White)||28|60654|Bachelors Degree|Single|Business: Mgt, Admin|60601|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502878273|31|0|2|37|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503484186|503355490|500706097|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|925|Red||2013-08-07|2013-08-26|2016-03-08|Child: Lost interest|Child: Lost interest||30.4||1|1|1|1|M|White||16|No|Mother|28273|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||63|28226|Masters Degree|Widowed|Business: Marketing||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503486052|1|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7671|13|1561|2|1|
501434147|501926474|500441566|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2542|Green||2010-03-16|2010-03-31|NaT||||83.5||1|1|1|1|M|Black||16|No|Mother|28212|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||26|28215|||Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|501434432|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501721527|501724420|500371546|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|135|Yellow||2009-06-29|2009-07-01|2009-11-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||4.4||1|1|1|1|M|White||16|No|Mother|28211|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||47|28270|Bachelors Degree|Married|Business: Marketing|28277|2|5|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500001281|501721867|1|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502850780|502835253|500604783|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|385|Red||2012-03-19|2012-04-06|2013-04-26|Child/Family: Moved|Child/Family: Moved||12.6||1|1|1|1|M|Black||16|No|Mother|28105|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community||Match Support|M|White||54|28173|Some College|Married|Unemployed||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|502852142|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501744683|501863268|500405317|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1118|Green||2009-11-03|2009-11-06|2012-11-28|Child/Family: Moved|Child/Family: Moved||36.7||1|1|1|1|M|Black||16|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||56|28270|Some College|Separated|Unknown|28277|7|7|BBBS National Site|Web Link|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500013781|501745023|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501721760|501755476|500368545|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2689|Green||2009-06-11|2009-06-22|2016-11-01|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||88.3||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||59|28269|Masters Degree|Married|Clergy||0|0|Coca Cola|Workplace Partner|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020752|501722098|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||9610|3|||1|
502591898|503002003|500620503|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1702|Green||2012-06-20|2012-07-18|NaT||||55.9||2|2|1|1|F|Black||16|No|Mother|28214|Two Parent|$40,000 to $44,999|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||29|28210|Masters Degree|Single|Medical: Healthcare Worker||1|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502592415|31|0|2|31|0|2|10|2|-2||2|1|500004640, 500005291|-2||-2|0|4|||7496|10|||1|
502591898|502476195|500539115|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|355|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-05-31|2011-06-04|2012-05-24|Volunteer: Moved|Volunteer: Moved||11.7||2|2|1|1|F|Black||16|No|Mother|28214|Two Parent|$40,000 to $44,999|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||28|28202|Bachelors Degree|Single|Finance: Banking|28210|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502592415|31|0|2|1|0|2|10|2|500004641||4|2|500004640, 500005291|-2||-2|0|4|||7496|10|||1|500004640, 500005291
502861536|502876160|500595490|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|282|Red||2012-02-01|2012-02-08|2012-11-16|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||9.3||1|1|1|1|F|Black||16|No|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||31|28213|Bachelors Degree|Single|Insurance|28262|3|0|BBBS National Site|Web Link|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500011349|502862935|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||46|2|||1|
501347097|501099568|500278256|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2269|Yellow||2008-07-17|2008-07-30|2014-10-16|Volunteer: Time constraint|Volunteer: Time constraint||74.5||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||35|28078|Bachelors Degree|Single|Finance: Banking||4|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500011349|501347376|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
502787401|503122442|500692539|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1279|Green||2013-04-11|2013-04-30|2016-10-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||42||1|1|1|1|F|Black||16|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||41|28105|High School Graduate|Divorced|Business: Mgt, Admin|28207|6|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502788587|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503326540|503459688|500699638|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|420|Red||2013-06-05|2013-06-24|2014-08-18|Volunteer: Time constraint|Volunteer: Time constraint||13.8||2|2|1|1|F|Black||16|No|Mother|28215|Two Parent|$50,000 to $59,999||||No||Self|General Community||Match Support|F|Black||30|28213|Some College|Single|Child/Day Care Worker||2|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503328374|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
503326540|503852999|500776439|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|549|Green||2014-09-17|2014-09-28|2016-03-30|Volunteer: Time constraint|Volunteer: Time constraint||18||2|2|1|1|F|Black||16|No|Mother|28215|Two Parent|$50,000 to $59,999||||No||Self|General Community||Match Support|F|White||26|28202|Bachelors Degree|Single|Business||11|10|Current/Previous Big|Other Big|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500013781|503328374|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||17159|12|||1|
501212662|501252394|500269647|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1764|Red|Amachi|2008-06-03|2008-06-23|2013-04-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||58||1|1|1|1|M|Multi-Race (None of the above)||16|Yes|Mother|28211|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Multi-Race (None of the above)||34|28205|Bachelors Degree|Single|Business: Sales|28210|0|10|Self|Self|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501212937|7|0|1|7|0|1|10|2|-2||4|3|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
504004117|503929259|500783097|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|857|Green||2014-10-13|2014-11-10|NaT||||28.2||1|1|1|1|F|Black||16|No|Mother|28262|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||26|28269|Masters Degree|Single|Human Services: Social Worker|28202|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504006132|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1|
502478700|502578355|500544505|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1192|Red|2010-2012 OJJDP JJI|2011-07-05|2011-08-09|2014-11-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||39.2||1|1|1|1|M|Black||16|No|Mother|28269|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|White||34|28027|Masters Degree|Single|Business: Engineer|28262|0|0|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Enrollment|0|1|1|0|277|60|598|500000170|500013781|502881024|31|0|1|1|0|1|10|2|-2||4|3|500005291|-2|500015184|-1|0|5|||7462|13|||1|500005291
502280284|502241391|500500329|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|961|Red|Project Big|2010-11-30|2010-12-13|2013-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.6||1|1|1|1|F|Black||16|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|White||31|28205|Associate Degree|Married|Business: Human Resources||3|0|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502280719|31|0|2|1|0|2|10|2|500004641||4|3|500004640|-2|500004640|-2|0|10|||46|2|||1|500004640
503373647|503377601|500688140|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|322|Yellow||2013-03-15|2013-03-21|2014-02-06|Child/Family: Moved|Child/Family: Moved||10.6||1|1|2|2|F|Black||16|No|Mother|28213|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||30|28213|Some College|Single|Medical|28209|1|4|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500015820|503375503|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502980965|503007163|500618600|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|205|Red||2012-06-08|2012-06-18|2013-01-09|Volunteer: Time constraint|Volunteer: Time constraint||6.7||2|2|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||40|28209|Bachelors Degree|Single|Finance: Banking|28255|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502982410|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
502980965|503091130|500676334|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1512|Green||2013-01-22|2013-01-24|NaT||||49.7||2|2|1|1|F|Black||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||32|28210|High School Graduate|Single|Business: Sales|28277|0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502982410|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502980958|503008664|500620394|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1703|Green||2012-06-19|2012-07-17|NaT||||56||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Sales|28273|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502982410|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502508499|502079235|500538672|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|450|Red|Project Big, 2010-2012 OJJDP JJI|2011-05-26|2011-06-06|2012-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.8||1|1|1|1|F|Black||16|No|Mother|28216|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|White||33|28209|Bachelors Degree|Single|Consultant||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502508948|31|0|2|1|0|2|5|2|-2||4|3|500004640, 500005291|-2||-2|0|10|||7496|10|||1|500004640, 500005291
502062624|502067861|500460279|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|842|Yellow||2010-07-08|2010-08-30|2012-12-19|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||27.7||1|1|1|1|F|Black||16|No|Mother|28081|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||32|28083|Bachelors Degree|Single|Tech: Computer/Programmer|28216|1|7|LPL Financial|Workplace Partner|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502063048|31|0|2|31|0|2|5|2|-2||4|2||-2||-2|0|10|||11247|3|||1|
500847570|500848661|500174103|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1562|Green|Amachi|2007-04-26|2007-05-07|2011-08-16|Volunteer: Time constraint|Volunteer: Time constraint||51.3||2|2|1|1|F|Black||16|Yes|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||53|28216||Married|Business: Clerical||4|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500188056|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
500847570|502542379|500592215|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1877|Yellow|Amachi|2012-01-18|2012-01-25|NaT||||61.7||2|2|1|1|F|Black||16|Yes|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||52|28227|Bachelors Degree|Married|Insurance|28277|14|0|AA Task Force|Special Event|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|500188056|31|0|2|31|0|2|10|2|500003586||2|2|500000294|-2|500000294|-2|0|10|||11098|8|||1|500000294
501842678|502335257|500542227|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1453|Yellow||2011-06-21|2011-06-27|2015-06-19|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||47.7||2|2|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|White||53|28117|Bachelors Degree|Married|Real Estate: Realtor|28031|0|0|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|0|1|0|1|277|60|598|500000170|500015820|501843047|31|0|1|1|0|1|10|2|-2||4|2||-2|500000294, 500004901|-2|0|10|||7464|9|||1|
501842678|500189254|500418168|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|333|Green||2009-12-03|2010-01-31|2010-12-30|Volunteer: Time constraint|Volunteer: Time constraint||10.9||2|2|2|2|M|Black||16|No|Mother|28216|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|M|White||48|28036|Masters Degree||Education: College Professor||0|0||High School Partner|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|501843047|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||0|4|||1|
501829369|501687434|500376549|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|890|Green||2009-08-03|2009-08-03|2012-01-10|Volunteer: Time constraint|Volunteer: Time constraint||29.2|Y|1|1|1|1|M|White||16|No|Mother|28027|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||61|28025||Married|Medical: Doctor, Provider||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501829737|1|0|1|1|0|1|10|2|500003586||4|1||-2||-2|0|10|||7464|9|||1|
502979759|503234517|500682418|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1065|Yellow||2013-02-15|2013-03-12|2016-02-10|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||35||1|1|1|1|M|Black||16||Mother|28211|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||29|28211|Bachelors Degree||Construction|28208|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502981210|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
500826603|501004437|500548053|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|447|Red||2011-07-29|2011-08-19|2012-11-08|Volunteer: Time constraint|Volunteer: Time constraint||14.7||3|3|2|2|F|Black||16|No|Mother|28226|Two Parent|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|F|Black||39|28105|Masters Degree|Single|Business: Mgt, Admin|28204|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|500826861|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|5|||46|2|||1|
500826603|502672644|500703783|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|554|Yellow||2013-07-16|2013-08-06|2015-02-11|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.2||3|3|2|2|F|Black||16|No|Mother|28226|Two Parent|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|F|Black||34|28215|Some College|Single|Finance: Banking|28270|1|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500011349|500826861|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|5|||7464|9|||1|
500826603|500864336|500177485|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1160|Red||2007-05-17|2007-05-25|2010-07-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||38.1||3|3|1|1|F|Black||16|No|Mother|28226|Two Parent|Less than $10,000|||Y|No||Therapist/Counselor|General Community||Match Support|F|White||34|28209|||Business: Clerical||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500826861|31|0|2|1|0|2|10|2|||4|3||-2||-2|0|5|||46|2|||1|
502489575|502432606|500541789|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|426|Red|Project Big, 2010-2012 OJJDP JJI|2011-06-16|2011-06-30|2012-08-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||14||1|1|2|2|M|Black||16|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes|TV|Media|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||44|28105|Masters Degree|Married|Business: Mgt, Admin|28202|3|6|Ally Financial|Workplace Partner|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500011746|502490022|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2||-1|56|1|||12831|3|1209, 635|1|1|500004640, 500005291
500850852|500834909|500172076|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1238|Green||2007-04-13|2007-04-19|2010-09-08|Child/Family: Moved|Child/Family: Moved||40.7||1|1|1|1|M|White||16|No|Mother|28105|One Parent: Female|$60,000 to $74,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||35|28277|||Finance: Banking||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500010765|500851121|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
503238896|503004093|500678152|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|399|Red||2013-01-29|2013-01-31|2014-03-06|Volunteer: Time constraint|Volunteer: Time constraint||13.1||1|1|1|1|F|Black||16|No|Mother|28278|One Parent: Female|Less than $10,000|Yes: Active|No|Y|Yes||Self|General Community||Enrollment|F|Black||27|28212|Bachelors Degree|Single|Finance: Banking||0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|503239061|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502552438|502549491|500538826|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2093|Green|Project Big, 2010-2012 OJJDP JJI|2011-05-27|2011-06-02|2017-02-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||68.8||1|1|1|1|M|Black||16|No|GrandMother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||36|28205|Masters Degree|Living w/ Significant Other|Journalist/Media|28202|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502552891|31|0|1|1|0|1|10|2|-2||4|1|500004640, 500005291|-2||-2|0|10|||7464|9|||1|500004640, 500005291
502613782|502719849|500568690|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|665|Red||2011-10-21|2011-11-17|2013-09-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.8||1|1|1|1|M|Black||16|No|Mother|28208|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28202|Bachelors Degree|Single|Consultant||12|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502614394|31|0|1|1|0|1|5|2|-2||4|3|500005291|-2||-2|0|10|||46|2|||1|
502637589|502619035|500545174|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1056|Green|2010-2012 OJJDP JJI|2011-07-12|2011-07-19|2014-06-09|Volunteer: Moved|Volunteer: Moved||34.7||1|1|1|1|F|Black||16|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|F|White||30|28203|Masters Degree|Single|Business: Marketing|28203|0|10|Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|502638284|31|0|2|1|0|2|5|2|-2||4|1|500005291|-2||-2|6854|8|||131|1|||1|500005291
503746685|503961087|500790718|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|620|Red|PERL 2014-2016|2014-10-31|2014-11-17|2016-07-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.4||1|1|1|1|F|Black||16|No|Mother|28277|One Parent: Female|$40,000 to $44,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||31|28209|Juris Doctorate (JD)|Single|Law|28210|1|1|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503755760|31|0|2|1|0|2|10|2|-2||4|3|500014681|-2|500014681|-2|34|2|||17159|12|||1|500014681
500961270|501079472|500230999|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|391|Green||2007-12-13|2007-12-18|2009-01-12|Volunteer: Moved|Volunteer: Moved||12.8||1|1|1|1|M|Black||16|No|Mother|28215|One Parent: Female|$35,000 to $39,999||||No||BBBS Board/Staff|General Community||RTBM|M|White||46|28173|Bachelors Degree|Married|Business: Mgt, Admin||2|0|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500961540|31|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|13|||7447|3|||1|
500765381|501579025|500342803|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2427|Green||2009-02-19|2009-02-26|2015-10-20|Volunteer: Moved|Volunteer: Moved||79.7||1|1|1|1|M|Black||16|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||33|10019|Bachelors Degree|Single|Business: Marketing|28202|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|500739190|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502828137|502446364|500607445|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1155|Green||2012-04-01|2012-04-30|2015-06-29|Child/Family: Moved|Child/Family: Moved||37.9||1|1|1|1|F|Multi-Race (None of the above)||16|No|Father|28214|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher|28078|0|8|Self|Self|Big|General Community|Project Big|Match Support|0|1|0|1|277|60|598|500000170|500008321|502829415|7|0|2|31|0|2|10|2|-2||4|1||-2|500004640|-2|0|10|||7464|9|||1|
502157842|502204211|500462416|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|447|Green||2010-07-23|2010-07-23|2011-10-13|Volunteer: Time constraint|Volunteer: Time constraint||14.7||1|1|2|2|F|Black||16|No|Mother|28205|One Parent: Female|$15,000 to $19,999||||Yes||Relative|General Community||Enrollment|F|Black||41|28213|Bachelors Degree|Single|Finance: Banking|28288|12|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011639|502158281|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
503010214|503306996|500683223|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|98|Yellow||2013-02-20|2013-03-13|2013-06-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||3.2||1|1|1|1|M|Black||16|No|Mother|28226|One Parent: Female|$45,000 to $49,999||||No||Self|General Community||Match Support|M|White||36|29708|Bachelors Degree|Married|Business: Sales|28216|10|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|503011744|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
502402515|502537081|500535130|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1686|Green|2010-2012 OJJDP JJI|2011-05-05|2011-05-17|2015-12-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||55.4||1|1|1|1|M|Black||16|No|Mother|28215|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||56|28215||Single|Law: Police Officer||14|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502402953|31|0|1|31|0|1|10|2|-2||4|1|500005291|-2||-2|34|2|||7464|9|||1|500005291
502244776|502143351|500511171|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2248|Green|2010-2012 OJJDP JJI|2011-01-14|2011-01-19|NaT||||73.9||1|1|2|2|F|Black||16|No|Mother|28216|Two Parent|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||31|28209|Bachelors Degree|Single|Law|28273|5|0|Relative|Relative|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500021785|502245202|31|0|2|1|0|2|10|2|-2||2|1|500005291|-2|500000294|-2|0|4|||17161|11|||1|500005291
502874168|503456011|500696583|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|292|Green||2013-05-13|2013-05-30|2014-03-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||9.6||2|2|1|1|F|Black||16|No|Mother|28217|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||31|28203|Bachelors Degree|Single|Business: Sales|28204|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502875571|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1|
502830103|502819928|500592797|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|121|Red||2012-01-20|2012-01-31|2012-05-31|Volunteer: Moved|Volunteer: Moved||4||1|1|1|1|F|Hispanic||16|No|Mother|28213|One Parent: Female|Less than $10,000||||Yes||Self|General Community|Amachi|RTBM|F|White||28|28205|Bachelors Degree|Single|Retail: Mgt|28056|0|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502831393|3|0|2|1|0|2|7|2|-2||4|3|500000294|-2||-2|0|10|||7464|9|||1|
503606415|503665457|500736909|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1149|Green||2013-12-05|2014-01-06|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||37.7||1|1|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||32|28270|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503608292|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
501574315|501567524|500338128|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|916|Green|Amachi|2009-02-03|2009-02-11|2011-08-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||30.1||1|1|1|1|M|Black||15|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Relative|General Community|Amachi|Enrollment|M|White||33|28269|Bachelors Degree|Single|Finance: Banking|28202|4|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500003657|501574611|31|0|1|1|0|1|5|2|500003586||4|1|500000294|-2|500000294|-2|0|3|||7464|9|||1|500000294
500947380|501390454|500299095|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|338|Green|Amachi|2008-10-14|2008-11-25|2009-10-29|Child/Family: Moved|Child/Family: Moved||11.1||1|1|1|1|M|Black||15|Yes|Foster Parent|28025|Foster Home|Unknown||||No||Self|General Community|Amachi|Match Support|M|Black||50|28027|Associate Degree|Married|Firefighter|28026|0|0|Other|BBBS Board/Staff|Big|General Community|Amachi|Enrollment|1|0|1|0|277|60|598|500000170|500001262|500947650|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7671|13|||1|500000294
503503500|503390470|500706999|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1240|Green||2013-08-16|2013-08-26|2017-01-17|Volunteer: Moved|Volunteer: Moved||40.7||1|1|1|1|F|Black||15|No|Mother|28216|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||37|28078|Bachelors Degree|Single|Medical|46285|6|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503505371|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501725168|501824761|500381463|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1570|Green||2009-08-28|2009-08-31|2013-12-18|Volunteer: Moved|Volunteer: Moved||51.6||2|2|1|1|F|Multi-Race (None of the above)||15|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||34|28269|Bachelors Degree|Married|Human Services: Non-Profit||2|6|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|501724831|7|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
501725168|503828482|500767445|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|972|Green||2014-06-23|2014-07-18|NaT||||31.9||2|2|1|1|F|Multi-Race (None of the above)||15|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||32|28209|Bachelors Degree|Single|Business: Sales|45236|0|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|501724831|7|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502530227|502531485|500532078|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1265|Red|2010-2012 OJJDP JJI|2011-04-20|2011-05-04|2014-10-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||41.6||1|1|1|1|F|Hispanic||15|No|Mother|28213|One Parent: Female|$10,000 to $14,999||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||30|28210|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502530676|3|0|2|3|0|2|10|2|-2||4|3|500005291|-2||-2|0|4|||7464|9|||1|500005291
503318447|503537303|500709889|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1245|Green||2013-09-10|2013-09-27|2017-02-23|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||40.9||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||47|28215|Bachelors Degree|Married|Finance: Banking|28269|13|6|Recruitment Event|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503320281|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7458|9|||1|
501853848|501839466|500405366|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1733|Red|Amachi|2009-11-03|2009-11-30|2014-08-29|Volunteer: Time constraint|Volunteer: Time constraint||56.9||1|1|1|1|M|Black||15|Yes|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|M|Black||33|28273|||Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|501854219|31|0|1|31|0|1|5|2|-2||4|3|500000294|-2||-2|0|10|||7464|9|||1|500000294
500861521|500922138|500186899|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|796|Red||2007-08-02|2007-08-16|2009-10-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||26.2||2|2|1|1|F|Black||15|No|Mother|28208|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Enrollment|F|White||34|28202|Masters Degree|Single|Finance: Accountant|28202|0|9|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500861790|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
504031334|503882331|500787330|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|869|Green||2014-10-23|2014-10-29|NaT||||28.6||1|1|1|1|F|Black||15|No|Mother|28262|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||37|28208|Bachelors Degree|Single|Tech: Research/Design|28202|3|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503917391|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|
501674139|501664714|500363753|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|306|Green|Amachi|2009-05-14|2009-06-03|2010-04-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.1||1|1|2|2|M|Black||15|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Black||44|28273|||Finance: Accountant||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|501674477|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501833026|502451325|500518305|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2039|Yellow|2010-2012 OJJDP JJI|2011-02-17|2011-03-02|2016-09-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||67||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||41|28205|Masters Degree|Single|Education: Teacher|2122|1|5|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|501833394|31|0|2|1|0|2|10|2|-2||4|2|500005291|-2|500000294|-2|0|10|||7464|9|||1|500005291
502307403|502523838|500538762|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|395|Red|Project Big, 2010-2012 OJJDP JJI|2011-05-26|2011-05-31|2012-06-29|Volunteer: Moved|Volunteer: Moved||13||2|2|1|1|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|White||31|28203|Masters Degree|Single|Finance|28203|0|8|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502307835|31|0|1|1|0|1|10|2|-2||4|3|500004640, 500005291|-2|500004640|-2|0|4|||7464|9|||1|500004640, 500005291
502307403|502312010|500487319|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|78|Green|Project Big|2010-10-28|2010-11-30|2011-02-16|Volunteer: Moved|Volunteer: Moved||2.6||2|2|1|1|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|M|Asian||28|28202|Bachelors Degree|Single|Finance|28202|0|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502307835|31|0|1|4|0|1|10|2|500004641||4|1|500004640, 500005291|-2||-2|0|4|||7462|13|||1|500004640
500796261|503790153|500767163|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|990|Green||2014-06-19|2014-06-30|NaT||||32.5||4|4|1|1|M|White||15|No|Mother|28031|One Parent: Female|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||59|28031|Bachelors Degree|Separated|Business: Mgt, Admin|28206|20|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|500796529|1|0|1|1|0|1|10|2|-2||2|1|500005291|-2||-2|34|2|||7496|10|||1|
500796261|501180716|500277571|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|805|Green||2008-07-14|2008-08-22|2010-11-05|Volunteer: Moved|Volunteer: Moved||26.4||4|4|1|1|M|White||15|No|Mother|28031|One Parent: Female|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||45|28078|Bachelors Degree|Divorced|Tech: Engineer|28117|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|500796529|1|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|34|2|||46|2|||1|
500796261|502492476|500523882|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|688|Green|2010-2012 OJJDP JJI|2011-03-08|2011-03-15|2013-01-31|Volunteer: Time constraint|Volunteer: Time constraint||22.6||4|4|1|1|M|White||15|No|Mother|28031|One Parent: Female|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|White||36|28078|Bachelors Degree|Single|Real Estate: Realtor|28269|0|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|500796529|1|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|34|2|||7464|9|||1|500005291
501194563|501486345|500357443|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1101|Green||2009-04-15|2009-04-21|2012-04-26|Volunteer: Time constraint|Volunteer: Time constraint||36.2||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$40,000 to $44,999||||Yes||Self|General Community||Match Support|M|White||37|28269|Masters Degree|Single|Tech: Management|28262|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501194837|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501194563|503477116|500700141|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1365|Green||2013-06-10|2013-06-20|NaT||||44.8||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$40,000 to $44,999||||Yes||Self|General Community||Match Support|M|Black||30|28205|Bachelors Degree|Single|Self-Employed, Entrepreneur|28206|5|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|501194837|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
500886374|500899924|500186914|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|878|Red||2007-08-02|2007-08-14|2010-01-08|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.8||1|1|1|1|F|Black||15|No|Mother|28216|One Parent: Female|Less than $10,000|||Y|No||Self|General Community||Enrollment|F|White||35|28202|Bachelors Degree|Single|Business: Sales||0|1|Coworker|Workplace Partner|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500886644|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|10|||7447|3|||1|
501543766|501422869|500383624|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|392|Red||2009-09-09|2009-09-29|2010-10-26|Volunteer: Moved|Volunteer: Moved||12.9||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||39|28078|Masters Degree|Single|Business: Mgt, Admin|28115|1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501544058|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
500560343|500464026|500138747|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|820|Green||2006-11-08|2006-11-08|2009-02-05|Vol: Other Reason|Vol: Other Reason||26.9||1|1|2|2|F|Black||15||GrandMother|28025|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||64|28027||Married|Business: Sales||0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500560595|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
503005868|502935610|500623124|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1678|Red||2012-07-06|2012-07-24|2017-02-26|Child: Lost interest|Child: Lost interest||55.1||1|1|1|1|M|Multi-race (Black & Hispanic)||15||Mother|28270|One Parent: Female|$25,000 to $29,999|||Y|No||Therapist/Counselor|General Community||Match Support|M|White||51|28173|Bachelors Degree|Married|Consultant|28173|1|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503007379|38|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|5|||7671|13|||1|
500496598|501383928|500299090|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3066|Yellow|Amachi, Cabarrus County|2008-10-14|2008-10-23|NaT||||100.7||2|2|1|1|M|White||15|Yes|Mother|28083|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community|Amachi, Cabarrus County|Match Support|M|White||35|28083|Masters Degree|Single|Business: Mgt, Admin|28027|2|3|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|500496849|1|0|1|1|0|1|10|2|500003586||2|2|500000294, 500016374|-2|500016374|-2|34|2|||7464|9|||1|500000294, 500016374
502548212|502469646|500531329|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|600|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-04-14|2011-04-29|2012-12-19|Volunteer: Moved|Volunteer: Moved||19.7||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||28|28210|Bachelors Degree|Single|Business: Marketing||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502548665|31|0|2|31|0|2|5|2|500004641||4|2|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291
500474841|500370830|500133665|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1886|Yellow||2006-10-26|2006-11-18|2012-01-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||62||1|1|2|2|F|Black||15||Mother|28208|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|Multi-Race (None of the above)||52|28227|Bachelors Degree|Single|Education: Admin||4|0|BBBS National Site|Web Link|Big|General Community||Enrollment|1|0|1|0|277|60|598|500000170|500013709|500474737|31|0|2|7|0|2|10|2|-2||4|2||-2||-2|34|2|||46|2|||1|
501177069|501613868|500361364|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|41|Green||2009-05-05|2009-05-13|2009-06-23|Child/Family: Infraction of match rules/agency policies Vol: Does Not Like Child or Parent|Child/Family: Infraction of match rules/agency policies|Vol: Does Not Like Child or Parent|1.3||2|2|2|2|M|Black||15|No|Mother|28210|One Parent: Female|$10,000 to $14,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||51|28278||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501177343|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
501177069|501385945|500326033|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|113|Green||2008-12-12|2009-01-12|2009-05-05|Vol: Other Reason|Vol: Other Reason||3.7||2|2|1|1|M|Black||15|No|Mother|28210|One Parent: Female|$10,000 to $14,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28209||Single|Medical: Doctor, Provider||0|1|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501177343|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7671|13|||1|
501201381|501248988|500318903|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|323|Green||2008-11-21|2008-12-08|2009-10-27|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||10.6||1|1|1|1|F|Hispanic||15|No|Aunt|28212|Two Parent|Unknown||||Yes||Service Organization|General Community||Match Support|F|White||39|28205||Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|501201651|3|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|11|||7464|9|||1|
502606280|501177078|500546219|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|168|Green|2010-2012 OJJDP JJI|2011-07-14|2011-07-21|2012-01-05|Child/Family: Time constraints|Child/Family: Time constraints||5.5||1|1|1|1|F|White||15|No|Mother|28081|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|2010-2012 OJJDP JJI|RTBM|F|White||45|28078|Bachelors Degree|Married|Business: Human Resources||2|0|BBBS National Site|Web Link|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500002335|502606797|1|0|2|1|0|2|7|2|-2||4|1|500005291|-2||-2|0|4|||46|2|||1|500005291
502838696|502445477|500582889|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|119|Red||2011-11-30|2011-11-30|2012-03-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.9||1|1|1|1|F|Hispanic||15|No|Mother|28031|Two Parent|Unknown||||Yes||School|General Community||Match Support|F|White||51|28031|Some College|Married|Real Estate: Realtor|28031|5|0||Relative|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500011746|502839988|3|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||0|11|||1|
503532788|503939365|500772617|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|936|Green|Cabarrus County|2014-08-18|2014-08-23|NaT||||30.8||1|1|1|1|F|Black||15|Yes|GrandMother|28075|Grandparents|$10,000 to $14,999|||Y|Yes||Relative|General Community|Amachi, Cabarrus County|Match Support|F|Black||33|28269|PHD|Single|Education: Admin|28081|4|0|Current/Previous Big|Other Big|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|503534663|31|0|2|31|0|2|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|3|||17159|12|||1|500016374
503346838|503369070|500693781|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|163|Yellow||2013-04-19|2013-05-29|2013-11-08|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||5.4||1|1|1|1|M|Black||15|Yes|Mother|28213|One Parent: Female|$50,000 to $59,999|||Y|No|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||49|28078|Masters Degree|Divorced|Finance||0|3|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500004169|503348683|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2||-2|34|2|||7464|9|||1|
502990571|503004889|500619186|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|330|Yellow||2012-06-13|2012-06-25|2013-05-21|Volunteer: Time constraint|Volunteer: Time constraint||10.8||2|2|1|1|F|Multi-race (Black & Hispanic)||15|Yes|Mother|28217|Two Parent|$35,000 to $39,999||||Yes||Self|General Community||Match Support|F|Black||29|28217|Bachelors Degree|Single|Business||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502992028|38|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502990571|503400909|500707095|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1077|Red||2013-08-19|2013-08-30|2016-08-11|Child/Family: Moved|Child/Family: Moved||35.4||2|2|1|1|F|Multi-race (Black & Hispanic)||15|Yes|Mother|28217|Two Parent|$35,000 to $39,999||||Yes||Self|General Community||Match Support|F|Black||28|28269|Bachelors Degree|Single|Business||0|7|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502992028|38|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502317500|502658498|500587614|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1269|Red|Project Big, Project Big AND Amachi|2011-12-16|2012-02-08|2015-07-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||41.7||1|1|2|2|M|Black||15|No|Mother|28214|One Parent: Female|Unknown||||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|M|White||33|28214|Associate Degree|Single|Law: Security Officer|28208|2|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502317931|31|0|1|1|0|1|10|2|-2||4|3|500004640, 500004901|-2||-2|0|4|||7464|9|||1|500004640, 500004901
501224282|501389463|500296679|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1337|Red|Amachi|2008-10-08|2008-10-16|2012-06-14|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||43.9||2|2|1|1|F|Black||15|Yes|Mother|28270|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||35|28215|Bachelors Degree|Single|Finance: Banking|28262|2|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500013781|501224558|31|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|5635|9|||7453|7|||1|500000294
501224282|503347558|500700583|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1365|Green|Amachi|2013-06-13|2013-06-20|NaT||||44.8||2|2|1|1|F|Black||15|Yes|Mother|28270|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||35|28205|Bachelors Degree|Married|Business: Mgt, Admin|28217|5|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|501224558|31|0|2|1|0|2|10|2|-2||2|1|500000294|-2||-2|5635|9|||46|2|||1|500000294
501015998|501322799|500292474|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|111|Green|Amachi|2008-09-29|2008-10-28|2009-02-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.6||1|1|1|1|M|Black||15|Yes|Mother|28212|One Parent: Female|Less than $10,000||||Yes||Self|General Community|Amachi|RTBM|M|Black||36|28226|Some College|Single|Business: Clerical||1|2|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500007521|501016267|31|0|1|31|0|1|7|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7462|13|||1|500000294
500545470|500815012|500173957|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3192|Red|Amachi|2007-04-26|2007-04-30|2016-01-25|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||104.9||1|1|1|1|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown||||No||Relative|General Community|Amachi|Match Support|M|White||34|29708|Bachelors Degree|Single|Self-Employed, Entrepreneur|29708|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|501750989|31|0|1|1|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|3|||2238|7|||1|500000294
503834613|503790527|500770182|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|219|Yellow||2014-07-22|2014-07-29|2015-03-05|Volunteer: Time constraint|Volunteer: Time constraint||7.2||1|1|1|1|M|White||15|No|Mother|28226|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||RTBM|M|White||73|28277|High School Graduate|Married|Arts, Entertainment, Sports||0|0|Radio|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|503836592|1|0|1|1|0|1|7|2|-2||4|2||-2||-2|0|10|||131|1|||1|
502763567|502672644|500587190|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|292|Red|Project Big|2011-12-15|2011-12-30|2012-10-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||9.6||1|1|2|2|F|Black||15|No|Mother|28211|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||34|28215|Some College|Single|Finance: Banking|28270|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502764479|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|500004640
502597596|502560341|500540008|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|286|Green|Project Big, 2010-2012 OJJDP JJI|2011-06-06|2011-06-30|2012-04-11|Child/Family: Moved|Child/Family: Moved||9.4||1|1|1|1|F|Black||15||Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||33|28273|Bachelors Degree|Single|Medical|28277|2|9|Self|Self|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500013709|502598113|31|0|2|31|0|2|10|2|-2||4|1|500004640, 500005291|-2||-1|0|4|||7464|9|||1|500004640, 500005291
502875276|502877270|500594084|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|486|Yellow||2012-01-26|2012-02-06|2013-06-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Enrollment|M|White||30|28031|Bachelors Degree|Single|Finance|28027|1|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502876679|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
502668768|502571563|500552927|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|423|Yellow||2011-09-01|2011-09-17|2012-11-13|Volunteer: Time constraint|Volunteer: Time constraint||13.9||1|1|1|1|F|Hispanic||15|No|Mother|28212|One Parent: Female|$10,000 to $14,999||||Yes||School|General Community||Match Support|F|Hispanic||30|28226|Bachelors Degree|Married|Law: Paralegal|28226|4|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502669595|3|0|2|3|0|2|10|2|-2||4|2||-2||-2|0|4|||7462|13|||1|
503533022|503534544|500718872|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|495|Green||2013-10-14|2013-10-24|2015-03-03|Volunteer: Moved|Volunteer: Moved||16.3||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||RTBM|M|Black||27|28216|Bachelors Degree|Single|Business: Engineer|28202|0|1|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|503534897|31|0|1|31|0|1|7|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
502378719|502454212|500518127|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|491|Green|2010-2012 OJJDP JJI|2011-02-16|2011-02-24|2012-06-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||16.1||1|1|1|1|F|Black||15|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|RTBM|F|White||30|28202|Bachelors Degree|Single|Business: Marketing||1|0|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500001281|502379157|31|0|2|1|0|2|7|2|-2||4|1|500005291|-2|500000294, 500004640|-2|0|10|||46|2|||1|500005291
501034365|501580873|500370326|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|583|Green|Amachi|2009-06-22|2009-07-06|2011-02-09|Volunteer: Health|Volunteer: Health||19.2||2|2|1|1|M|Black||15|Yes|Mother|28216|One Parent: Female|$30,000 to $34,999||||No|BBBS National Site|Web Link|General Community|Amachi|Enrollment|M|Black||52|28262|Associate Degree|Married|Finance: Banking||7|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501034638|31|0|1|31|0|1|5|2|-2||4|1|500000294|-2|500000294|-2|34|2|||7453|7|||1|500000294
502859187|503090888|500658723|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1573|Green|VOL - PreMatch|2012-11-12|2012-11-24|NaT||||51.7||2|2|1|1|F|Black||15|No|GrandMother|28205|Grandparents|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||31|28209|Associate Degree|Married|Retail: Mgt|28134|4|3|UNCC|College Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|500187987|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||9221|5|||1|500007920
502859187|502849360|500597086|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|78|Red||2012-02-08|2012-03-14|2012-05-31|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||2.6||2|2|2|2|F|Black||15|No|GrandMother|28205|Grandparents|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||28|28213|Bachelors Degree|Single|Medical: Nurse||0|4|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|500187987|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502030263|501923553|500438867|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2542|Green||2010-03-03|2010-03-31|NaT||||83.5||1|1|1|1|M|White||15|No|Mother|29710|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Community||Match Support|M|White||38|28210|||Business||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502030662|1|0|1|1|0|1|10|2|-2||2|1||-2||-2|6855|8|||7464|9|||1|
501247269|501914025|500515263|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2215|Green|2010-2012 OJJDP JJI, Cabarrus County|2011-02-03|2011-02-21|NaT||||72.8||2|2|1|1|F|White||15|No|Father|28025|One Parent: Male|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|White||43|28027|Associate Degree|Married|Student: College||4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|500341682|1|0|2|1|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7496|10|||1|500005291, 500016374
501247269|501444307|500339623|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|331|Green||2009-02-09|2009-02-17|2010-01-14|Volunteer: Time constraint|Volunteer: Time constraint||10.9||2|2|1|1|F|White||15|No|Father|28025|One Parent: Male|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|White||33|28083|Bachelors Degree|Married|Student: College|28233|0|3|Recruitment Event|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|500341682|1|0|2|1|0|2|10|2|-2||4|1|500016374|-2||-2|0|10|||7458|9|||1|
501536365|501443152|500336020|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1990|Red|Amachi|2009-01-27|2009-02-03|2014-07-17|Volunteer: Time constraint|Volunteer: Time constraint||65.4||1|1|1|1|M|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|M|Black||57|28105|Some College|Married|Retail: Sales|28105|10|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|501536657|31|0|1|31|0|1|5|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||7453|7|||1|500000294
501691220|501721806|500367645|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1154|Green||2009-06-05|2009-07-02|2012-08-29|Child/Family: Moved|Child/Family: Moved||37.9||1|1|2|3|M|White||15|No|Mother|27949|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree||Business: Marketing|28031|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501691558|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502809446|502909383|500608444|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1530|Yellow|Amachi|2012-04-05|2012-04-12|2016-06-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||50.3||1|1|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Multi-race (Black & White)||33|28269|Bachelors Degree|Single|Business: Mgt, Admin||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502810724|31|0|2|36|0|2|10|2|500003586||4|2|500000294|-2||-2|0|10|||7462|13|||1|500000294
500570756|502889143|500703847|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1333|Green||2013-07-17|2013-07-22|NaT||||43.8||4|5|2|2|F|Black||15||Aunt|28213|Two Parent|Unknown||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Black||24|28262|Some College|Single|Student: College|28216|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|500214349|31|0|2|31|0|2|10|2|-2||2|1|500004640, 500005291|-2||-2|0|4|||7464|9|||1|
502551047|503347969|500681888|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|209|Green||2013-02-13|2013-02-21|2013-09-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.9||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Enrollment|M|White||28|28262|Some College|Single|Military|27260|6|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502551498|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
501190199|500839927|500408132|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|91|Green||2009-11-09|2009-12-04|2010-03-05|Volunteer: Time constraint|Volunteer: Time constraint||3||2|2|2|2|F|Black||15|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|F|White||32|28075|Bachelors Degree||Child/Day Care Worker|28075|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501190473|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501190199|501093278|500244944|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|470|Green||2008-02-13|2008-03-04|2009-06-17|Match Successful: Support No Longer Needed|Match Successful: Support No Longer Needed||15.4||2|2|1|1|F|Black||15|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|F|Black||31|28027|Some College|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|501190473|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502247579|502681447|500575685|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1621|Green|Amachi, Project Big, Project Big AND Amachi|2011-11-08|2011-12-02|2016-05-10|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||53.3||2|2|1|1|F|Black||15|Yes|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||47|28226|Bachelors Degree|Single|Education: Teacher||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502248010|31|0|2|31|0|2|10|2|500003586||4|1|500000294, 500004640, 500004901|-2||-2|0|10|||2238|7|||1|500000294, 500004640, 500004901
502247579|502322424|500483853|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|360|Yellow|Amachi, Project Big, Project Big AND Amachi|2010-10-21|2010-10-30|2011-10-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.8||2|2|1|1|F|Black||15|Yes|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||29|28203||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502248010|31|0|2|1|0|2|10|2|500004772||4|2|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7496|10|||1|500000294, 500004640, 500004901
502051702|503378835|500690864|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1430|Yellow|Amachi|2013-04-01|2013-04-16|NaT||||47||1|1|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||31|28262|Bachelors Degree|Single|Finance|28281|5|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501977740|31|0|2|31|0|2|10|2|-2||2|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
501865540|501645618|500425153|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|280|Red||2010-01-07|2010-01-19|2010-10-26|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||9.2||1|1|1|1|F|White||15||Relative: Other|28208|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||49|28273|||Business: Human Resources|28036|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501865913|1|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501253195|500395148|500282924|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3065|Green|Amachi|2008-08-21|2008-10-24|NaT||||100.7||1|1|2|2|M|Black||15|Yes|Mother|28230|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||37|28203|Masters Degree|Single|Medical: Doctor, Provider|28211|6|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|501253471|31|0|1|1|0|1|10|2|500003586||2|1||-2||-2|0|10|||7464|9|||1|500000294
503569117|503583743|500735247|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|448|Green||2013-11-27|2013-12-19|2015-03-12|Child/Family: Moved|Child/Family: Moved||14.7||1|1|1|1|F|Black||15|No|Mother|2649|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||32|28203|Doctor of Medicine (MD)|Living w/ Significant Other|Medical|28112|1|2|other|College Partner|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500015820|503570990|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7670|5|||1|
502549826|503431300|500693780|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1388|Green||2013-04-19|2013-05-28|NaT||||45.6||4|4|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|Black||38|28215|Bachelors Degree|Single|Business: Mgt, Admin|28210|11|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502550279|31|0|2|31|0|2|10|2|-2||3|1|500014505, 500015184|-1||-2|0|4|||7464|9|||1|
502549826|502584664|500537198|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|625|Red|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|2011-05-20|2011-06-13|2013-02-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||20.5||4|4|1|1|F|Black||15|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|mentor2.0, mentor2.0 2015|Match Support|F|White||32|28209|Bachelors Degree|Single|Law: Paralegal|28204|1|5||Relative|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011349|502550279|31|0|2|1|0|2|10|2|500004772||4|3|500014505, 500015184|-1|500004640|-2|0|4|||0|11|||1|500000294, 500004640, 500004901, 500005291
503831166|503861120|500772203|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|523|Green||2014-08-13|2014-08-21|2016-01-26|Volunteer: Time constraint|Volunteer: Time constraint||17.2||1|1|1|1|M|Black||15|No|Mother|28227|One Parent: Female|$60,000 to $74,999||||No|AARTF|BBBS Board/Staff|General Community||Match Support|M|Black||23|28227|Some College|Single|Student: College|28078|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503833145|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|7294|13|||7496|10|||1|
502699353|503945609|500783805|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|870|Green|PERL 2014-2016|2014-10-15|2014-10-28|NaT||||28.6||2|2|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown||||No||School|General Community|PERL 2014-2016, Project Big|Match Support|F|Black||50|28278|Bachelors Degree|Single|Finance: Banking|29715|15|2|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|502700198|31|0|2|31|0|2|10|2|-2||2|1|500004640, 500014681|-2|500000294, 500014681|-2|0|4|||7496|10|||1|500014681
502699353|502530062|500568290|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|822|Yellow|Project Big|2011-10-20|2011-10-31|2014-01-30|Volunteer: Moved|Volunteer: Moved||27||2|2|1|1|F|Black||15|No|Mother|28208|One Parent: Female|Unknown||||No||School|General Community|PERL 2014-2016, Project Big|Match Support|F|White||29|28204|Bachelors Degree|Single|Business|28255|0|2|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500015820|502700198|31|0|2|1|0|2|10|2|-2||4|2|500004640, 500014681|-2|500000294|-2|0|4|||7464|9|||1|500004640
501989028|503039778|500641725|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1408|Yellow||2012-10-04|2012-10-22|2016-08-30|Child/Family: Moved|Child/Family: Moved||46.3||2|2|1|1|M|Black||15|No|Mother|28273|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28273|Juris Doctorate (JD)|Single|Law: Lawyer||0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502425720|31|0|1|31|0|1|10|2|-2||4|2|500005291|-2||-2|6855|8|||7496|10|635|1|1|
501989028|502346780|500521737|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|377|Red|2010-2012 OJJDP JJI|2011-03-04|2011-03-16|2012-03-27|Volunteer: Time constraint|Volunteer: Time constraint||12.4||2|2|1|1|M|Black||15|No|Mother|28273|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|M|Black|Other African|44|28212|Bachelors Degree|Married|Business: Marketing||12|0|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011746|502425720|31|0|1|31|31|1|10|2|-2||4|3|500005291|-2|500000294|-2|6855|8|||7671|13|||1|500005291
502972004|502908172|500617689|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|139|Red||2012-06-04|2012-06-29|2012-11-15|Volunteer: Time constraint|Volunteer: Time constraint||4.6||1|1|1|1|F|Black||15|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes|AARTF|BBBS Board/Staff|General Community||Match Support|F|Black||57|28273|Masters Degree|Single|Business|28210|5|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502973441|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|7294|13|||7462|13|||1|
503023832|503139766|500692957|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1385|Green||2013-04-15|2013-05-31|NaT||||45.5||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||33|28278|Bachelors Degree|Single|Arts, Entertainment, Sports|28269|0|4|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503025372|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1|
501730492|501595189|500367450|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|60|Green||2009-06-04|2009-06-19|2009-08-18|Volunteer: Time constraint|Volunteer: Time constraint||2||1|1|1|1|F|Black||15|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|White||33|28210|||Unknown||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501730818|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503831971|504011759|500788190|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|225|Yellow||2014-10-27|2014-11-17|2015-06-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.4||1|1|2|2|M|Black||15|Yes|Mother|28269|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|Hispanic||31|28209|High School Graduate|Single|Finance|28262|1|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|503833950|31|0|1|3|0|1|10|2|-2||4|2|500000294|-2||-2|0|10|||46|2|||1|
502255225|502312682|500487118|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2118|Red||2010-10-28|2010-11-08|2016-08-26|Volunteer: Moved|Volunteer: Moved||69.6||1|1|1|1|M|Hispanic||15||Mother|28212|One Parent: Female|Unknown||||No|Spanish Radio|Media|General Community||Match Support|M|White||33|28226|Bachelors Degree|Single|Education: Teacher||3|0|Spanish Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502255655|3|0|1|1|0|1|10|2|-2||4|3||-2||-2|7068|1|||11662|1|||1|
502845758|502944923|500606912|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1245|Red||2012-03-28|2012-04-19|2015-09-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||40.9||1|1|1|1|M|Black||15|No|Mother|28202|One Parent: Male|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||30|28277||Single|Business||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502847118|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
501811395|500876892|500436702|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2563|Green|Cabarrus County|2010-02-23|2010-03-10|NaT||||84.2||1|1|1|1|F|Black||15|No|Mother|28027|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|F|Black||60|28213||Married|Business: Clerical||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|501811730|31|0|2|31|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|6854|8|||2238|7|||1|500016374
503452081|503371848|500694854|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|529|Green||2013-04-29|2013-05-09|2014-10-20|Volunteer: Moved|Volunteer: Moved||17.4||1|1|1|1|M|White||15|No|Mother|28227|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|White||26|28269|Bachelors Degree|Single|Business: Engineer||0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503453947|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501332658|501814288|500384166|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2669|Green|Amachi|2009-09-11|2009-09-29|2017-01-19|Child: Severity of challenges|Child: Severity of challenges||87.7||1|1|1|1|M|Black||15|Yes|GrandMother|28213|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||46|28227|High School Graduate|Single|Medical: Healthcare Worker|28269|4|0|Coworker|Workplace Partner|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|0|1|277|60|598|500000170|500020752|501332937|31|0|1|1|0|1|10|2|-2||4|1|500000294|-2|500007920, 500011315, 500011316|-2|6854|8|||7447|3|||1|500000294
502495501|502508181|500531873|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2127|Green|2010-2012 OJJDP JJI|2011-04-19|2011-05-20|NaT||||69.9||1|1|1|1|M|White||15|No|Mother|28226|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||55|28210|Bachelors Degree|Married|Finance|28203|1|6|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|0|1|277|60|598|500000170|500018851|502495950|1|0|1|1|0|1|10|2|-2||2|1|500005291|-2|500005291|-2|0|10|||7464|9|||1|500005291
501810015|501646021|500391598|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|843|Green||2009-10-06|2009-10-19|2012-02-09|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||27.7||1|1|2|2|M|Hispanic||15|No|Mother|28210|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501810370|3|0|1|3|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503803718|503930530|500783205|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|854|Green||2014-10-13|2014-11-13|NaT||||28.1||1|1|1|1|M|Black||15|No|Mother|28208|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Some Other Race||33|28056|Doctor of Medicine (MD)|Single|Medical: Doctor, Provider|28204|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503805695|31|0|1|41|0|1|10|2|-2||2|1||-2||-2|34|2|||46|2|||1|
502983808|503140432|500668771|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1152|Yellow|Amachi|2012-12-11|2012-12-15|2016-02-10|Volunteer: Time constraint|Volunteer: Time constraint||37.8||1|1|1|1|M|Black||15|Yes|Mother|28205|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community|Amachi|Match Support|M|White||27|28203|Bachelors Degree|Single|Business||0|2|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|502985262|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2|500000294|-2|0|4|||7464|9|||1|500000294
503041998|503110820|500638908|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1612|Yellow||2012-09-26|2012-10-16|NaT||||53||1|1|1|1|M|Black||15|No|Mother|28214|One Parent: Female|$45,000 to $49,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||34|28207|Masters Degree|Married|Finance|28273|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503043639|31|0|1|1|0|1|10|2|-2||2|2||-2||-2|34|2|||7464|9|||1|
502146600|503483337|500760757|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1051|Green||2014-04-23|2014-04-30|NaT||||34.5||1|1|2|2|F|Black||15|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||45|28227|Bachelors Degree|Married|Customer Service|28262|18|0|Big For A Day|Special Event|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|502932575|31|0|2|31|0|2|10|2|-2||2|1||-2|500000294|-2|6854|8|||16422|8|||1|
501604446|501832854|500396125|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|215|Yellow||2009-10-16|2009-10-22|2010-05-25|Volunteer: Time constraint|Volunteer: Time constraint||7.1||2|2|2|2|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||65|28213|Bachelors Degree|Married|Tech: Engineer|28213|2|9|TV|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500001281|501604760|31|0|1|1|0|1|10|2|-2||4|2|500005291|-2|500000294|-2|0|10|||130|1|||1|
501604446|502664359|500555050|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2005|Green|2010-2012 OJJDP JJI|2011-09-15|2011-09-19|NaT||||65.9||2|2|1|1|M|Black||15|No|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28213|Bachelors Degree|Married|Tech: Support, Writing|28273|11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501604760|31|0|1|31|0|1|10|2|-2||2|1|500005291|-2||-2|0|10|||7462|13|||1|500005291
502093473|502256927|500468462|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|391|Green|Amachi|2010-09-01|2010-09-29|2011-10-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.8||2|2|1|1|F|Black||15|Yes|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|White||33|28203|Bachelors Degree|Single|Business: Mgt, Admin|28273|0|8|Self|Self|Big|General Community|Amachi, Project Big AND Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502093897|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294, 500004901|-2|34|2|||7464|9|||1|500000294
502093473|502080552|500447214|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|110|Green||2010-04-14|2010-04-28|2010-08-16|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.6||2|2|1|1|F|Black||15|Yes|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|White||29|28227||Married|Student: College||0|0|TV|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|502093897|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||130|1|||1|
502612404|503790988|500773744|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|233|Red|PERL 2014-2016|2014-08-28|2014-10-06|2015-05-27|Volunteer: Moved|Volunteer: Moved||7.7||2|2|1|1|F|Some Other Race||15|No|Aunt|28217|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||26|28217|Bachelors Degree|Single|Business|28277|0|8|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|500188044|41|0|2|31|0|2|10|2|-2||4|3||-2|500014681|-2|0|10|||46|2|||1|500014681
501750505|501777375|500375403|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1063|Green||2009-07-24|2009-07-31|2012-06-28|Volunteer: Moved|Volunteer: Moved||34.9||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|Black||32|28205|Bachelors Degree|Single|Finance: Banking||3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501750847|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502663937|503296990|500684232|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1478|Green||2013-02-25|2013-02-27|NaT||||48.6||1|1|1|1|M|Black||15|No|Mother|28212|Two Parent|$35,000 to $39,999|Yes: Active|Yes||No||Relative|General Community||Match Support|M|White||30|28105|Bachelors Degree|Single|Business: Sales|17001|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502664764|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|3|||7496|10|||1|
500864335|500873774|500176256|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|799|Yellow||2007-05-09|2007-05-23|2009-07-30|Volunteer: Time constraint|Volunteer: Time constraint||26.3||1|1|1|1|F|Black||15||Mother|28215|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||38|28269|Bachelors Degree|Single|Medical: Healthcare Worker||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009007|500864598|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|4|||7464|9|||1|
502980163|502949611|500626324|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|385|Red||2012-07-26|2012-08-10|2013-08-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.6||1|1|1|1|M|Black||15|No|Mother|28105|One Parent: Female|$25,000 to $29,999|||Y|No||Self|General Community||Match Support|M|Black||39|28110|Some College|Married|Business||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|502981615|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502637403|502883455|500613355|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|676|Green|Amachi|2012-05-04|2012-05-24|2014-03-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||22.2||1|1|1|1|F|Black||15|Yes|Mother|28278|One Parent: Female|$30,000 to $34,999||||No||School|General Community|Amachi|Match Support|F|White||24|28105|Some College||Student: College||0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500008321|502638098|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|4|||46|2|||1|500000294
501641325|501715652|500366872|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2231|Green||2009-06-01|2009-06-24|2015-08-03|Volunteer: Time constraint|Volunteer: Time constraint||73.3||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Multi-race (Asian & White)||34|28205|Bachelors Degree|Single|Tech: Research/Design|28255|3|1|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500011349|501641648|31|0|1|37|0|1|10|2|-2||4|1|500000294|-2|500000294|-2|6854|8|||7464|9|||1|
501627668|503921388|500773645|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|392|Red||2014-08-27|2014-09-15|2015-10-12|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12.9||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||40|28217|Masters Degree|Single|Finance: Accountant|28034|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|501627988|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||17159|12|||1|
501627668|501865457|500423715|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|962|Yellow||2009-12-23|2010-01-26|2012-09-14|Volunteer: Moved|Volunteer: Moved||31.6||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||38|28209|Bachelors Degree|Single|Business|28277|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501627988|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
502537639|502387375|500533008|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|401|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-04-23|2011-04-26|2012-05-31|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||13.2||1|1|1|1|F|Black||15|No|Mother|28208|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|White||39|28209|Bachelors Degree|Single|Finance: Banking|28202|9|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013709|502538092|31|0|2|1|0|2|5|2|-2||4|2|500004640, 500005291|-2||-2|0|4|||46|2|||1|500004640, 500005291
502270499|502376097|500501731|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|91|Green||2010-12-03|2010-12-28|2011-03-29|Volunteer: Time constraint|Volunteer: Time constraint||3||2|2|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||67|28207|Bachelors Degree|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502231230|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|5635|9|||7464|9|||1|
502270499|502510107|500536754|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2122|Green|Amachi|2011-05-18|2011-05-25|NaT||||69.7||2|2|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Match Support|F|White||34|28203|Masters Degree|Single|Business: Mgt, Admin|28273|0|7|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502231230|31|0|2|1|0|2|10|2|500003586||2|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
501010684|502570658|500549074|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|575|Red|2010-2012 OJJDP JJI|2011-08-08|2011-08-17|2013-03-14|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||18.9||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Less than $10,000||||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|White||46|28227|Bachelors Degree|Married|Business: Mgt, Admin|28277|10|0|Local Print|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|503560069|31|0|1|1|0|1|10|2|-2||4|3|500005291|-2||-2|7016|11|||7439|1|||1|500005291
501010684|503491643|500710107|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1220|Green||2013-09-10|2013-10-22|2017-02-23|Volunteer: Time constraint|Volunteer: Time constraint||40.1||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|Less than $10,000||||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|M|White||41|28269|Bachelors Degree|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503560069|31|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|7016|11|||7464|9|||1|
501123191|502153920|500478644|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1888|Green||2010-10-11|2010-10-20|2015-12-21|Child/Family: Moved|Child/Family: Moved||62||2|2|1|1|F|Black||15|No|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||48|28210|Some College|Single|Human Services||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|500915629|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501123191|500898008|500234534|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|888|Green||2007-12-21|2007-12-21|2010-05-27|Volunteer: Moved|Volunteer: Moved||29.2||2|2|1|1|F|Black||15|No|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||33|28202|Bachelors Degree|Living w/ Significant Other|Journalist/Media|28203|0|10|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500915629|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503425373|500967139|500699541|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|366|Red||2013-06-05|2013-06-24|2014-06-25|Child/Family: Moved|Child/Family: Moved||12||1|1|2|2|M|Multi-race (Black & White)||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||60|28269|Bachelors Degree|Married|Business: Sales|28079|9|0|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503427238|36|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||4748|14|||1|
502180724|502391505|500505039|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2268|Green|Amachi, Project Big, Project Big AND Amachi|2010-12-13|2010-12-30|NaT||||74.5|Y|2|2|2|2|M|Black||15|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||38|28210|Bachelors Degree|Married|Business||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|502181148|31|0|1|31|0|2|10|2|500004772||2|1|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||7438|1|||1|500000294, 500004640, 500004901
502180724|502176723|500457633|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|150|Green|Amachi|2010-06-22|2010-06-25|2010-11-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.9||2|2|1|1|M|Black||15|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|M|Hispanic||32|28269|Some College|Single|Customer Service||0|0|UnitedMethodistChrch|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|502181148|31|0|1|3|0|1|10|2|500003586||4|1|500000294, 500004640, 500004901|-2|500000294|-2|0|10|||8529|7|||1|500000294
500784687|503531111|500709609|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|826|Red||2013-09-09|2013-10-01|2016-01-05|Volunteer: Time constraint|Volunteer: Time constraint||27.1||2|2|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|No||Therapist/Counselor|General Community||Match Support|M|Black||32|28277|Bachelors Degree|Single|Construction|28211|0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|500784955|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|5|||7464|9|||1|
502287066|502501212|500532817|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1220|Green|2010-2012 OJJDP JJI|2011-04-21|2011-05-03|2014-09-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||40.1||2|2|1|1|M|Black||15||GrandMother|28227|One Parent: Female|Unknown|||Y|Yes|AARTF|BBBS Board/Staff|General Community|2010-2012 OJJDP JJI|Enrollment|M|White||37|28215|Associate Degree|Married|Medical: Nurse||3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502287498|31|0|1|1|0|1|5|2|-2||4|1|500005291|-2||-2|7294|13|||7464|9|||1|500005291
501575257|501234758|500348757|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1651|Red||2009-03-11|2009-03-18|2013-09-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||54.2||1|1|1|1|M|Black||15|No|Mother|28079|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||38|28079||Married|Law: Police Officer|28211|5|0|Recruitment Event|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500004169|501575553|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7458|9|||1|
503230648|503169561|500700323|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1338|Green||2013-06-12|2013-07-17|NaT||||44||1|1|1|1|F|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|Black||39|28214|Bachelors Degree|Single|Govt||1|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|502841119|31|0|2|31|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
501611456|501876475|500450969|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2484|Green||2010-05-03|2010-05-28|NaT||||81.6||1|1|1|1|M|Black||15|No|Mother|28262|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black|Other African|32|28262||Married|Law: Police Officer||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501611776|31|0|1|31|31|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503523387|503537943|500720846|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|388|Green||2013-10-18|2013-10-29|2014-11-21|Child/Family: Moved|Child/Family: Moved||12.7||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||29|28262|Juris Doctorate (JD)|Single|Law: Lawyer||0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|503525262|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503246887|503253208|500690197|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1141|Green|Amachi|2013-03-27|2013-04-10|2016-05-25|Volunteer: Moved|Volunteer: Moved||37.5||1|1|1|1|M|Black||15|No|Mother|28212|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||27|28209|Bachelors Degree|Single|Finance|28255|1|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|503248691|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||46|2|||1|500000294
501372080|501347529|500292730|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1111|Green||2008-09-29|2008-10-10|2011-10-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||36.5||2|2|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|M|White||39|28203|Bachelors Degree|Single|Finance: Banking|28255|2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008629|501372359|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|3|||7496|10|||1|
501372080|502500246|500640327|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1269|Yellow||2012-10-01|2012-10-31|2016-04-22|Child/Family: Moved|Child/Family: Moved||41.7||2|2|2|2|M|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Relative|General Community||Match Support|M|White||31|28269|Masters Degree|Single|Insurance|28262|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501372359|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|3|||7496|10|||1|
501809541|501620528|500375025|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2778|Green||2009-07-22|2009-08-07|NaT||||91.3||1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||49|28031|Bachelors Degree|Married|Transport: Pilot|40223|9|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501809896|36|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502415267|502657931|500550917|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|444|Red|2010-2012 OJJDP JJI|2011-08-19|2011-09-19|2012-12-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||14.6||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|$25,000 to $29,999|||Y|Yes||Therapist/Counselor|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||53|28269|Some College|Single|Unknown||0|0|Radio|Media|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500015820|502415705|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2||-2|0|5|||131|1|||1|500005291
501585465|501613868|500350872|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|4|Green||2009-03-19|2009-03-23|2009-03-27|Vol: Does Not Like Child or Parent|Vol: Does Not Like Child or Parent||0.1||1|1|2|2|M|Black||15|No|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|Black||51|28278||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501585785|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501762789|501663549|500378602|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|210|Green||2009-08-13|2009-08-13|2010-03-11|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.9||1|1|1|1|M|Black||15|No|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|White||37|28278||Single|Finance: Banking|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009242|501763124|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
501365904|501459709|500353421|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1234|Yellow||2009-03-30|2009-04-20|2012-09-05|Child/Family: Moved|Child/Family: Moved||40.5||1|1|1|1|M|Black||15|No|Mother|28269|One Parent: Female|Unknown|||Y|No||Self|General Community||Enrollment|M|Black||48|28269|Some College|Married|Business: Engineer|28262|20|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501366183|31|0|1|31|0|1|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502252828|502602451|500547383|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1532|Green|2010-2012 OJJDP JJI|2011-07-25|2011-08-03|2015-10-13|Volunteer: Time constraint|Volunteer: Time constraint||50.3||1|1|1|1|M|Black||15||GrandMother|28227|Grandparents|Unknown||||No||Self|General Community|PERL 2014-2016|RTBM|M|White||27|28205|Associate Degree|Single|Law: Police Officer||0|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|0|1|277|60|598|500000170|500017777|502253254|31|0|1|1|0|1|7|2|-2||4|1|500014681|-2|500005291|-2|0|10|||7496|10|||1|500005291
500791645|501365854|500307006|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|393|Green||2008-10-29|2008-11-17|2009-12-15|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||12.9||4|4|1|1|F|Multi-Race (None of the above)||15||Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Multi-race (Black & White)||33|28269|Bachelors Degree|Single|Business: Sales|28213|1|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500187654|7|0|2|36|0|2|10|2|-2||4|1|500005291|-2||-2|0|10|||7464|9|||1|
500791645|503313689|500682785|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|188|Yellow||2013-02-19|2013-02-22|2013-08-29|Volunteer: Time constraint|Volunteer: Time constraint||6.2||4|4|1|1|F|Multi-Race (None of the above)||15||Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||32|28202|Juris Doctorate (JD)|Single|Law: Lawyer|28209|2|5|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|500187654|7|0|2|1|0|2|10|2|-2||4|2|500005291|-2|500000294|-2|0|10|||7496|10|||1|
500791645|502524278|500529175|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|518|Red|2010-2012 OJJDP JJI|2011-04-04|2011-04-28|2012-09-27|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17||4|4|1|1|F|Multi-Race (None of the above)||15||Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||27|28213|Some College|Single|Education|28235|0|6||Relative|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500012459|500187654|7|0|2|31|0|2|10|2|-2||4|3|500005291|-2||-2|0|10|||0|11|||1|500005291
500998933|502274159|500497430|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1113|Red|Amachi|2010-11-18|2010-11-19|2013-12-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||36.6||1|1|1|1|F|Black||15|Yes|Mother|28212|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|Amachi|Match Support|F|White||37|28210|Masters Degree|Single|Medical|28210|1|10|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500015820|500999202|31|0|2|1|0|2|10|2|500003586||4|3|500000294|-2|500000294, 500004640|-2|0|10|||7496|10|||1|500000294
500940594|501174997|500263752|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|267|Red||2008-04-29|2008-05-07|2009-01-29|Child/Family: Time constraints|Child/Family: Time constraints||8.8||1|1|2|2|M|Black||15|No|Mother|28215|One Parent: Female|$25,000 to $29,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||42|28269|Bachelors Degree|Married|Business: Mgt, Admin|28215|10|2|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001267|500940864|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
501716720|501878786|500435676|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2533|Red|Cabarrus County|2010-02-18|2010-03-02|2017-02-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||83.2||1|1|1|1|M|Black||15|No|Mother|28083|One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|Black||52|28075||Married|Medical: Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|501716992|31|0|1|31|0|1|10|2|500016307||4|3|500016374|-2|500016374|-2|6854|8|||7464|9|||1|500016374
503728057|503788318|500763247|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|578|Yellow|Amachi|2014-05-14|2014-05-22|2015-12-21|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||19||1|1|2|2|M|Black||15|Yes|Mother|28227|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||30|28213|Masters Degree|Single|Education|28217|0|7|Recruitment Event|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|503730029|31|0|1|31|0|1|10|2|-2||4|2||-2|500007920, 500011315, 500011316, 500016374|-2|0|10|||7458|9|||1|500000294
502274030|502133187|500477736|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|591|Red||2010-10-07|2010-10-18|2012-05-31|Volunteer: Moved|Volunteer: Moved||19.4||1|1|1|1|F|White||15|No|Mother|28270|One Parent: Female|Unknown||||Yes||Relative|General Community||Enrollment|F|White||38|28205|Bachelors Degree|Married|Tech: Engineer||3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502274462|1|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|3|||7464|9|||1|
503899239|503871007|500770094|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|911|Green||2014-07-21|2014-07-30|2017-01-26|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||29.9||1|1|1|1|M|Black||15|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||38|28269|Some College|Married|Tech: Management|28273|3|1|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503901239|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||17101|1|||1|
503722616|503707316|500759403|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|543|Green||2014-04-11|2014-04-24|2015-10-19|Volunteer: Moved|Volunteer: Moved||17.8||2|2|1|1|F|Multi-race (Black & White)||15|No|Mother|28134|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||55|28217|Some College|Married|Retail: Mgt|28217|14|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503724588|36|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501574833|502189570|500465030|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|381|Green||2010-08-09|2010-08-17|2011-09-02|Volunteer: Time constraint|Volunteer: Time constraint||12.5||2|2|1|1|F|Black||15|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|White||46|28202|Some College|Divorced|Medical: Healthcare Worker|29732|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011184|501575129|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501574833|501452632|500349109|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|498|Green||2009-03-12|2009-03-23|2010-08-03|Volunteer: Time constraint|Volunteer: Time constraint||16.4||2|2|1|1|F|Black||15|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|White||34|28205|Masters Degree|Single|Finance: Accountant|28217|0|3|Recruitment Event|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501575129|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7460|12|||1|
501198008|501043465|500257446|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1165|Green||2008-04-08|2008-04-08|2011-06-17|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38.3||1|1|1|1|F|White||15|No|Mother|28110|One Parent: Female|Unknown||||No||Relative|General Community||Match Support|F|Asian|Indian|33|28105|Bachelors Degree|Single|Business: Clerical||5|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501197566|1|0|2|4|18|2|10|2|-2||4|1||-2||-2|0|3|||46|2|||1|
501247286|501247141|500264655|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|3100|Green||2008-05-05|2008-05-14|2016-11-08|Volunteer: Time constraint|Volunteer: Time constraint||101.8||1|1|1|1|M|White||15|No|Father|28025|One Parent: Male|Unknown||||No||Self|General Community|Cabarrus County|Enrollment|M|White||49|27103|Masters Degree|Single|Education: Teacher|27282|0|0|Other|Service Organization|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500020753|500341682|1|0|1|1|0|1|5|2|-2||4|1|500016374|-2|500016374|-2|0|10|||7452|6|||1|
502328599|502732347|500594124|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|982|Red||2012-01-26|2012-02-22|2014-10-31|Volunteer: Time constraint|Volunteer: Time constraint||32.3||1|1|1|1|M|Black||15|No|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||73|28226|Bachelors Degree|Widowed|Construction||7|0|Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502329034|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|10|||131|1|||1|
501390344|501380163|500342682|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2940|Green|Amachi|2009-02-18|2009-02-26|NaT||||96.6||1|1|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||37|28210|Bachelors Degree|Single|Tech: Computer/Programmer||0|5|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|501390617|31|0|1|1|0|1|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501390345|502966998|500609269|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1773|Green|Amachi|2012-04-11|2012-05-08|NaT||||58.3||2|2|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||35|28206|Bachelors Degree|Single|Business: Sales|28117|4|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|501390617|31|0|1|1|0|1|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501390345|501474303|500342705|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|918|Green|Amachi|2009-02-18|2009-02-26|2011-09-02|Volunteer: Moved|Volunteer: Moved||30.2||2|2|1|1|M|Black||15|Yes|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||29|28206|Some College|Single|Retail: Sales||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011184|501390617|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
503044619|503021454|500624634|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1504|Green||2012-07-18|2012-08-03|2016-09-15|Child/Family: Moved|Child/Family: Moved||49.4||1|1|1|1|M|Black||15|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||29|28202|Bachelors Degree|Single|Finance: Banking|28202|0|7|Self|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500020910|503046265|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
503396873|503381783|500701243|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|175|Green||2013-06-19|2013-08-09|2014-01-31|Child: Lost interest|Child: Lost interest||5.7||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||33|28202|Masters Degree|Single|Arts, Entertainment, Sports||0|0|BBBS National Site|Web Link|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|503398730|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
503043863|502996721|500629081|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|541|Red||2012-08-16|2012-09-04|2014-02-27|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||17.8||1|1|1|1|M|Hispanic||15|No|Mother|28211|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|Asian||32|28204|Bachelors Degree|Single|Medical: Admin|28203|0|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|503045507|3|0|1|4|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501831581|500715453|500387624|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2725|Green|Amachi|2009-09-24|2009-09-29|NaT||||89.5||1|1|2|3|F|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||38|28273||Single|Tech: Engineer||0|8|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501831944|31|0|2|31|0|2|10|2|500003586||2|1|500000294|-2||-2|0|10|||46|2|||1|500000294
502118927|502069043|500455591|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|700|Green||2010-06-04|2010-06-23|2012-05-23|Child/Family: Moved|Child/Family: Moved||23||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||38|28202||Single|Customer Service||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|502099867|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
503071479|503051382|500629193|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1628|Green||2012-08-17|2012-09-30|NaT||||53.5||1|1|1|1|M|Black||15|No|Mother|28216|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||28|28269|Some College|Single|Business: Clerical||0|3|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503069483|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1|
502221871|501239584|500465188|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|128|Yellow||2010-08-10|2010-08-30|2011-01-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.2||2|2|1|1|F|Black||15|No|GrandMother|28216|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||33|28075|Masters Degree|Single|Medical: Healthcare Worker||1|2|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010355|502222302|31|0|2|31|0|2|10|2|-2||4|2|500005291|-2||-2|7016|11|||7496|10|||1|
502221871|501349106|500512728|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|401|Red|2010-2012 OJJDP JJI|2011-01-24|2011-02-24|2012-03-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||13.2||2|2|1|1|F|Black||15|No|GrandMother|28216|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community|2010-2012 OJJDP JJI|Match Support|F|Some Other Race||33|28031|Some College|Single|Tech: Sales, Mktg||1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013709|502222302|31|0|2|41|0|2|10|2|-2||4|3|500005291|-2||-2|7016|11|||7496|10|||1|500005291
501529924|501526581|500338425|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|550|Yellow||2009-02-04|2009-02-06|2010-08-10|Volunteer: Moved|Volunteer: Moved||18.1||2|2|1|1|F|Black||15|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||31|10016|Bachelors Degree|Single|Finance: Banking|28217|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501530213|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501529924|502199360|500465517|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2377|Green||2010-08-12|2010-08-27|2017-02-28|Volunteer: Time constraint|Volunteer: Time constraint||78.1||2|2|1|1|F|Black||15|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||30|28209|Bachelors Degree|Single|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501530213|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
502569117|502538689|500536957|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2116|Green|Amachi, 2010-2012 OJJDP JJI|2011-05-19|2011-05-31|NaT||||69.5||1|1|1|1|F|Black||15|Yes|Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|No||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||40|28269|Masters Degree|Single|Tech: Engineer|77058|6|6|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502569571|31|0|2|31|0|2|10|2|500003586||2|1|500005291|-2||-2|0|10|||17161|11|||1|500000294, 500005291
501261979|500418936|500278634|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2274|Green||2008-07-21|2008-07-22|2014-10-13|Volunteer: Moved|Volunteer: Moved||74.7||1|1|3|3|F|Black||15|No|Mother|28134|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||55|28173||Married|Human Services: Non-Profit|28205|0|0|Coworker|Workplace Partner|Big|General Community|VOL - Maximizing Match Impact|Match Support|1|0|1|0|277|60|598|500000170|500011349|501262256|31|0|2|31|0|2|10|2|-2||4|1||-2|500011314|-2|0|10|||7447|3|||1|
502581001|502650916|500547358|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|917|Red||2011-07-25|2011-07-28|2014-01-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||30.1||1|1|1|1|M|Black||15|No|Mother|28210|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|2010-2012 OJJDP JJI|Match Support|M|Black||37|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28210|0|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500013781|502581504|31|0|1|31|0|1|10|2|-2||4|3|500005291|-2|500000294|-2|34|2|||7496|10|||1|
501536733|501418563|500320917|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2994|Red|Cabarrus County|2008-11-26|2008-11-26|2017-02-06|Child: Severity of challenges|Child: Severity of challenges||98.4||3|3|1|1|F|White||15||Father|28025|One Parent: Male|Unknown||||No||School|General Site|Cabarrus County|Match Support|F|White||44|28037|Bachelors Degree|Married|Business: Sales|28027|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|1|0|0|1|277|60|598|500000170|500022817|501537025|1|0|2|1|0|2|10|2|500016307||4|3|500016374|-1|500016374|-2|0|4|||7464|9|||1|500016374
501220307|501085735|500262676|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1143|Green||2008-04-24|2008-04-30|2011-06-17|Volunteer: Moved|Volunteer: Moved||37.6||1|1|1|1|M|Multi-race (Black & Hispanic)||15|No|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||35|28207|Bachelors Degree|Married|Tech: Engineer||2|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500008062|501220583|38|0|1|1|0|1|10|2|||4|1||-2||-2|0|10|||46|2|||1|
501454635|500188923|500424889|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1350|Red||2010-01-06|2010-01-19|2013-09-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||44.4||1|1|2|2|M|Black||15|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Some Other Race||40|28216|Bachelors Degree|Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|501454920|31|0|1|41|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
501185592|501255830|500270254|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2810|Green||2008-06-06|2008-06-23|2016-03-03|Child: Family structure changed|Child: Family structure changed||92.3|Y|1|1|1|1|M|Multi-race (Black & White)||15|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||45|28211||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501185866|36|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
501771263|501622704|500379993|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2709|Green||2009-08-19|2009-09-29|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||89||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||31|28262|Bachelors Degree|Single|Medical: Admin|28216|0|8|Recruitment Event|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501741899|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7443|2|||1|
503770826|503820142|500761166|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|366|Green||2014-04-25|2014-04-29|2015-04-30|Volunteer: Time constraint|Volunteer: Time constraint||12||1|1|1|1|M|White||15|No|Mother|28211|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||63|28105|Bachelors Degree|Married|Self-Employed, Entrepreneur|28105|7|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503772799|1|0|1|1|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
503328958|503574852|500733114|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1198|Green||2013-11-20|2013-12-04|NaT||||39.4||1|1|1|1|M|Black||15|No|Mother|28213|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||31|28203||Single|Law|28202|3|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|503330792|31|0|1|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
501160611|501508941|500334882|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|189|Green|Amachi|2009-01-22|2009-01-30|2009-08-07|Child/Family: Moved|Child/Family: Moved||6.2||2|2|2|2|M|Black||15|Yes|Mother|28217|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||36|28278|Bachelors Degree|Single|Retail: Sales|30071|5|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|501160885|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501253965|501454688|500327880|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|231|Green|Amachi|2008-12-17|2008-12-18|2009-08-06|Child/Family: Moved|Child/Family: Moved||7.6||3|3|2|2|F|Black||15|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|No||Self|General Community|Amachi|Enrollment|F|White||35|28277|||Education: Teacher|28025|0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001262|503287812|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501253965|502985911|500613577|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1436|Green||2012-05-07|2012-06-11|2016-05-17|Volunteer: Time constraint|Volunteer: Time constraint||47.2||3|3|1|1|F|Black||15|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|No||Self|General Community|Amachi|Enrollment|F|Black||34|28215|Some College|Single|Customer Service||0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503287812|31|0|2|31|0|2|5|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|
502619301|502590110|500552773|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|314|Red|2010-2012 OJJDP JJI|2011-08-31|2011-09-21|2012-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.3||1|1|1|1|F|Hispanic||15|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||RTBM|F|Hispanic||34|28078|Some College|Single|Education: Teacher|28269|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502619917|3|0|2|3|0|2|7|2|500003586||4|3||-2|500004640|-2|0|10|||7462|13|||1|500005291
501526664|501233757|500332719|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1455|Yellow|Amachi|2009-01-14|2009-02-25|2013-02-19|Volunteer: Moved|Volunteer: Moved||47.8||1|1|1|1|F|White||15|Yes|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|F|White||35|28269|Bachelors Degree|Single|Business: Sales|33609|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|501526956|1|0|2|1|0|2|5|2|500003586||4|2|500000294|-2||-2|0|10|||7496|10|||1|500000294
500961274|500403000|500186952|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3489|Green|Amachi|2007-08-02|2007-08-27|NaT||||114.6||1|1|2|2|F|Black||15|Yes|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|Black||51|28216|Bachelors Degree|Divorced|Business: Clerical|28204|20|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|500934638|31|0|2|31|0|2|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
503758675|503792275|500756323|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1085|Green||2014-03-24|2014-03-27|NaT||||35.6||1|1|1|1|M|Black||15|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Black||30|28202|Bachelors Degree|Single|Consultant|28281|2|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503760648|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503704573|503883049|500776636|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|890|Green|PERL 2014-2016|2014-09-18|2014-10-08|NaT||||29.2||1|1|1|1|M|Black||15|No|Mother|28273|One Parent: Female|$20,000 to $24,999||||No||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28277|Bachelors Degree|Single|Business: Marketing|29067|0|3|Man Up Campaign|Media|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|503706538|31|0|1|1|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||17101|1|||1|500014681
502183217|501733851|500462588|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2415|Green|Amachi|2010-07-26|2010-08-05|NaT||||79.3||1|1|2|2|M|Black||15|Yes|Mother|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|Black||50|28078|||Service: Restaurant|28082|0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|502183646|31|0|1|31|0|1|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
503707241|503767700|500759405|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|330|Green||2014-04-11|2014-04-30|2015-03-26|Volunteer: Time constraint|Volunteer: Time constraint||10.8||1|1|1|1|F|Black||15|Yes|Mother|28214|One Parent: Female|$35,000 to $39,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Some Other Race||34|28216|Masters Degree|Living w/ Significant Other|Finance: Banking|28216|0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018850|503709207|31|0|2|41|0|2|5|2|-2||4|1|500000294|-2||-2|34|2|||7464|9|||1|
502896719|502959645|500614239|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1174|Yellow||2012-05-11|2012-06-01|2015-08-19|Volunteer: Moved|Volunteer: Moved||38.6||1|1|1|1|F|Black||15|No|Mother|28269|One Parent: Female|$20,000 to $24,999||||No||Self|General Community||Match Support|F|White||27|28269|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502898127|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
503318449|500716763|500694861|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|280|Green||2013-04-29|2013-05-06|2014-02-10|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||9.2||2|2|2|2|F|Black||15|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||28|28213|Masters Degree|Single|Student: College||0|0||Law Student Association|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503320281|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||0|15|||1|
503318449|503775488|500766059|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|996|Green||2014-06-10|2014-06-24|NaT||||32.7||2|2|1|1|F|Black||15|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||27|28209|Bachelors Degree|Single|Finance|28202|2|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503320281|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501599416|500188567|500357914|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2879|Green||2009-04-17|2009-04-28|NaT||||94.6||1|1|1|1|M|White||14|No|Mother|28262|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||46|28078|Masters Degree|Single|Retail: Mgt|28207|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|501599736|1|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501561529|501333443|500359635|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1206|Green||2009-04-27|2009-05-11|2012-08-29|Volunteer: Moved|Volunteer: Moved||39.6||1|1|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||36|28202|Masters Degree|Single|Business: Sales|28202|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501561821|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502183053|503073638|500621039|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1722|Green||2012-06-22|2012-06-28|NaT||||56.6||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||46|28134|Bachelors Degree|Married|Finance|28105|1|6|Alpha Phi Alpha|Fraternity/Sorority|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|502183482|31|0|1|31|0|1|10|2|-2||2|1||-2|500014681|-2|0|10|||4748|14|633|1|1|
502566369|503065299|500622859|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1703|Green||2012-07-05|2012-07-17|NaT||||56||2|2|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||49|28215|Bachelors Degree|Married|Business: Mgt, Admin|28277|13|0|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502566823|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7439|1|||1|
502566369|502484867|500534744|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|348|Yellow|2010-2012 OJJDP JJI|2011-05-03|2011-05-18|2012-04-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.4||2|2|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||31|28105|Bachelors Degree|Single|Tech: Production Line|28203|3|8|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500011746|502566823|31|0|2|31|0|2|10|2|-2||4|2||-2|500005291|-2|0|10|||7464|9|||1|500005291
503219503|503589945|500746532|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1086|Green||2014-02-03|2014-02-05|2017-01-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.7||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Multi-race (Hispanic & White)||33|28226|Some College|Single|Tech: Management|28277|1|7|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503221284|31|0|1|35|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503816186|501675299|500764043|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|144|Yellow||2014-05-21|2014-05-29|2014-10-20|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||4.7||2|2|1|1|F|Black||14|No|Mother|28206|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||30|28226|Bachelors Degree|Single|Business: Human Resources|28203|0|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|501097065|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502920377|502942994|500620441|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1705|Green||2012-06-19|2012-06-29|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||56||1|1|1|1|F|Black||14|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||31|28211|Bachelors Degree|Single|Real Estate: Realtor|19137|2|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502921794|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501446827|501725833|500368690|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|41|Green||2009-06-12|2009-06-18|2009-07-29|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||1.3||1|1|1|1|M|Black||14|No|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|Black||46|28262|Some College|Divorced|Business|28208|0|8|Local TV|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501447112|31|0|1|31|0|1|5|2|-2||4|1||-2|500000294|-2|0|10|||7438|1|||1|
501215084|501923058|500426321|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|333|Yellow||2010-01-12|2010-01-22|2010-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.9||1|1|1|1|M|Black||14|No|GrandMother|28216|Grandparents|$50,000 to $59,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||33|28078|Bachelors Degree|Divorced|Firefighter||5|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501215360|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|34|2|||7464|9|||1|
503511553|503504991|500702866|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1334|Green||2013-07-08|2013-07-21|NaT||||43.8||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||28|28273|Bachelors Degree||Business|28217|2|0|Elevation Church|Faith Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503513424|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||16414|7|||1|
501553185|501556179|500342698|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1222|Green||2009-02-18|2009-02-23|2012-06-29|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||40.1||1|1|1|1|M|Black||14|No|Mother|28277|One Parent: Female|Unknown||||No|Brochure|Media|General Community||Match Support|M|Black||47|28262|Juris Doctorate (JD)|Married|Law: Lawyer|28262|10|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501553481|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|51|1|||7464|9|||1|
500868942|500947018|500195082|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3465|Green||2007-09-12|2007-09-20|NaT||||113.8|Y|1|1|1|1|M|Black||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999||||No||Self|General Community||Match Support|M|White||54|28207||Married|Business: Sales||0|0|Recruitment Event|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500017732|500869211|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7458|9|||1|
502643010|503262615|500686907|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|488|Yellow||2013-03-08|2013-03-30|2014-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||16||1|1|1|1|M|Black||14|Yes|Mother|28262|One Parent: Female|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Enrollment|M|Black||30|28203|Bachelors Degree|Single|Finance|28255|3|5|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|502643706|31|0|1|31|0|1|5|2|500003586||4|2|500000294|-2|500000294|-2|6854|8|||6247|12|||1|
503110829|503130981|500687926|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1154|Yellow||2013-03-14|2013-03-27|2016-05-24|Volunteer: Moved|Volunteer: Moved||37.9||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|$45,000 to $49,999||||No||Self|General Community||Match Support|M|White||30|28210|Bachelors Degree|Single|Business: Mgt, Admin|28217|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503112489|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502229042|503507627|500704987|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|325|Red||2013-07-26|2013-08-19|2014-07-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.7||3|3|1|1|F|Black||14|No|Mother|28269|Two Parent|Unknown||||Yes||Relative|General Community||Match Support|F|White||54|28210|Some College|Single|Finance: Banking||25|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502172965|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|3|||7464|9|||1|
502229042|502272069|500470500|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|876|Yellow||2010-09-15|2010-09-30|2013-02-22|Volunteer: Time constraint|Volunteer: Time constraint||28.8||3|3|1|1|F|Black||14|No|Mother|28269|Two Parent|Unknown||||Yes||Relative|General Community||Match Support|F|White||35|28211||Single|Business: Sales||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013781|502172965|31|0|2|1|0|2|10|2|-2||4|2||-2|500000294|-2|0|3|||7496|10|||1|
502229042|503849760|500785297|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|243|Red||2014-10-20|2014-10-31|2015-07-01|Volunteer: Moved|Volunteer: Moved||8||3|3|1|1|F|Black||14|No|Mother|28269|Two Parent|Unknown||||Yes||Relative|General Community||Match Support|F|Black||29|28262||Single|Military|28308|5|0|Local TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502172965|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|3|||7438|1|||1|
503634718|503595858|500746721|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1113|Green|Cabarrus County|2014-02-04|2014-02-27|NaT||||36.6||1|1|1|1|F|White||14|No|Father|28081|One Parent: Male|$15,000 to $19,999||||Yes||Self|General Community|Cabarrus County|Match Support|F|White||28|28209|Bachelors Degree|Single|Finance|28217|3|0|Recruitment Event|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500013781|503636659|1|0|2|1|0|2|10|2|-2||2|1|500016374|-2|500016374|-2|0|10|||7458|9|||1|500016374
503961917|504052039|500788399|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|867|Green|PERL 2014-2016, Cabarrus County|2014-10-27|2014-10-31|NaT||||28.5||1|1|1|1|M|White||14|No|Father|28081|One Parent: Male|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|White||28|28277|Bachelors Degree||Finance|28255|0|4|Current/Previous Big|Other Big|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|503636659|1|0|1|1|0|1|10|2|-2||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|5|||17159|12|||1|500014681, 500016374
501160887|501615415|500447312|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1110|Green|Amachi|2010-04-14|2010-04-30|2013-05-14|Volunteer: Time constraint|Volunteer: Time constraint||36.5||2|2|1|1|F|Black||14|Yes|Mother|28208|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Enrollment|F|White||58|28226|||Education: Teacher Asst/Aid|28203|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|501016235|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501160887|501126847|500242032|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|604|Green|Amachi|2008-02-04|2008-02-12|2009-10-08|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||19.8||2|2|1|1|F|Black||14|Yes|Mother|28208|One Parent: Female|Unknown|||Y|No||Self|General Community|Amachi|Enrollment|F|White||31|28227|Bachelors Degree|Single|Medical: Healthcare Worker|28277|0|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501016235|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501938282|502356100|500493871|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2311|Green|Amachi, Cabarrus County|2010-11-11|2010-11-17|NaT||||75.9||1|1|1|1|F|White||14|Yes|Mother|28025|Two Parent|Unknown|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||63|28027|High School Graduate|Married|Self-Employed, Entrepreneur|28027|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|501938680|1|0|2|1|0|2|10|2|500016307||2|1|500000294, 500016374|-2|500016374|-2|0|10|||7464|9|||1|500000294, 500016374
502245129|502670839|500551050|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2033|Green|Amachi|2011-08-22|2011-08-22|NaT||||66.8||1|1|1|1|M|Multi-race (Black & Hispanic)||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||28|28262|High School Graduate|Single|Laborer||0|8|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502245570|38|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1|500000294
500934911|500359073|500221619|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|530|Green|Amachi|2007-11-19|2007-12-06|2009-05-19|Volunteer: Lost contact with child/agency Volunteer: Health|Volunteer: Lost contact with child/agency|Volunteer: Health|17.4||1|1|3|3|M|Black||14|Yes|Mother|28216|One Parent: Female|Less than $10,000|||Y|No||Faith Organization|General Community|Amachi|Enrollment|M|Black||60|28202|Bachelors Degree|Divorced|Tech: Engineer||10|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500935173|31|0|1|31|0|1|5|2|500003586||4|1|500000294|-2|500000294|-2|0|9|||2238|7|||1|500000294
503492214|503551073|500711788|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|49|Red||2013-09-18|2013-10-24|2013-12-12|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||1.6||2|2|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Site|Amachi, mentor2.0, mentor2.0 2016|Match Support|F|White||50|28216|Bachelors Degree|Married|Business: Human Resources|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503494082|31|0|2|1|0|2|10|2|-2||4|3|500000294, 500014505, 500016394|-1||-2|0|10|||7464|9|||1|
503021417|503115600|500631553|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1130|Yellow||2012-08-30|2012-09-11|2015-10-16|Child/Family: Moved|Child/Family: Moved||37.1||1|1|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||32|28204|Bachelors Degree|Single|Business: Marketing|29730|0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|501428579|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502179818|502057930|500460281|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|956|Yellow|Amachi|2010-07-08|2010-07-16|2013-02-26|Volunteer: Moved|Volunteer: Moved||31.4||1|1|1|1|F|Black||14|Yes|GrandMother|28216|Grandparents|Unknown||||Yes|Other|Faith Organization|General Community|Amachi|Enrollment|F|Black||28|28216||Single|Student: College||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|502180247|31|0|2|31|0|2|5|2|500003586||4|2|500000294|-2|500000294|-2|5635|9|||7464|9|||1|500000294
501615769|501567383|500350987|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|124|Green||2009-03-20|2009-04-02|2009-08-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.1||1|1|1|1|F|Black||14|No|Mother|28262|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|F|White||38|28205|Some College||Business: Mgt, Admin|28202|2|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501616089|31|0|2|1|0|2|7|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501662021|502902255|500627357|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|556|Green||2012-08-03|2012-08-14|2014-02-21|Volunteer: Moved|Volunteer: Moved||18.3||2|2|1|1|M|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|Black||50|28269|Some College|Divorced|Retired||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011349|501090456|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501662021|503759352|500757152|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|838|Green||2014-03-27|2014-04-16|2016-08-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||27.5||2|2|1|1|M|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|Black||32|28209|Masters Degree||Finance|28217|0|9|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501090456|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501091420|503668132|500738168|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|265|Green||2013-12-11|2013-12-31|2014-09-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.7||4|4|1|1|M|Black||14||Mother|28206|One Parent: Female|Unknown||||No||School|General Community|PERL 2014-2016|Match Support|M|Black||38|29730|Masters Degree|Married|Human Services: Non-Profit|28212|4|0|TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|501091694|31|0|1|31|0|1|10|2|-2||4|1|500014681|-2||-2|0|4|||130|1|||1|
501091420|503946168|500783556|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|874|Green|PERL 2014-2016|2014-10-14|2014-10-24|NaT||||28.7||4|4|1|1|M|Black||14||Mother|28206|One Parent: Female|Unknown||||No||School|General Community|PERL 2014-2016|Match Support|M|White||29|28205|Bachelors Degree|Single|Finance: Banking|28262|4|0|Man Up Campaign|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|501091694|31|0|1|1|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17100|2|||1|500014681
504081573|503880925|500796131|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|296|Green||2014-11-17|2014-11-25|2015-09-17|Volunteer: Moved|Volunteer: Moved||9.7||2|2|1|1|F|Black||14|No|Mother|28206|One Parent: Female|Unknown|||Y|No||Relative|General Community||Enrollment|F|White||27|28278|Bachelors Degree|Single|Education: Teacher|28056|1|9|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|501091694|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|3|||17159|12|||1|
502000252|502127058|500465318|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2398|Green||2010-08-11|2010-08-22|NaT||||78.8||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||34|28216|Some College||Unemployed||0|0|TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502000651|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||130|1|||1|
502902247|502801082|500619356|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1709|Green||2012-06-14|2012-07-11|NaT||||56.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||30|28203|Bachelors Degree|Single|Business: Marketing|28117|0|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502903657|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502758832|502666962|500586238|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1041|Green||2011-12-12|2011-12-17|2014-10-23|Child: Family structure changed|Child: Family structure changed||34.2||1|1|1|1|F|White||14|No|Mother|28027|One Parent: Female|$50,000 to $59,999||||No||Relative|General Community||Match Support|F|White||33|28027|Masters Degree|Single|Education: Teacher|28027|5|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502759744|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
502569411|502642653|500550403|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|462|Yellow|Amachi, 2010-2012 OJJDP JJI|2011-08-16|2011-09-14|2012-12-19|Child/Family: Time constraints|Child/Family: Time constraints||15.2||1|1|1|1|F|American Indian or Alaska Native||14|Yes|Mother|28213|One Parent: Female|Unknown||||Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|F|White||45|28027|||Medical: Nurse|28144|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502569865|6|0|2|1|0|2|10|2|500003586||4|2|500005291|-2||-2|0|10|||7496|10|||1|500000294, 500005291
502008563|503400112|500730792|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|728|Green||2013-11-13|2013-11-21|2015-11-19|Volunteer: Time constraint|Volunteer: Time constraint||23.9||2|2|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||32|28210|Some College||Business||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|502008962|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
502008563|502053340|500453826|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1153|Green||2010-05-21|2010-06-02|2013-07-29|Volunteer: Moved|Volunteer: Moved||37.9||2|2|1|1|M|Black||14|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||31|28210|Bachelors Degree|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502008962|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501147999|503112265|500665633|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|737|Green||2012-12-03|2013-01-26|2015-02-02|Volunteer: Time constraint|Volunteer: Time constraint||24.2||2|2|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Unknown||||No||School|General Community||Match Support|F|Black||35|28262|Bachelors Degree|Single|Insurance||6|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|501148273|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502700503|502931327|500605634|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1812|Green||2012-03-22|2012-03-30|NaT||||59.5||1|1|1|1|M|Black||14|No|Mother|28217|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||36|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502701348|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503813952|503829786|500763221|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|350|Green||2014-05-13|2014-05-29|2015-05-14|Volunteer: Time constraint|Volunteer: Time constraint||11.5||1|1|1|1|F|Black||14|No|Mother|28262|One Parent: Female|$20,000 to $24,999|||Y|No|BBBS National Site|Web Link|General Community||Enrollment|F|White||28|28202|Masters Degree|Single|Finance: Banking|28205|0|1|Other|Service Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503969639|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|34|2|||7452|6|||1|
501273088|503079327|500659156|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1553|Green||2012-11-13|2012-11-28|2017-02-28|Volunteer: Time constraint|Volunteer: Time constraint||51||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|F|Black||48|28213|Bachelors Degree|Single|Finance: Accountant||8|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501273365|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
501273088|501205202|500277761|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|675|Yellow||2008-07-15|2008-08-23|2010-06-29|Child: Family structure changed|Child: Family structure changed||22.2||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|F|White||38|28210|Masters Degree|Married|Tech: Sales, Mktg|28226|4|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|501273365|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|3|||7464|9|||1|
503952645|503942996|500772607|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|876|Green|PERL 2014-2016, Cabarrus County|2014-08-18|2014-10-22|NaT||||28.8||1|1|1|1|F|White||14|No|Father|28025|One Parent: Male|$40,000 to $44,999|||Y|No|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||31|28025|Bachelors Degree|Married|Business: Mgt, Admin|28027|4|7|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|503954653|1|0|2|31|0|2|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|34|2|||7464|9|||1|500014681, 500016374
502636177|502643313|500551053|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|752|Green||2011-08-22|2011-08-29|2013-09-19|Volunteer: Moved|Volunteer: Moved||24.7||1|1|1|1|F|Black||14|No|GrandMother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|Black||30|28212||Single|Medical||0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502636872|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
501635933|502887536|500601528|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|709|Red||2012-03-01|2012-03-19|2014-02-26|Volunteer: Time constraint|Volunteer: Time constraint||23.3||1|1|1|1|M|Black||14|No|Mother|28202|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||29|28078|Bachelors Degree|Single|Finance|28205|1|0|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501636256|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|10|||7438|1|||1|
501581313|501653852|500360630|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|251|Green||2009-04-30|2009-05-28|2010-02-03|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.2||1|1|1|1|M|Black||14|No|Mother|28211|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||39|28211|||Real Estate: Realtor|28217|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501581615|31|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503838769|503948333|500772925|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|382|Red||2014-08-20|2014-08-30|2015-09-16|Child/Family: Moved|Child/Family: Moved||12.6||1|1|1|1|M|Black||14|No|Mother|28269|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|M|Black||62|28210|Bachelors Degree|Divorced|Business|28202|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503840748|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7671|13|||1|
501069450|500887364|500212043|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3401|Green|Amachi|2007-10-30|2007-11-07|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||111.7||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|M|Black||66|28075||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|501048131|31|0|1|31|0|1|10|2|-2||4|1|500000294|-2||-2|5635|9|||7464|9|||1|500000294
503361148|502459922|500710308|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1269|Green||2013-09-11|2013-09-24|NaT||||41.7||1|1|2|2|M|Multi-race (Black & Hispanic)||14|No|Mother|28273|One Parent: Female|$50,000 to $59,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||59|28226|Bachelors Degree|Married|Business: Sales||0|0|Self|Self|Big|General Community|Project Big|Match Support|0|1|0|1|277|60|598|500000170|500008321|503362993|38|0|1|1|0|1|10|2|-2||2|1||-2|500004640|-2|34|2|||7464|9|||1|
502544579|501718489|500532120|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|735|Yellow|Project Big, 2010-2012 OJJDP JJI|2011-04-20|2011-04-21|2013-04-25|Volunteer: Time constraint|Volunteer: Time constraint||24.1||1|1|1|1|F|Hispanic||14|No|Mother|28213|Two Parent|Unknown||||No||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|Hispanic||35|28078|Bachelors Degree|Married|Human Services: Social Worker|28208|3|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502540313|3|0|2|3|0|2|10|2|500004641||4|2|500004640, 500005291|-2||-2|0|4|||7464|9|||1|500004640, 500005291
502863776|503029273|500622877|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1689|Green||2012-07-05|2012-07-31|NaT||||55.5||1|1|1|1|F|Black||14|No|Mother|28031|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Mgt, Admin|28078|1|11|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502865175|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501014187|501404007|500306699|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3051|Green|Amachi|2008-10-28|2008-11-07|NaT||||100.2||2|2|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|F|White||48|28205|Bachelors Degree|Living w/ Significant Other|Human Services: Non-Profit|28205|3|0|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500013781|500948399|31|0|2|1|0|2|10|2|500003586||2|1|500000294|-2||-2|0|10|||7671|13|||1|500000294
502303088|502445797|500533193|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1890|Green|Project Big|2011-04-25|2011-06-27|2016-08-29|Volunteer: Time constraint|Volunteer: Time constraint||62.1||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community|Project Big|Enrollment|F|Black||33|28215|Bachelors Degree|Single|Human Services: Social Worker|28217|2|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500017777|502303520|31|0|2|31|0|2|5|2|-2||4|1|500004640|-2|500000294, 500004640|-2|6854|8|||7464|9|||1|500004640
502335675|502305990|500495220|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2132|Red|Amachi, Project Big, Project Big AND Amachi|2010-11-16|2010-12-30|2016-10-31|Child: Lost interest|Child: Lost interest||70||1|1|1|1|M|Black||14|Yes|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community|Project Big AND Amachi|Match Support|M|White||27|28262||Single|Self-Employed, Entrepreneur||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500008321|502336110|31|0|1|1|0|1|10|2|500004772||4|3|500004901|-2|500000294, 500004640|-2|0|4|||7496|10|||1|500000294, 500004640, 500004901
503849038|503930671|500778856|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|439|Green||2014-09-29|2014-10-15|2015-12-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.4||1|1|1|1|M|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999||||No||Self|General Community||Match Support|M|Black||32|28202|Bachelors Degree|Single|Consultant|28202|0|9|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503851023|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||17101|1|||1|
502858216|503376842|500687641|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1458|Green||2013-03-13|2013-03-19|NaT||||47.9||1|1|1|1|M|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||32|29708|Bachelors Degree|Married|Finance||0|9|Local TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502859613|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7438|1|||1|
501213488|501225276|500262655|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3223|Green||2008-04-24|2008-05-19|NaT||||105.9||1|1|1|1|F|White||14|No|Father|28207|One Parent: Male|Unknown||||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Finance: Banking|28255|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501213764|1|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
503587461|503541106|500718377|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|595|Green||2013-10-11|2013-10-30|2015-06-17|Child/Family: Time constraints|Child/Family: Time constraints||19.5||1|1|1|1|F|Black||14|Yes|Mother|28262|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||25|28202|Bachelors Degree|Single|Finance|28202|0|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503587387|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502254067|503047588|500677904|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|406|Yellow||2013-01-29|2013-01-31|2014-03-13|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.3||3|3|1|1|F|Black||14|No|Mother|28209|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|Black||39|28213|Bachelors Degree|Married|Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502254499|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502254067|502214352|500466835|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|846|Yellow||2010-08-24|2010-09-10|2013-01-03|Volunteer: Time constraint|Volunteer: Time constraint||27.8||3|3|1|1|F|Black||14|No|Mother|28209|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|Black||37|28210|Bachelors Degree|Single|Insurance||1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502254499|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502254067|503590595|500758482|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1044|Green||2014-04-07|2014-05-07|NaT||||34.3||3|3|1|1|F|Black||14|No|Mother|28209|One Parent: Female|Unknown|||Y|No||Self|General Community||Match Support|F|White||32|28277|Bachelors Degree|Single|Real Estate: Realtor|28202|1|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|502254499|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
502002990|502912865|500599902|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|519|Red||2012-02-23|2012-03-28|2013-08-29|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||17.1||1|1|1|1|M|Black||14||Non-Relative: Other|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes|AARTF|Neighbor/Friend|General Community||Enrollment|M|Asian||32|28204|Bachelors Degree|Single|Finance: Banking||4|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502003389|31|0|1|4|0|1|5|2|500003586||4|3||-2||-2|6855|8|||7496|10|||1|
501537655|501518919|500344393|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|164|Red||2009-02-24|2009-03-13|2009-08-24|Volunteer: Time constraint|Volunteer: Time constraint||5.4||1|1|1|1|M|White||14|No||28027|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||32|28097|Bachelors Degree|Single|Human Services: Non-Profit|28025|0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001262|501537947|1|0|1|1|0|1|7|2|-2||4|3||-2||-2|0|10|||7671|13|||1|
501092822|503854063|500768017|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|968|Green||2014-06-27|2014-07-22|NaT||||31.8||3|4|2|2|F|Black||14|No|Mother|28217|Two Parent|$15,000 to $19,999|||Y|No||School|General Site|mentor2.0, mentor2.0 2016|Match Support|F|White||31|28203|High School Graduate|Single|Business: Sales|28281|3|3|BBBS National Site|Web Link|Big|General Site|mentor2.0, mentor2.0 2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|501093096|31|0|2|1|0|2|10|2|-2||2|1|500014505, 500016394|-1|500014505, 500016394|-1|0|4|||46|2|||1|
503441472|503551607|500738115|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|802|Green||2013-12-11|2014-02-21|2016-05-03|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||26.3||1|1|1|1|F|Black||14|No|Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|No||School|General Community||Match Support|F|Black||28|28216|Masters Degree|Single|Consultant|28205|0|0|Recruitment Event|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500021785|501290021|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||7458|9|||1|
502467122|502658498|500550136|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|39|Green|Amachi|2011-08-15|2011-08-28|2011-10-06|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||1.3||1|1|2|2|M|Black||14|Yes|Mother|28214|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||33|28214|Associate Degree|Single|Law: Security Officer|28208|2|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012319|502467569|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
502034144|502212267|500460434|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1598|Green||2010-07-09|2010-07-20|2014-12-04|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||52.5||1|1|1|1|M|Black||14|No|Mother|28262|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||RTBM|M|Some Other Race||45|28210|Bachelors Degree|Married|Education: Teacher||0|0|CIS/Hidden Valley|Service Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018987|502034543|31|0|1|41|0|1|7|2|||4|1||-2||-2|34|2|||11522|6|||1|
502340295|502881673|500594127|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|22|Green||2012-01-26|2012-02-23|2012-03-16|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||0.7||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Single|Business: Marketing|28036|5|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502340731|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500969483|501344571|500302356|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|269|Green||2008-10-21|2008-11-03|2009-07-30|Volunteer: Time constraint|Volunteer: Time constraint||8.8||2|2|1|1|F|Black||14|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|No||Therapist/Counselor|General Community||Enrollment|F|Black||50|28278|Bachelors Degree|Married|Tech: Engineer|28262|16|0|Volunteer Match|Web Link|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500009007|500969749|31|0|2|31|0|2|5|2|-2||4|1||-2|500000294|-2|0|5|||7444|2|||1|
502545184|501284967|500530934|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|287|Green|2010-2012 OJJDP JJI|2011-04-13|2011-04-15|2012-01-27|Volunteer: Moved|Volunteer: Moved||9.4||1|1|1|1|F|Black||14|No|Mother|28269|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||33|28269|Masters Degree|Single|Business|28269|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502535785|31|0|2|31|0|2|10|2|-2||4|1|500005291|-2||-2|6854|8|||46|2|||1|500005291
502619926|502642260|500548116|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1365|Green|Project Big|2011-07-29|2011-08-09|2015-05-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||44.8||2|2|1|1|F|Black||14|No|GrandMother|28206|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||38|28205|Bachelors Degree|Single|Law: Lawyer|28202|2|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502620542|31|0|2|1|0|2|10|2|500004641||4|1||-2||-2|0|10|||7464|9|||1|500004640
502273093|502252422|500471568|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1642|Green||2010-09-20|2010-10-01|2015-03-31|Child/Family: Moved|Child/Family: Moved||53.9||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||37|28277|PHD|Single|Medical: Healthcare Worker||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|502273525|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|4|||7496|10|||1|
502183420|502264770|500473793|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1570|Yellow|Amachi|2010-09-27|2010-09-28|2015-01-15|Volunteer: Time constraint|Volunteer: Time constraint||51.6||2|2|1|1|M|Multi-race (Black & White)||14|Yes|GrandMother|28215|Grandparents|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|White||58|28226|Masters Degree|Married|Tech: Sales, Mktg|28202|6|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|502183840|36|0|1|1|0|1|10|2|500003586||4|2|500000294|-2||-2|7016|11|||7464|9|||1|500000294
502183420|502202642|500459613|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|11|Green||2010-06-30|2010-07-20|2010-07-31|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||0.4||2|2|1|1|M|Multi-race (Black & White)||14|Yes|GrandMother|28215|Grandparents|Unknown||||Yes|A Child's Place|Service Organization|General Community|Amachi|Match Support|M|Black||54|28212|Some College|Single|Construction||0|0|ACT|Special Event|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|502183840|36|0|1|31|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|7016|11|||7455|8|||1|
503937201|503582646|500772180|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|474|Red||2014-08-13|2014-08-22|2015-12-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||15.6||1|1|1|1|F|Black||14|No|Mother|28031|Two Parent|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|F|White||49|28115|High School Graduate|Single|Customer Service|28115|13|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503939209|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
503913977|503898216|500767515|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|680|Yellow||2014-06-24|2014-06-24|2016-05-04|Child: Family structure changed|Child: Family structure changed||22.3||2|2|2|2|M|White||14|No|GrandMother|28031|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|M|White||61|28202|Masters Degree|Married|Retired||0|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503915984|1|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|4|||17101|1|||1|
501130375|501127478|500245574|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1194|Green|Amachi|2008-02-15|2008-02-15|2011-05-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||39.2||1|1|1|1|M|Black||14|No|Mother|28213|One Parent: Female|Less than $10,000|||Y|Yes||BBBS Board/Staff|General Community|Amachi|Match Support|M|White||33|28202|Masters Degree|Single|Finance: Accountant|28244|0|4|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501130628|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2|500000294|-2|0|13|||2238|7|||1|500000294
502513881|502393006|500615307|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|823|Green||2012-05-17|2012-06-21|2014-09-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27||2|2|3|3|F|Hispanic||14|No|Mother|28262|One Parent: Female|Unknown||||No||School|General Community||Enrollment|F|Black||49|28213|Juris Doctorate (JD)|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502514330|3|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502829894|503443998|500696822|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1385|Yellow||2013-05-14|2013-05-31|NaT||||45.5||2|2|1|1|F|Hispanic||14|No|Mother|28269|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Hispanic||41|28079|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502831178|3|0|2|3|0|2|10|2|-2||2|2||-2||-2|0|4|||7464|9|||1|
502549830|502462453|500538768|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2086|Green|Amachi, Project Big, Project Big AND Amachi|2011-05-26|2011-06-30|NaT||||68.5||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Site|Amachi, Project Big, Project Big AND Amachi|Match Support|M|Black||25|28211||Single|Transport: Driver||0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502550279|31|0|1|31|0|1|10|2|500004772||2|1|500000294, 500004640, 500004901|-1||-2|0|4|||7464|9|||1|500000294, 500004640, 500004901
502560948|502578527|500546411|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|396|Green||2011-07-15|2011-07-31|2012-08-30|Volunteer: Moved|Volunteer: Moved||13||2|2|1|1|F|Black||14|No|Mother|28031|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||39|28078|Masters Degree|Single|Business: Human Resources|28145|5|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|500191427|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502560948|503643705|500742977|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|204|Red||2014-01-15|2014-02-06|2014-08-29|Volunteer: Moved|Volunteer: Moved||6.7||2|2|1|1|F|Black||14|No|Mother|28031|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||25|28031|Some College|Single|Student: College|28031|0|4|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|500191427|31|0|2|31|0|2|5|2|-2||4|3||-2|500000294|-2|0|10|||46|2|||1|
501375862|501832854|500380761|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|30|Green||2009-08-25|2009-08-31|2009-09-30|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||1||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||65|28213|Bachelors Degree|Married|Tech: Engineer|28213|2|9|TV|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500009242|501376141|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||130|1|||1|
502359051|502242295|500483954|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2315|Red|Amachi, Project Big, Project Big AND Amachi|2010-10-21|2010-10-28|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||76.1||1|1|1|1|F|Black||14|Yes|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|Black||35|28213|Masters Degree|Married|Business: Clerical||3|6|Radio|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502359489|31|0|2|31|0|2|10|2|500004772||4|3|500000294, 500004640, 500004901|-2||-2|0|10|||131|1|||1|500000294, 500004640, 500004901
501788776|501698382|500418170|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2607|Green|Amachi|2009-12-03|2010-01-25|NaT||||85.7||1|1|1|1|M|Black||14|Yes|Mother|28214|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||64|28117||Married|Business: Sales|28031|0|0|Alpha Kappa Alpha|Fraternity/Sorority|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501789128|31|0|1|1|0|1|10|2|500003586||2|1|500000294|-2||-2|0|10|||8697|14|||1|500000294
502825916|502367677|500589764|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1879|Yellow|Amachi|2012-01-04|2012-01-23|NaT||||61.7||1|1|2|2|F|Black||14|Yes|Mother|28273|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||36|28208|Some College|Single|Education: Teacher|28226|1|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500008321|502827199|31|0|2|31|0|2|10|2|-2||2|2|500000294|-2|500000294, 500004640|-2|0|10|||7464|9|||1|500000294
502753873|503146044|500691867|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1424|Green||2013-04-08|2013-04-22|NaT||||46.8||2|2|1|1|F|Hispanic||14|No|Mother|28262|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||43|28216|Masters Degree|Single|Finance: Accountant|28685|1|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502751081|3|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
502753873|502896683|500596765|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|359|Yellow||2012-02-07|2012-02-29|2013-02-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.8||2|2|1|1|F|Hispanic||14|No|Mother|28262|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||27|28269|Bachelors Degree|Single|Finance|28227|0|5|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502751081|3|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
502186245|502268901|500470155|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|316|Yellow||2010-09-13|2010-09-15|2011-07-28|Volunteer: Time constraint|Volunteer: Time constraint||10.4||3|3|1|1|F|Black||14|No|Mother|28216|Two Parent|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||37|28211||Single|Business: Mgt, Admin||10|2|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501610196|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502186245|502605983|500548277|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|735|Green|Project Big|2011-08-01|2011-08-18|2013-08-22|Volunteer: Moved|Volunteer: Moved||24.1||3|3|1|1|F|Black||14|No|Mother|28216|Two Parent|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|White||33|28203||Single|Business|28211|3|6|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500004169|501610196|31|0|2|1|0|2|10|2|500004641||4|1||-2|500000294, 500004640|-2|0|10|||7464|9|||1|500004640
503016111|503135600|500636811|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1607|Red||2012-09-19|2012-09-30|2017-02-23|Volunteer: Time constraint|Volunteer: Time constraint||52.8||1|1|1|1|M|Black||14|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|Black||32|28216|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|503013381|31|0|1|31|0|1|10|2|500003586||4|3|500000294|-2|500000294|-2|0|10|||7496|10|||1|
502436198|502446619|500520591|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|594|Green||2011-02-28|2011-03-17|2012-10-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.5||2|2|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||51|28205|Masters Degree|Married|Education: Teacher|28212|14|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502436641|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
502436198|503255826|500701262|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1358|Green||2013-06-19|2013-06-27|NaT||||44.6||2|2|1|1|F|Black||14|No|Mother|28212|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||31|28209|Masters Degree|Single|Medical|28207|0|5|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502436641|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1|
502567552|502208867|500538510|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|420|Red|Amachi, Project Big, Project Big AND Amachi|2011-05-25|2011-06-07|2012-07-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||13.8||1|1|2|2|F|Hispanic||14|Yes|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||25|28262||Single|Student: College||0|0|Self|Self|Big|General Community|Project Big AND Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011746|502568002|3|0|2|31|0|2|10|2|500004772||4|3|500004640, 500004901|-2|500004901|-2|0|4|||7464|9|||1|500000294, 500004640, 500004901
502404516|502624164|500548056|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|666|Red||2011-07-29|2011-08-23|2013-06-19|Volunteer: Moved|Volunteer: Moved||21.9||1|1|1|1|M|White||14|No|Mother|28273|One Parent: Female|Unknown||||No|Yahoo!|Web Link|General Community||Enrollment|M|White||49|19711|Bachelors Degree|Living w/ Significant Other|Business: Marketing|28278|15|2|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500004169|502404954|1|0|1|1|0|1|5|2|-2||4|3||-2|500004640|-2|30|2|||7464|9|||1|
503643026|503377601|500761779|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|535|Red||2014-04-30|2014-05-09|2015-10-26|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17.6||3|3|2|2|F|Black||14|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||30|28213|Some College|Single|Medical|28209|1|4|Self|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500020990|503644986|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503643026|503603792|500731516|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|107|Yellow||2013-11-15|2013-11-26|2014-03-13|Volunteer: Time constraint|Volunteer: Time constraint||3.5||3|3|1|1|F|Black||14|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Business: Human Resources||1|3|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|503644986|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7671|13|||1|
501143676|503315012|500683363|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|866|Red||2013-02-21|2013-02-28|2015-07-14|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||28.5||1|1|1|1|M|Black||14|No|Mother|28213|One Parent: Female|$10,000 to $14,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||50|28269|Associate Degree|Married|Self-Employed, Entrepreneur||12|0|Newspaper|Media|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|501143950|31|0|1|31|0|1|10|2|-2||4|3||-2|500000294|-2|34|2|||129|1|||1|
503803127|503866013|500766041|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|993|Green||2014-06-10|2014-06-27|NaT||||32.6||1|1|1|1|M|Black||14|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Match Support|M|Black||42|28270|Bachelors Degree|Married|Unknown||0|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503798593|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|4|||17101|1|||1|
502261654|502264865|500470591|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|388|Green||2010-09-15|2010-09-20|2011-10-13|Volunteer: Time constraint|Volunteer: Time constraint||12.7|Y|1|1|1|1|M|Black||14|No|Mother|28209|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||37|28211|Bachelors Degree|Married|Business: Mgt, Admin|28210|7|0|Big Champions|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011639|502262086|31|0|1|1|0|2|5|2|-2||4|1||-2||-2|6854|8|||7461|12|||1|
501295653|501374940|500331192|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|970|Green||2009-01-08|2009-01-15|2011-09-12|Volunteer: Time constraint|Volunteer: Time constraint||31.9||1|1|1|1|M|White||14|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|White||43|28025|Some College|Divorced|Business: Mgt, Admin|28107|3|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501295931|1|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
503524258|500497043|500713184|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|848|Green||2013-09-25|2013-09-30|2016-01-26|Volunteer: Moved|Volunteer: Moved||27.9||1|1|3|3|F|Black||14|No|Mother|28217|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|Black||34|28273|Bachelors Degree|Single|Retail: Mgt|28217|5|6|AA Task Force|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503526133|31|0|2|31|0|2|5|2|-2||4|1|500000294|-2||-2|34|2|||6247|12|||1|
503544893|503844843|500777054|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|375|Yellow||2014-09-19|2014-09-26|2015-10-06|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.3||1|1|2|2|F|Black||14|No|Mother|28227|One Parent: Female|$20,000 to $24,999|Yes: Active|No|Y|Yes||Self|General Community||Match Support|F|Black||46|28216|Bachelors Degree|Single|Business: Marketing|28036|0|3|Self|Self|Big|General Community|VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500012459|503546768|31|0|2|31|0|2|10|2|-2||4|2||-2|500007920, 500011312, 500011315, 500011316|-2|0|10|||7464|9|||1|
502255156|502946412|500608992|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1787|Green|Amachi|2012-04-10|2012-04-24|NaT||||58.7||2|2|1|1|F|Black||14|Yes|Relative: Other|28227|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|White||35|28277|Masters Degree|Single|Education: Admin||8|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502255582|31|0|2|1|0|2|10|2|500003586||2|1|500000294|-2||-2|0|5|||7462|13|||1|500000294
502255156|502165697|500512286|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|330|Green|Amachi|2011-01-20|2011-02-14|2012-01-10|Volunteer: Moved|Volunteer: Moved||10.8||2|2|1|1|F|Black||14|Yes|Relative: Other|28227|One Parent: Female|Unknown||||Yes||Therapist/Counselor|General Community|Amachi|Match Support|F|Black||34|28227|Some College|Single|Medical: Healthcare Worker||0|7|AA Task Force|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502255582|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|5|||6247|12|||1|500000294
502529397|500188946|500548763|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2044|Green|Project Big|2011-08-04|2011-08-11|NaT||||67.2||1|1|2|2|M|Black||14|No|Mother|28216|One Parent: Female|$30,000 to $34,999||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||48|28216|Bachelors Degree|Married|Finance: Banking|28255|8|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502529850|31|0|1|31|0|1|10|2|500004641||2|1||-2||-2|6854|8|||7464|9|||1|500004640
503479095|503915425|500768983|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|621|Green||2014-07-09|2014-07-17|2016-03-29|Volunteer: Moved|Volunteer: Moved||20.4||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Enrollment|M|White||28|28270|Bachelors Degree|Married|Real Estate: Realtor|28203|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503480961|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501863951|501601161|500421259|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1988|Red||2009-12-14|2009-12-18|2015-05-29|Child: Lost interest|Child: Lost interest||65.3||1|1|2|2|F|Black||14|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Black||37|28078|Bachelors Degree|Single|Business: Human Resources|28226|0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501864324|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503021552|502951522|500618601|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1220|Yellow||2012-06-08|2012-06-19|2015-10-22|Volunteer: Moved|Volunteer: Moved||40.1||1|1|1|1|F|Black||14|No|Mother|28270|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Multi-Race (None of the above)||28|28215|Some College|Single|Insurance||0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503023091|31|0|2|7|0|2|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503497835|503507978|500710423|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1274|Green||2013-09-11|2013-09-19|NaT||||41.9||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|Black||26|28209|Bachelors Degree|Single|Retail: Sales|28210|0|10|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503499703|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503470435|503597172|500757513|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|91|Green||2014-03-31|2014-03-31|2014-06-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3||1|1|1|1|M|White||14|No|Mother|28214|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||40|28205|Bachelors Degree|Separated|Construction|28205|4|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017732|503472301|1|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
503429736|503850437|500760086|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1052|Green||2014-04-17|2014-04-29|NaT||||34.6||1|1|1|1|M|Black||14|No|Mother|28216|One Parent: Female|$60,000 to $74,999|Yes: Active|Yes||No|AARTF|Neighbor/Friend|General Community||Match Support|M|White||27|28217|Masters Degree|Single|Finance|28202|0|7|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503431601|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|6855|8|||17159|12|||1|
501345383|501083988|500325591|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|154|Green|Amachi|2008-12-11|2008-12-18|2009-05-21|Vol: Other Reason Child/Family: Feels incompatible with volunteer|Vol: Other Reason|Child/Family: Feels incompatible with volunteer|5.1||2|2|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||41|28278|Associate Degree|Single|Human Services: Social Worker|28211|1|4|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|501345662|31|0|2|1|0|2|10|2|500003586||4|1|500000294|-2||-2|34|2|||7464|9|||1|500000294
501345383|501484003|500392320|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1141|Yellow|Amachi|2009-10-07|2009-10-28|2012-12-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||37.5||2|2|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|White||31|28273|Bachelors Degree|Single|Service: Restaurant|28269|0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|501345662|31|0|2|1|0|2|10|2|500003586||4|2|500000294|-2||-2|34|2|||7462|13|||1|500000294
502943644|503899413|500771637|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|431|Red||2014-08-07|2014-08-25|2015-10-30|Volunteer: Time constraint|Volunteer: Time constraint||14.2||2|2|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|Black||23|28213||Single|Arts, Entertainment, Sports||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502945070|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503166335|503335465|500683005|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|554|Red||2013-02-20|2013-03-19|2014-09-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.2||2|2|1|1|F|White||14|No|Mother|28031|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|F|White||34|28031|Bachelors Degree|Single|Business: Marketing|28031|6|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503168022|1|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503166335|503729353|500796127|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|410|Yellow||2014-11-17|2014-11-24|2016-01-08|Child: Lost interest|Child: Lost interest||13.5||2|2|1|1|F|White||14|No|Mother|28031|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|F|White||31|28036|Associate Degree|Single|Medical|28202|6|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503168022|1|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502672482|502621665|500566301|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|681|Red|Project Big|2011-10-17|2011-10-18|2013-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||22.4||1|1|1|1|M|Hispanic||14|No|Mother|28208|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Project Big|Match Support|M|White||27|28209|Bachelors Degree|Single|Tech: Support, Writing|29707|0|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502673310|3|0|1|1|0|1|10|2|500004641||4|3|500004640|-2||-2|0|10|||7464|9|||1|500004640
502635070|502823119|500581061|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|239|Green|Amachi|2011-11-22|2012-01-05|2012-08-31|Volunteer: Time constraint|Volunteer: Time constraint||7.9||1|1|1|1|M|Multi-race (Black & Hispanic)||14|Yes|Mother|28269|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community|Amachi|RTBM|M|White||31|28202|Masters Degree|Single|Finance: Auditor|28202|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502635764|38|0|1|1|0|1|7|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
502875279|502864263|500600651|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1003|Red||2012-02-27|2012-03-19|2014-12-17|Volunteer: Time constraint|Volunteer: Time constraint||33||2|2|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||32|28210|Bachelors Degree|Single|Business: Sales||2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502876679|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502934735|502992001|500660486|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|211|Yellow||2012-11-15|2012-11-19|2013-06-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.9||1|1|1|1|F|Black||14|No|Mother|28269|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|F|White||51|28031|Some College|Married|Finance: Banking||7|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502936158|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503017622|503095382|500631726|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1639|Green||2012-08-31|2012-09-19|NaT||||53.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|$30,000 to $34,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|F|White||33|28207|Bachelors Degree|Married|Business||0|7|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503019155|31|0|2|1|0|2|10|2|-2||3|1||-2||-2|34|2|||7464|9|||1|
501704517|501775116|500375074|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|329|Red||2009-07-22|2009-07-29|2010-06-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.8||1|1|1|1|M|Black||14|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|Black||47|28215||Single|Unknown||0|0|Other|BBBS Board/Staff|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500008629|501704855|31|0|1|31|0|1|5|2|-2||4|3||-2|500000294|-2|0|10|||7671|13|||1|
502945480|502919780|500603409|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1813|Green||2012-03-12|2012-03-29|NaT||||59.6||1|1|1|1|F|Black||14|No|Mother|28215|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||54|28262|Bachelors Degree|Single|Business: Mgt, Admin||0|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502946906|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501142903|501236825|500268808|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3206|Green|Amachi|2008-05-28|2008-06-05|NaT||||105.3||1|1|1|1|M|Black||14|Yes|GrandMother|28208|One Parent: Female|Less than $10,000||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Match Support|M|White||53|28204|Juris Doctorate (JD)|Married|Law: Lawyer|28244|16|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|501143177|31|0|1|1|0|1|10|2|500003586||2|1|500000294|-2|500000294|-2|7294|13|||2238|7|||1|500000294
501721579|501687513|500375006|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2520|Red|Amachi|2009-07-22|2009-07-24|2016-06-17|Volunteer: Moved|Volunteer: Moved||82.8||2|2|1|1|F|Multi-Race (None of the above)||14|No|Mother|28211|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||50|28227|Some College|Single|Human Services: Social Worker||2|5|St. Paul Baptist|Faith Organization|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|501721919|7|0|2|31|0|2|10|2|500003586||4|3|500000294|-2|500000294|-2|5635|9|||9609|7|||1|500000294
501721579|501351593|500357749|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|91|Green|Amachi|2009-04-16|2009-04-21|2009-07-21|Volunteer: Time constraint|Volunteer: Time constraint||3||2|2|1|1|F|Multi-Race (None of the above)||14|No|Mother|28211|One Parent: Female|Unknown||||No|Other|Faith Organization|General Community|Amachi|Match Support|F|Black||37|28216|Bachelors Degree|Single|Medical: Admin|28203|10|0|Recruitment Event|Workplace Partner|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500003657|501721919|7|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|5635|9|||7446|3|||1|500000294
502902269|501631588|500677452|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|391|Yellow||2013-01-26|2013-01-26|2014-02-21|Child: Lost interest|Child: Lost interest||12.8||1|1|3|3|M|Black||14|No|Mother|28215|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Enrollment|M|Black||31|28203|Juris Doctorate (JD)||Law: Lawyer|28203|1|0|Self|Self|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500011349|502903679|31|0|1|31|0|1|5|2|-2||4|2||-2|500015184|-1|0|10|||7464|9|||1|
503381531|500540549|500762593|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1015|Green||2014-05-08|2014-06-05|NaT||||33.3||1|1|2|2|M|Black||14|No|Mother|28206|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||66|28269||Married|Retired||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503383388|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503070961|503034904|500628328|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|764|Red|Amachi|2012-08-13|2012-08-21|2014-09-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||25.1||1|1|1|1|F|Black||14|Yes|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community|Amachi|Match Support|F|White||29|28209|||Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503072625|31|0|2|1|0|2|10|2|-2||4|3|500000294|-2||-2|0|4|||7464|9|||1|500000294
501397326|501371039|500336441|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|150|Green|Amachi|2009-01-28|2009-02-20|2009-07-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||4.9||1|1|1|1|M|Black||14|Yes|Mother|28025|One Parent: Female|Unknown|||Y|Yes|Other|Faith Organization|General Community|Amachi|Enrollment|M|Black||56|28075||Married|Unknown||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500001262|501397607|31|0|1|31|0|1|5|2|500003586||4|1|500000294|-2|500000294|-2|5635|9|||7453|7|||1|500000294
502264663|502080569|500503506|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|229|Green||2010-12-08|2010-12-30|2011-08-16|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||7.5||2|2|2|2|F|Multi-race (Black & White)||14|No|Mother|28206|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community||Match Support|F|White||33|28078|High School Graduate|Single|Self-Employed, Entrepreneur|28269|0|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|502265095|36|0|2|1|0|2|10|2|-2||4|1||-2||-2|5635|9|||7464|9|||1|
502264663|502590405|500562787|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|369|Green||2011-10-07|2012-01-06|2013-01-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.1||2|2|1|1|F|Multi-race (Black & White)||14|No|Mother|28206|One Parent: Female|Unknown||||Yes|Other|Faith Organization|General Community||Match Support|F|White||32|28205|Bachelors Degree|Single|Human Services: Youth Worker|28203|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502265095|36|0|2|1|0|2|10|2|-2||4|1||-2||-2|5635|9|||7496|10|||1|
502570185|502191626|500542078|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1050|Yellow|Amachi, Project Big, Project Big AND Amachi, 2010-2012 OJJDP JJI|2011-06-20|2011-06-30|2014-05-15|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.5||1|1|1|1|F|Black||14|No|Mother|28206|Other/Unknown|Unknown||||Yes||Relative|General Community|2010-2012 OJJDP JJI, Project Big|Enrollment|F|Black||58|28226|Masters Degree|Single|Tech: Management|28078|0|2|BBBS National Site|Web Link|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500017777|502570639|31|0|2|31|0|2|5|2|500004641||4|2|500004640, 500005291|-2|500004640|-2|0|3|459|3|46|2|||1|500000294, 500004640, 500004901, 500005291
501721762|502884274|500612996|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|113|Green||2012-05-02|2012-05-15|2012-09-05|Volunteer: Moved|Volunteer: Moved||3.7||3|3|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||41|28278|Masters Degree|Living w/ Significant Other|Tech: Computer/Programmer|30005|5|0|BBBS National Site|Web Link|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|501722098|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501721762|503471102|500700196|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1359|Green||2013-06-11|2013-06-26|NaT||||44.6||3|3|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||39|28211||Single|Retail: Sales||0|11|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501722098|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501721762|501278761|500368878|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|932|Green||2009-06-15|2009-06-22|2012-01-10|Volunteer: Time constraint|Volunteer: Time constraint||30.6||3|3|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||36|28213|Some College|Married|Customer Service|28262|1|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008629|501722098|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
501721761|501951880|500432328|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|350|Red||2010-02-04|2010-02-24|2011-02-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||11.5||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||31|28213|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501722098|31|0|1|1|0|1|7|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501721761|503023854|500618753|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1127|Yellow||2012-06-11|2012-06-25|2015-07-27|Volunteer: Time constraint|Volunteer: Time constraint||37||2|2|1|1|M|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||31|28210|Bachelors Degree|Single|Retail: Sales||1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|501722098|31|0|1|1|0|1|7|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502236953|502232559|500464143|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1627|Red||2010-08-04|2010-08-17|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||53.5||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||50|28212|Some College|Married|Law: Police Officer||2|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|502237384|31|0|1|31|0|1|10|2|-2||4|3||-2|500000294|-2|0|10|||7464|9|||1|
502495686|502755977|500581022|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|175|Yellow||2011-11-22|2011-12-16|2012-06-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||5.7||1|1|1|1|M|Hispanic||14|No|Mother|28212|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|M|Hispanic||28|28212||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502496135|3|0|1|3|0|1|10|2|-2||4|2||-2||-2|0|4|||7464|9|||1|
502308197|502325667|500493122|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1984|Green||2010-11-10|2010-12-03|2016-05-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||65.2||1|1|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|F|White||35|28210|Bachelors Degree|Living w/ Significant Other|Business: Sales|18034|2|7|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big AND Amachi|Match Support|0|1|0|1|277|60|598|500000170|500021785|502308629|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294, 500004901|-2|0|10|||7496|10|||1|
502506397|503039829|500619509|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1585|Yellow||2012-06-15|2012-06-30|2016-11-01|Child: Severity of challenges|Child: Severity of challenges||52.1||1|1|1|1|F|White||14|No|Mother|28210|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||33|28277|Bachelors Degree|Single|Consultant|28202|1|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502506846|1|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502794252|503351102|500696692|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|455|Red||2013-05-13|2013-05-31|2014-08-29|Volunteer: Time constraint|Volunteer: Time constraint||14.9||2|2|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|White||30|28202|Bachelors Degree|Single|Business|28203|1|6|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|502129968|31|0|2|1|0|2|5|2|-2||4|3||-2|500000294|-2|0|10|||7464|9|||1|
502794252|502725901|500584551|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|333|Green||2011-12-06|2011-12-16|2012-11-13|Volunteer: Time constraint|Volunteer: Time constraint||10.9||2|2|1|1|F|Black||14|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|Black||28|28212|Some College|Single|Customer Service||0|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502129968|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
502507408|502673562|500559678|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1775|Yellow|2010-2012 OJJDP JJI|2011-09-29|2011-10-13|2016-08-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||58.3||1|1|1|1|M|Black||14|No|Mother|28226|One Parent: Female|Less than $10,000||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||71|28277|Bachelors Degree|Married|Retired||0|0||Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502507857|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|34|2|||0|11|||1|500005291
503170936|503258884|500674088|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|8|Green||2013-01-10|2013-01-23|2013-01-31|Child: Severity of challenges|Child: Severity of challenges||0.3||1|1|2|2|M|White||14|No|Mother|28277|Grandparents|Less than $10,000||||Yes||Therapist/Counselor|General Community||Match Support|M|Asian|Indian|27|28277|Bachelors Degree|Single|Business|28277|0|2||Relative|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500004169|503172623|1|0|1|4|18|1|10|2|-2||4|1||-2||-2|0|5|||0|11|||1|
501615994|500757448|500370013|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|413|Green|Amachi|2009-06-18|2009-06-22|2010-08-09|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.6|Y|1|1|2|2|M|Black||14|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|RTBM|F|Black||59|28216||Married|Business: Human Resources||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500003657|501616314|31|0|1|31|0|2|7|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501295538|501207855|500265791|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1001|Green||2008-05-13|2008-05-13|2011-02-08|Volunteer: Time constraint|Volunteer: Time constraint||32.9||2|2|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|Black||33|28217|Bachelors Degree|Single|Business: Clerical||0|7|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500740560|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
501295538|502897530|500603727|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1812|Green||2012-03-13|2012-03-30|NaT||||59.5||2|2|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||31|28078|Bachelors Degree||Medical||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|500740560|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503756716|503596238|500754325|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|654|Green||2014-03-12|2014-03-31|2016-01-14|Child: Lost interest|Child: Lost interest||21.5||1|1|1|1|F|Black||14|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||29|28270||Single|Unemployed||0|0|Self|Self|Big|General Community|Amachi|Enrollment|0|1|0|1|277|60|598|500000170|500020990|503758688|31|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
503061519|503115965|500646319|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|651|Green||2012-10-16|2012-10-31|2014-08-13|Child/Family: Moved|Child/Family: Moved||21.4||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||27|28031|Bachelors Degree|Married|Business: Mgt, Admin|28205|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|503063175|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|34|2|||7496|10|||1|
501209738|501608996|500380528|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|412|Green|Amachi|2009-08-24|2009-09-09|2010-10-26|Volunteer: Moved|Volunteer: Moved||13.5||2|2|1|1|F|Black||14|Yes|Mother|28206|One Parent: Female|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Enrollment|F|White||33|28211|||Consultant|28202|0|0|Self|Self|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500003657|501210012|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|7294|13|||7464|9|||1|500000294
501209738|502351250|500502375|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|699|Yellow|Amachi|2010-12-06|2011-01-24|2012-12-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||23||2|2|1|1|F|Black||14|Yes|Mother|28206|One Parent: Female|Unknown||||Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Enrollment|F|White||29|28211|Some College|Single|Student: College||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|501210012|31|0|2|1|0|2|5|2|-2||4|2|500000294|-2|500000294|-2|7294|13|||7464|9|||1|500000294
502225378|502245842|500509780|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2241|Green||2011-01-07|2011-01-26|NaT||||73.6||1|1|1|1|M|White||14|No|Mother|28277|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||67|28277|Bachelors Degree|Divorced|Tech: Sales, Mktg||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|502225809|1|0|1|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
503452963|503489818|500705904|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|517|Red||2013-08-06|2013-08-22|2015-01-21|Volunteer: Time constraint|Volunteer: Time constraint||17||1|1|1|1|M|Black||14|No|Mother|28211|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|Black||41|28216|Bachelors Degree|Single|Customer Service|28262|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503430105|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
503717073|503853194|500762798|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|882|Green||2014-05-09|2014-05-16|2016-10-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||29||1|1|1|2|M|Black||14|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|Black||54|28277|Bachelors Degree|Single|Consultant|28202|7|6|Man Up Campaign|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Pending Match|0|1|0|1|277|60|598|500000170|500020910|503719040|31|0|1|31|0|1|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|4|||17101|1|||1|
502336272|503743688|500752685|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1093|Green||2014-03-04|2014-03-19|NaT||||35.9||2|2|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||35|27713|Associate Degree|Single|Business|28216|0|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502336707|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|6854|8|||7464|9|||1|
502336272|502363052|500502396|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1049|Yellow||2010-12-06|2011-01-07|2013-11-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||34.5||2|2|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||31|28208|Bachelors Degree|Single|Business: Sales||0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502336707|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1|
501222138|500189173|500447311|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1833|Yellow|Amachi|2010-04-14|2010-04-30|2015-05-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||60.2||2|2|2|3|F|Black||14|Yes|GrandMother|28227|Grandparents|Unknown||||No||Self|General Community|Amachi|Enrollment|F|Black||53|28269|Some College|Married|Business: Sales|28227|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500012459|501222414|31|0|2|31|0|2|5|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
501222138|501238738|500268752|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|389|Green|Amachi|2008-05-28|2008-05-30|2009-06-23|Volunteer: Moved|Volunteer: Moved||12.8||2|2|1|1|F|Black||14|Yes|GrandMother|28227|Grandparents|Unknown||||No||Self|General Community|Amachi|Enrollment|F|White||36|28277|Bachelors Degree|Single|Unknown||5|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|501222414|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||2238|7|||1|500000294
503972507|500189600|500780309|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|868|Green||2014-10-03|2014-10-13|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||28.5||1|1|2|2|F|Black||14|Yes|Mother|28278|One Parent: Female|$50,000 to $59,999|||Y|No||Self|General Community||Match Support|M|Black||46|28214|Bachelors Degree|Single|Finance: Economist|28217|14|0|Brochure|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503974518|31|0|2|31|0|1|10|2|500003586||4|1||-2||-2|0|10|||127|1|||1|
502222545|502196116|500462566|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|2366|Green||2010-07-26|2010-08-03|2017-01-24|Volunteer: Time constraint|Volunteer: Time constraint||77.7||1|1|1|1|F|Black||14|No|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|F|White||37|28208|Masters Degree|Single|Education: Teacher||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|502222979|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502255210|502255794|500470233|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2362|Green||2010-09-14|2010-09-27|NaT||||77.6||1|1|1|1|M|Black||14|No|Mother|28214|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||29|28210|Bachelors Degree|Married|Business: Mgt, Admin|97224|6|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020752|500910307|31|0|1|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7496|10|||1|
501955315|501972860|500427129|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|150|Red||2010-01-15|2010-01-29|2010-06-28|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||4.9||1|1|1|1|M|Black||14|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|Black||61|28212|||Retired||0|0|Local TV|Media|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010765|501955713|31|0|1|31|0|1|7|2|-2||4|3||-2|500000294|-2|0|10|||7438|1|||1|
501254255|501356688|500282157|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3080|Green||2008-08-15|2008-09-23|2017-02-28|Volunteer: Moved|Volunteer: Moved||101.2||1|1|1|1|F|Black||14|No|Mother|28230|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||34|28205|Masters Degree|Single|Finance: Banking|28217|0|4|Yahoo!|Web Link|Big|General Community|Amachi|Match Support|1|0|0|1|277|60|598|500000170|500013781|501254531|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||32|2|||1|
502568949|502626358|500547244|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|245|Green|Amachi|2011-07-22|2011-07-29|2012-03-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||8||1|1|1|1|M|Black||14|Yes|Mother|28208|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community|Amachi|Match Support|M|White||30|28202|Masters Degree|Single|Finance|28202|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502569403|31|0|1|1|0|1|10|2|500003586||4|1|500000294|-2||-2|0|10|||7496|10|||1|500000294
502866443|502920462|500613414|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|831|Red||2012-05-04|2012-06-14|2014-09-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27.3||1|1|1|1|F|Black||14|No|Mother|28262|One Parent: Female|$30,000 to $34,999|||Y|No||Self|General Community||Match Support|F|Black||38|28212|Some College|Single|Business: Mgt, Admin|28270|7|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502867844|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502197486|502870668|500597982|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1849|Green||2012-02-13|2012-02-22|NaT||||60.7||1|1|1|1|M|Black||14|No|Mother|28212|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||30|28209|Bachelors Degree|Single|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502197915|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|
503953654|503976139|500775808|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|888|Green|PERL 2014-2016|2014-09-15|2014-10-10|NaT||||29.2||1|1|1|1|M|Black||14|Yes|Mother|28208|One Parent: Female|Less than $10,000|||Y|No||Therapist/Counselor|General Community|Amachi, PERL 2014-2016|Match Support|M|White||28|28209|Bachelors Degree|Single|Tech: Engineer||0|5|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020752|503955662|31|0|1|1|0|1|10|2|-2||2|1|500000294, 500014681|-2|500014681|-2|0|5|||46|2|||1|500014681
502255223|501823103|500463922|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2409|Green||2010-08-03|2010-08-11|NaT||||79.1||1|1|1|1|F|Hispanic||14|No|Mother|28212|One Parent: Female|Unknown|||Y|No|Spanish Radio|Media|General Community||Match Support|F|White||33|28209||Single|Education: Teacher||0|0||High School Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502255655|3|0|2|1|0|2|10|2|-2||2|1||-2||-2|7068|1|||0|4|||1|
502583662|503943422|500783380|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|211|Yellow||2014-10-14|2014-10-28|2015-05-27|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||6.9||3|3|1|1|F|Black||14|No|GrandMother|28215|Grandparents|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|F|Black||50|28215|Associate Degree|Married|Medical: Nurse||2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502584168|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|4|||7464|9|||1|
502583662|503515217|500706497|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|293|Red||2013-08-12|2013-08-30|2014-06-19|Volunteer: Time constraint|Volunteer: Time constraint||9.6||3|3|1|1|F|Black||14|No|GrandMother|28215|Grandparents|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|F|Black||45|28204|Some College|Married|Finance: Banking|29715|4|0|Big For A Day|Special Event|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502584168|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|4|||16422|8|||1|
502583660|503944507|500775919|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|589|Yellow||2014-09-15|2014-10-06|2016-05-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.4||2|2|1|1|F|Black||14|No|GrandMother|28215|Grandparents|$30,000 to $34,999|||Y|Yes||School|General Community||RTBM|F|White||35|28205|Masters Degree|Single|Education: Teacher|28273|3|6|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|502584168|31|0|2|1|0|2|7|2|500003586||4|2||-2|500000294|-2|0|4|||46|2|||1|
502583660|503286709|500701403|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|365|Red||2013-06-20|2013-06-26|2014-06-26|Volunteer: Time constraint|Volunteer: Time constraint||12||2|2|1|1|F|Black||14|No|GrandMother|28215|Grandparents|$30,000 to $34,999|||Y|Yes||School|General Community||RTBM|F|White||32|28211|Bachelors Degree|Single|Business|28211|3|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502584168|31|0|2|1|0|2|7|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
502320003|502810883|500606071|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|877|Red||2012-03-26|2012-04-30|2014-09-24|Volunteer: Moved|Volunteer: Moved||28.8||1|1|1|1|F|Black||14|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||30|28216||Single|Tech: Research/Design||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502320438|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|6854|8|||7464|9|||1|
502681380|502847991|500603939|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1002|Green||2012-03-14|2012-03-21|2014-12-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||32.9||1|1|1|1|M|White||14|No|Mother|28075|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|M|White||29|28277|Bachelors Degree|Single|Insurance|28262|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502682208|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
502236255|502436546|500518376|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1375|Red||2011-02-17|2011-02-24|2014-11-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||45.2||1|1|1|1|M|Black||14|No|Father|28214|Two Parent|Unknown||||Yes||Relative|General Community||Match Support|M|White||64|28207|Masters Degree|Married|Education: Teacher||0|0|Radio|Media|Big|General Site|mentor2.0 2015|Enrollment|0|1|1|0|277|60|598|500000170|500013781|502236686|31|0|1|1|0|1|10|2|-2||4|3||-2|500015184|-1|0|3|||131|1|||1|
502278985|500220237|500599107|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1841|Green|Project Big|2012-02-17|2012-03-01|NaT||||60.5||1|1|2|2|M|Black||14|No|Mother|28213|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||40|28269||Married|Business: Marketing||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|502279417|31|0|1|31|0|1|10|2|-2||2|1||-2|500000294|-2|6854|8|||2238|7|||1|500004640
503552606|501052547|500794702|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|846|Green||2014-11-12|2014-11-21|NaT||||27.8||1|1|2|2|M|Black||14|No|Mother|28079|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||45|28079|Bachelors Degree|Married|Business||13|6|Other|BBBS Board/Staff|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|503554481|31|0|1|31|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7671|13|||1|
503755565|503814505|500763994|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|434|Yellow||2014-05-21|2014-05-29|2015-08-06|Volunteer: Time constraint|Volunteer: Time constraint||14.3||1|1|1|1|M|Black||13|No|Mother|28227|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Enrollment|M|White||55|28031|Bachelors Degree|Separated|Business: Sales|53964|3|3|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|503757537|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7439|1|||1|
503632799|503567146|500763613|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1020|Green||2014-05-16|2014-05-31|NaT||||33.5||1|1|1|1|F|Black||13|No|Mother|28269|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||59|28209|Bachelors Degree|Divorced|Medical|28209|1|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503634738|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501332660|503579743|500715179|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|531|Green||2013-10-02|2013-10-24|2015-04-08|Volunteer: Moved|Volunteer: Moved||17.4||2|2|1|1|M|Black||13||GrandMother|28213|Grandparents|Unknown||||Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||42|28212|Bachelors Degree|Married|Arts, Entertainment, Sports|28202|2|11|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500011349|501332937|31|0|1|31|0|1|10|2|-2||4|1|500000294|-2||-2|6854|8|||7464|9|||1|
502605331|503090281|500627504|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1676|Red|Cabarrus County|2012-08-06|2012-08-13|NaT||||55.1||1|1|1|1|M|Hispanic||13|No|Mother|28027|One Parent: Female|$25,000 to $29,999||||No|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|White||33|28036|Bachelors Degree|Married|Business||2|5|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502605848|3|0|1|1|0|1|10|2|500016307||2|3|500016374|-2|500016374|-2|34|2|||7464|9|||1|500016374
501561525|501627716|500371266|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|443|Yellow||2009-06-26|2009-07-06|2010-09-22|Volunteer: Moved|Volunteer: Moved||14.6||1|1|1|1|M|Black||13|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|M|White||31|28202|||Consultant|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501561821|31|0|1|1|0|1|7|2|||4|2||-2||-2|0|10|||7464|9|||1|
501252806|501320197|500310204|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3033|Green||2008-11-04|2008-11-25|NaT||||99.6||1|1|1|1|M|Black||13|No|Mother|28078|One Parent: Female|Unknown||||No||Relative|General Community||Match Support|M|Black||45|28262|Bachelors Degree|Married|Business: Mgt, Admin||0|6|AA Task Force|Other Big|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501253082|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|3|||6247|12|||1|
503617980|503573243|500730441|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|772|Green||2013-11-13|2013-11-25|2016-01-06|Child/Family: Moved|Child/Family: Moved||25.4||1|1|1|1|F|Black||13|No|Mother|28217|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||25|28134|Some College|Single|Child/Day Care Worker||0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503619857|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
501445192|501508141|500343010|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|593|Green|Amachi|2009-02-19|2009-03-12|2010-10-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||19.5||1|1|1|1|M|Black||13|Yes|Mother|28202|One Parent: Female|Unknown||||Yes||Relative|General Community|Amachi|Match Support|M|Black||35|28212|Some College|Single|Finance: Banking|28204|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501445477|31|0|1|31|0|1|10|2|500003586||4|1|500000294|-2||-2|0|3|||7464|9|||1|500000294
502083465|502591360|500557052|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|609|Green||2011-09-22|2011-10-06|2013-06-06|Child/Family: Moved|Child/Family: Moved||20||1|1|2|2|F|Black||13|No|Mother|28025|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||69|28027||Married|Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|1|0|277|60|598|500000170|500012459|502083880|31|0|2|31|0|2|10|2|-2||4|1||-2|500016374|-2|0|10|||7464|9|||1|
503421607|503520561|500711787|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1251|Green||2013-09-18|2013-09-26|2017-02-28|Child: Family structure changed|Child: Family structure changed||41.1||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28214|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|Black||49|28273|Associate Degree|Single|Finance: Accountant|28273|7|0|Agency Sponsored|Special Event|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|503423471|36|0|2|31|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||16426|8|||1|
502346286|502726270|500564990|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|207|Yellow|Project Big|2011-10-13|2011-10-31|2012-05-25|Volunteer: Moved|Volunteer: Moved||6.8||1|1|1|1|M|Black||13|No|Mother|28214|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community|Project Big|Match Support|M|Black||44|28202||Single|Unknown||0|0|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500001281|502346724|31|0|1|31|0|1|10|2|500004641||4|2|500004640|-2|500004640|-2|6854|8|||7464|9|||1|500004640
501314104|501170940|500315948|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3024|Yellow||2008-11-17|2008-12-04|NaT||||99.4||1|1|1|1|M|Black||13|No|Mother|28217|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||39|28134|Bachelors Degree|Single|Business: Mgt, Admin||6|0|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500008321|501314382|31|0|1|1|0|1|10|2|-2||2|2||-2||-2|0|10|||7464|9|||1|
501662033|500459674|500597964|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|747|Green||2012-02-13|2012-03-03|2014-03-20|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||24.5||2|2|4|4|F|Black||13|No|Mother|28215|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Enrollment|F|Black||38|28219||Single|Finance: Banking|28273|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011349|501090456|31|0|2|31|0|2|5|2|-2||4|1||-2|500000294|-2|0|10|||2238|7|||1|
501662033|503655814|500767861|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|253|Green||2014-06-26|2014-06-30|2015-03-10|Volunteer: Moved|Volunteer: Moved||8.3||2|2|1|1|F|Black||13|No|Mother|28215|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Enrollment|F|White||27|28203|Bachelors Degree|Single|Finance: Banking|28211|2|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500011349|501090456|31|0|2|1|0|2|5|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
503977573|504047655|500801295|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|336|Red|PERL 2014-2016|2014-12-04|2014-12-29|2015-11-30|Volunteer: Moved|Volunteer: Moved||11||2|2|1|1|F|Black||13|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||29|28277|Bachelors Degree|Single|Business: Clerical|28202|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503980164|31|0|2|31|0|2|10|2|-2||4|3||-2|500014681|-2|0|10|||17159|12|||1|500014681
503662377|503573326|500743531|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1124|Green||2014-01-17|2014-01-31|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||36.9||1|1|1|1|F|Black||13|No|Mother|28216|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|F|White||28|28031|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503664337|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503052850|503028888|500626321|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1628|Green||2012-07-26|2012-09-30|NaT||||53.5||1|1|1|1|F|Hispanic||13|No|Mother|28277|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||31|28210|Bachelors Degree|Single|Education: Teacher|29710|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503027860|3|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
503959684|503985328|500775400|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|409|Green||2014-09-11|2014-09-15|2015-10-29|Child/Family: Moved|Child/Family: Moved||13.4||1|1|1|1|F|Black||13|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||26|28207|Masters Degree||Finance: Accountant|28202|0|11|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503961693|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503535102|503882165|500774003|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|239|Yellow||2014-09-02|2014-09-17|2015-05-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.9||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|Black||26|28214|Bachelors Degree|Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503536977|36|0|2|31|0|2|5|2|-2||4|2||-2||-2|0|10|||46|2|||1|
501704180|501216868|500435681|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|369|Green||2010-02-18|2010-02-25|2011-03-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||12.1||1|1|3|3|M|Black||13|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||32|28078||Single|Education: Teacher||0|0|other|College Partner|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500002335|501704518|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7670|5|||1|
502528776|502588092|500539956|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|126|Yellow||2011-06-06|2011-06-16|2011-10-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.1||1|1|1|1|F|Hispanic||13|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes|Come Out and Play|Special Event|General Community||RTBM|F|Hispanic||27|28031|Some College|Divorced|Retail: Mgt|28117|4|9|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502529226|3|0|2|3|0|2|7|2|-2||4|2||-2||-2|2203|12|||46|2|||1|
502225262|500205341|500459723|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|14|Green||2010-07-01|2010-07-15|2010-07-29|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||0.5||2|2|3|4|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown|||Y|Yes|AARTF|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||48|28213|Masters Degree|Divorced|Finance: Economist|28202|13|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|502225693|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|6855|8|||46|2|||1|
502225262|502244560|500463849|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|933|Yellow|Amachi|2010-08-02|2010-08-10|2013-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||30.7||2|2|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown|||Y|Yes|AARTF|Neighbor/Friend|General Community|Amachi|Match Support|F|Black||33|28204|Bachelors Degree|Single|Education: Teacher||0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|502225693|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2|500000294|-2|6855|8|||7496|10|||1|500000294
503989203|504066226|500799476|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|822|Green|PERL 2014-2016|2014-11-26|2014-12-15|NaT||||27||1|1|1|1|M|White||13|No|Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|Yes||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|White||33|28203|Bachelors Degree|Single|Finance: Banking|28203|7|8|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|503991217|1|0|1|1|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|0|5|||17159|12|||1|500014681
503268271|502993922|500669147|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|965|Red||2012-12-12|2012-12-27|2015-08-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.7||1|1|1|1|F|Black||13|No|Mother|28226|One Parent: Female|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||40|28273|Some College|Married|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503270085|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|6854|8|||7496|10|3|3|1|
502868923|502832013|500591320|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1372|Green|Project Big|2012-01-12|2012-01-27|2015-10-30|Volunteer: Moved|Volunteer: Moved||45.1||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||||Yes||School|General Community|Project Big|Match Support|F|Black||28|28262|Bachelors Degree|Single|Finance: Banking||0|0|AA Task Force|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502870324|31|0|2|31|0|2|10|2|500004641||4|1|500004640|-2||-2|0|4|||11098|8|||1|500004640
502605248|503049689|500623109|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|569|Green||2012-07-06|2012-08-07|2014-02-27|Volunteer: Time constraint|Volunteer: Time constraint||18.7||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|Unknown||||Yes||Relative|General Community|Project Big|Enrollment|M|White||36|28205|Masters Degree|Single|Finance: Banking||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502137975|31|0|1|1|0|1|5|2|-2||4|1|500004640|-2||-2|0|3|||7496|10|||1|
501674143|501474438|500365029|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|307|Green|Amachi|2009-05-22|2009-06-03|2010-04-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.1||1|1|1|1|F|Black||13|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||29|28273|Bachelors Degree|Single|Child/Day Care Worker|28209|5|0|BBBS National Site|Web Link|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500010355|501674477|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||46|2|||1|500000294
501755470|502038804|500456645|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2451|Green||2010-06-14|2010-06-30|NaT||||80.5||2|2|2|2|F|Black||13|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||Match Support|F|Black||51|28269||Married|Finance: Auditor||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|501755813|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
501755470|501595590|500373938|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|233|Red||2009-07-14|2009-07-22|2010-03-12|Volunteer: Time constraint|Volunteer: Time constraint||7.7||2|2|1|1|F|Black||13|No|GrandMother|28269|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||Match Support|F|White||30|28214|||Retail: Sales|28273|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501755813|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503328946|503371779|500703253|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1117|Green||2013-07-10|2013-07-19|2016-08-09|Volunteer: Moved|Volunteer: Moved||36.7||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Enrollment|M|Black||26|28217|Bachelors Degree|Single|Business: Marketing|28217|4|0|Coworker|Workplace Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503330792|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|10|||7447|3|||1|
501614593|500896567|500358150|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|350|Green||2009-04-20|2009-04-28|2010-04-13|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||11.5||1|1|2|2|M|Black||13|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|Black||68|28215||Married|Retired||0|0|Other Church Partner|Faith Organization|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500008629|501614913|31|0|1|31|0|1|5|2|-2||4|1||-2|500000294|-2|0|10|||7453|7|||1|
501319029|501130547|500306707|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|860|Green|Amachi|2008-10-28|2008-11-21|2011-03-31|Volunteer: Moved|Volunteer: Moved||28.3||4|4|2|2|F|Black||13|Yes|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||33|28202|Bachelors Degree|Single|Medical: Admin||0|9|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500003657|500948399|31|0|2|1|0|2|5|2|500003586||4|1|500014681|-2||-2|0|10|||46|2|||1|500000294
501319029|502425995|500534754|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|370|Red|Amachi|2011-05-03|2011-05-27|2012-05-31|Volunteer: Moved|Volunteer: Moved||12.2||4|4|1|1|F|Black||13|Yes|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||28|28203|Bachelors Degree|Single|Business: Sales|10595|0|8|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|500948399|31|0|2|1|0|2|5|2|500003586||4|3|500014681|-2||-2|0|10|||7464|9|||1|500000294
501319029|503078205|500673752|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1222|Red||2013-01-09|2013-01-31|2016-06-06|Volunteer: Moved|Volunteer: Moved||40.1||4|4|1|1|F|Black||13|Yes|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||28|28212|Bachelors Degree|Married|Child/Day Care Worker||0|3|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|500948399|31|0|2|1|0|2|5|2|-2||4|3|500014681|-2||-2|0|10|||7439|1|||1|
502866083|503378884|500688846|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1451|Green||2013-03-19|2013-03-26|NaT||||47.7||1|1|1|1|M|White||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||32|28104|Bachelors Degree|Single|Business|20785|0|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502867478|1|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502866079|503378886|500686789|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1451|Green||2013-03-08|2013-03-26|NaT||||47.7||1|1|1|1|M|White||13|No|Mother|28213|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|White||32|28210|Bachelors Degree|Single|Business: Sales||4|6|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020752|502867478|1|0|1|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
502477677|502621765|500545314|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|755|Red||2011-07-13|2011-07-29|2013-08-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.8||1|1|1|1|M|Black||13|No|Mother|28273|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|Black||31|28217|Bachelors Degree|Single|Business: Engineer|28273|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|502478124|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|5|||7496|10|||1|
501722052|502030533|500450450|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1725|Green|Amachi|2010-04-29|2010-05-11|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||56.7||2|2|1|1|F|White||13|Yes|GrandMother|28083|Grandparents|Unknown||||No||Self|General Community||Enrollment|F|White||40|28027||Single|Customer Service|28027|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|501227925|1|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|12|3|1|500000294
501722052|501737001|500363616|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|58|Green||2009-05-13|2009-05-18|2009-07-15|Volunteer: Health|Volunteer: Health||1.9||2|2|1|1|F|White||13|Yes|GrandMother|28083|Grandparents|Unknown||||No||Self|General Community||Enrollment|F|White||33|28078||Single|Business: Mgt, Admin||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501227925|1|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502435258|502670193|500589905|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1022|Green||2012-01-05|2012-01-12|2014-10-30|Volunteer: Time constraint|Volunteer: Time constraint||33.6||2|2|1|1|F|Black||13|No|Relative: Other|28081|Other Relative|Unknown|||Y|Yes||Self|General Community||Enrollment|F|Black||31|28025|Bachelors Degree|Single|Child/Day Care Worker|28027|5|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502435701|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
502435258|502449877|500520542|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|295|Green||2011-02-28|2011-03-16|2012-01-05|Volunteer: Moved|Volunteer: Moved||9.7||2|2|1|1|F|Black||13|No|Relative: Other|28081|Other Relative|Unknown|||Y|Yes||Self|General Community||Enrollment|F|White||30|28036||Single|Finance||0|0|Big Champions|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|502435701|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7461|12|||1|
501597169|501563612|500352827|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2612|Green||2009-03-26|2009-04-06|2016-05-31|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||85.8||1|1|1|1|M|Black||13||Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|Black||54|28262|High School Graduate|Married|Disabled||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|501597489|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503628199|503966130|500775002|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|169|Green||2014-09-09|2014-09-18|2015-03-06|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.6||1|1|1|1|M|Black||13|No|Mother|28273|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||54|28226|Masters Degree|Single|Tech: Computer/Programmer|28202|0|3|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|503630137|31|0|1|1|0|1|10|2|-2||4|1|500014681|-2|500000294|-2|0|10|||17159|12|||1|
501663584|501579777|500355189|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|179|Green||2009-04-03|2009-04-27|2009-10-23|Child/Family: Moved|Child/Family: Moved||5.9||1|1|1|1|M|White||13|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||32|28027|Bachelors Degree|Married|Finance: Banking||0|6|Recruitment Event|Workplace Partner|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500001262|501663922|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7446|3|||1|
503880559|503860995|500768591|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|43|Green||2014-07-03|2014-07-23|2014-09-04|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||1.4||1|1|2|2|F|Black||13|Yes|Father|28027|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Enrollment|F|Black||38|28269|Masters Degree|Single|Business|28262|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500002335|503882555|31|0|2|31|0|2|5|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|10|||46|2|||1|
502917069|502883342|500602923|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|272|Green||2012-03-08|2012-03-20|2012-12-17|Child/Family: Moved|Child/Family: Moved||8.9||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||29|28212|Masters Degree||Finance: Accountant||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008629|502918486|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|6854|8|||7464|9|||1|
502093515|502190908|500459974|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|567|Green|Amachi|2010-07-06|2010-07-13|2012-01-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.6||1|1|1|1|F|Black||13|Yes|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Enrollment|F|White||30|28203|Bachelors Degree|Single|Education||0|2|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013709|502093897|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|34|2|||7464|9|||1|500000294
502728289|502339145|500565493|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1952|Green||2011-10-14|2011-11-04|2017-03-09|Child/Family: Moved|Child/Family: Moved||64.1||1|1|1|1|F|Hispanic||13|No|Mother|28278|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|F|White||32|28211||Married|Finance||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|502729186|3|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|0|3|||7496|10|||1|
502721278|502701096|500560499|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1982|Green|Amachi, Cabarrus County|2011-10-03|2011-10-12|NaT||||65.1||1|1|1|1|M|White||13|Yes|Mother|28025|One Parent: Female|Unknown||||Yes||School|General Community|Cabarrus County|Match Support|M|White||47|28025||Single|Tech: Support, Writing|28026|0|2|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|501938680|1|0|1|1|0|1|10|2|500003586||2|1|500016374|-2|500016374|-2|0|4|||7464|9|||1|500000294, 500016374
502700500|502824634|500589524|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1889|Green||2012-01-03|2012-01-13|NaT||||62.1||1|1|1|1|M|Black||13|No|Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||30|28202|Bachelors Degree|Single|Business: Sales|28212|0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502701345|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502551048|501472128|500554178|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1184|Yellow||2011-09-12|2011-10-19|2015-01-15|Volunteer: Moved|Volunteer: Moved||38.9||1|1|2|2|F|Hispanic||13|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Enrollment|F|Black||52|30080|Bachelors Degree|Single|Consultant|2451|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|502551498|3|0|2|31|0|2|5|2|-2||4|2||-2||-2|0|4|||7464|9|||1|
502912138|502881673|500610045|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|427|Red||2012-04-16|2012-04-27|2013-06-28|Volunteer: Moved|Volunteer: Moved||14||3|3|2|2|M|Black||13|No|Mother|28216|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||33|28078|Bachelors Degree|Single|Business: Marketing|28036|5|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502913549|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
502912138|503541787|500704406|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|112|Red||2013-07-23|2013-08-22|2013-12-12|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.7||3|3|1|1|M|Black||13|No|Mother|28216|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|Black||31|28262|Bachelors Degree|Single|Business|28025|5|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502913549|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
502912138|503857059|500767007|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|368|Red||2014-06-18|2014-06-20|2015-06-23|Volunteer: Time constraint|Volunteer: Time constraint||12.1||3|3|1|1|M|Black||13|No|Mother|28216|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||28|28209|Bachelors Degree|Single|Business|28278|2|2|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502913549|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|34|2|||46|2|||1|
502763968|502939016|500608284|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1592|Red||2012-04-05|2012-04-30|2016-09-08|Volunteer: Moved|Volunteer: Moved||52.3||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Enrollment|M|White||38|28206|Bachelors Degree|Divorced|Business: Mgt, Admin|28164|3|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502764880|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
502338766|502249870|500526448|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|168|Green|Amachi, Project Big, Project Big AND Amachi|2011-03-21|2011-03-31|2011-09-15|Volunteer: Time constraint|Volunteer: Time constraint||5.5||1|1|1|1|M|Black||13|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||School|General Community|Project Big AND Amachi|Enrollment|M|Some Other Race||38|28226|Bachelors Degree|Single|Real Estate: Realtor||5|0||Relative|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502339202|31|0|1|41|0|1|5|2|500004772||4|1|500004901|-2|500004640|-2|0|4|||0|11|||1|500000294, 500004640, 500004901
503915384|503995835|500787470|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|872|Green|PERL 2014-2016|2014-10-23|2014-10-26|NaT||||28.6||1|1|1|1|M|Black||13|No|Mother|28262|One Parent: Female|$20,000 to $24,999||||Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|Multi-race (Asian & White)||36|28203|Masters Degree|Married|Finance: Banking|20815|11|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500018851|503917391|31|0|1|37|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|34|2|||7464|9|||1|500014681
503879123|503889097|500766443|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|999|Green||2014-06-12|2014-06-21|NaT||||32.8||1|1|1|1|M|Black||13|No|Mother|28212|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||33|28202|Masters Degree|Single|Finance: Banking|28244|0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503881119|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1|
503688885|503606993|500738203|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1184|Green||2013-12-11|2013-12-18|NaT||||38.9||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||35|28204|Bachelors Degree|Single|Retail: Mgt|28273|1|10|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503690850|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
503898651|503494199|500773073|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|530|Red||2014-08-21|2014-09-17|2016-02-29|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.4||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||40|28056|Some College|Single|Real Estate: Realtor|28202|2|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503891857|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
501712048|502405439|500516322|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2214|Green|Amachi|2011-02-09|2011-02-22|NaT||||72.7||1|1|1|1|M|Black||13|Yes|Mother|28134|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|M|White||29|28273|Some College|Single|Govt: Mgmt/Admin|28208|2|0|Relative|Relative|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020752|501712386|31|0|1|1|0|1|10|2|500003586||2|1|500000294|-2|500000294|-2|0|10|||17161|11|||1|500000294
502597599|500747912|500540004|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|369|Green|Project Big|2011-06-06|2011-06-30|2012-07-03|Child/Family: Moved|Child/Family: Moved||12.1||1|1|1|1|F|Black||13||Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big, Project Big AND Amachi|Match Support|F|White||28|28202|Bachelors Degree|Single|Finance: Banking|28255|1|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502598113|31|0|2|1|0|2|10|2|500004641||4|1|500004640, 500004901|-2||-2|0|10|||7462|13|||1|500004640
501938014|501874077|500426161|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1181|Green||2010-01-12|2010-01-15|2013-04-10|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||38.8||1|1|1|1|M|White||13|No|Mother|28083|One Parent: Female|Unknown|||Y|Yes||School|General Community|Cabarrus County, PERL 2014-2016|RTBM|M|Hispanic||44|28081|Bachelors Degree|Single|Business: Mgt, Admin|28025|2|10|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002335|501938412|1|0|1|3|0|1|7|2|-2||4|1|500014681, 500016374|-2||-2|0|4|||7464|9|||1|
502353937|501672025|500487322|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2306|Green|Amachi, Project Big, Project Big AND Amachi|2010-10-28|2010-11-22|NaT||||75.8||1|1|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown|||Y|Yes||School|General Community|Amachi, Project Big, Project Big AND Amachi|Match Support|F|White||31|29605|Bachelors Degree|Single|Business: Human Resources|29615|1|0|Local TV|Media|Big|General Community|Project Big AND Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|502354375|31|0|2|1|0|2|10|2|500004772||2|1|500000294, 500004640, 500004901|-2|500004901|-2|0|4|||7438|1|||1|500000294, 500004640, 500004901
503723868|503940354|500779635|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|367|Red||2014-10-01|2014-10-13|2015-10-15|Volunteer: Moved|Volunteer: Moved||12.1||1|1|1|1|M|Black||13|Yes|Mother|28215|One Parent: Female|$10,000 to $14,999||||Yes||Self|General Community||Enrollment|M|Black||25|28205|Bachelors Degree|Single|Tech: Research/Design|28202|0|11|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503725860|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|0|10|||17159|12|||1|
503034234|503070689|500639279|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|779|Green||2012-09-27|2012-10-29|2014-12-17|Volunteer: Moved|Volunteer: Moved||25.6||1|1|1|1|M|Hispanic||13|No|Mother|28078|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Enrollment|M|White||30|28031|Bachelors Degree|Married|Finance|28036|4|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503035830|3|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502249189|502485458|500523907|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|2010|Green||2011-03-08|2011-03-23|2016-09-22|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||66||1|1|1|1|M|Black||13|No|Mother|28277|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||34|28262||Married|Finance|29715|6|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500017732|502249620|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|34|2|||7462|13|||1|
503405468|502944301|500699540|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|793|Yellow||2013-06-05|2013-07-30|2015-10-01|Volunteer: Time constraint|Volunteer: Time constraint||26.1||2|2|2|2|F|White||13|No|Father|28211|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|White||58|28277|High School Graduate|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503407325|1|0|2|1|0|2|10|2|-2||4|2|500014681|-2||-2|0|10|||7464|9|||1|
503743876|503908096|500769242|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|691|Green||2014-07-11|2014-09-10|2016-08-01|Child/Family: Moved|Child/Family: Moved||22.7||1|1|1|1|M|Black||13|No|Mother|28212|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Enrollment|M|White||44|28203|Masters Degree|Single|Finance|29715|10|0|Igniting Breakfast|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503261158|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||17266|8|||1|
503851354|503962684|500774775|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|396|Red||2014-09-08|2014-09-29|2015-10-30|Volunteer: Moved|Volunteer: Moved||13||1|1|1|1|M|Black||13|Yes|Mother|28227|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|White||34|28209|Masters Degree|Single|Finance: Accountant|28210|2|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|503853343|31|0|1|1|0|1|10|2|-2||4|3||-2|500000294|-2|0|10|||46|2|||1|
502217146|502209019|500464101|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|657|Red|Amachi|2010-08-04|2010-08-13|2012-05-31|Volunteer: Time constraint|Volunteer: Time constraint||21.6||1|1|1|1|F|Black||13|Yes|Mother|28213|One Parent: Female|Unknown||||Yes|A Child's Place|Service Organization|General Community||Match Support|F|Multi-Race (None of the above)||28|28216||Single|Student: College||0|0||Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501364150|31|0|2|7|0|2|10|2|500003586||4|3||-2||-2|7016|11|||0|11|||1|500000294
503506115|503552068|500718774|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1070|Red||2013-10-14|2013-10-23|2016-09-27|Child: Family structure changed|Child: Family structure changed||35.2||1|1|1|1|M|Black||13|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Asian||54|28211|Masters Degree|Married|Self-Employed, Entrepreneur|28211|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503507986|31|0|1|4|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501868355|502820280|500592823|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|136|Red||2012-01-20|2012-02-13|2012-06-28|Volunteer: Time constraint|Volunteer: Time constraint||4.5||1|1|1|1|M|Black||13|No|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Enrollment|M|White||37|28277|Bachelors Degree|Single|Finance|91311|1|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501868724|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
502987717|503559146|500753781|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|372|Green||2014-03-10|2014-03-19|2015-03-26|Child/Family: Moved|Child/Family: Moved||12.2||1|1|1|1|F|Black||13|No|Mother|28134|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||37|28209|Bachelors Degree|Divorced|Medical|28078|5|6|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|502989174|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
502296291|502277214|500475457|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1029|Green||2010-09-30|2010-10-21|2013-08-15|Volunteer: Moved|Volunteer: Moved||33.8||1|1|1|1|M|White||13|No|Mother|28270|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||34|28278||Married|Self-Employed, Entrepreneur||4|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502296723|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502939347|503598887|500748884|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|597|Green||2014-02-13|2014-02-25|2015-10-15|Child/Family: Moved|Child/Family: Moved||19.6||1|1|1|1|F|Black||13|No|Mother|28052|Two Parent|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||32|28202|Masters Degree|Single|Medical: Doctor, Provider|28204|0|11|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|502940773|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502997224|502939526|500613729|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1057|Green||2012-05-08|2012-05-21|2015-04-13|Volunteer: Time constraint|Volunteer: Time constraint||34.7||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||32|28210|Bachelors Degree|Married|Business: Human Resources|28269|0|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500011349|502998689|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502576641|502537061|500535114|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2122|Green||2011-05-05|2011-05-25|NaT||||69.7||1|1|1|1|F|Black||13|No|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community||Match Support|F|White||41|28207|Masters Degree|Married|Business: Marketing|28202|2|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502577144|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|
502471024|502685747|500552890|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1788|Green||2011-09-01|2011-09-09|2016-08-01|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||58.7|Y|1|1|1|1|M|Black||13|Yes|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||51|28205|Bachelors Degree|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502471471|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502073665|502183515|500458730|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|699|Yellow||2010-06-28|2010-07-16|2012-06-14|Volunteer: Time constraint|Volunteer: Time constraint||23||2|2|1|1|F|Black||13|No|Mother|29732|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|F|White||31|28203|Masters Degree|Single|Finance: Accountant||1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502074089|31|0|2|1|0|2|7|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502073665|503245956|500696434|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|989|Red||2013-05-10|2013-05-21|2016-02-04|Child/Family: Moved|Child/Family: Moved||32.5||2|2|1|1|F|Black||13|No|Mother|29732|One Parent: Female|Unknown||||Yes||Self|General Community||RTBM|F|White||31|28226|Bachelors Degree|Single|Medical: Healthcare Worker|28211|0|3|Self|Self|Big|General Community|Amachi|Enrollment|0|1|0|1|277|60|598|500000170|500013781|502074089|31|0|2|1|0|2|7|2|-2||4|3||-2|500000294|-2|0|10|||7464|9|||1|
501750647|501584134|500374039|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1424|Red||2009-07-15|2009-08-31|2013-07-25|Volunteer: Time constraint|Volunteer: Time constraint||46.8||2|2|1|1|F|Black||13|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Site||Match Support|F|White||31|28207||Single|Medical: Nurse|28054|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501750989|31|0|2|1|0|2|10|2|-2||4|3||-1||-2|0|10|||7464|9|||1|
502217873|502223367|500478268|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|944|Red||2010-10-08|2010-10-27|2013-05-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31||1|1|1|1|F|Hispanic||13|No|Mother|28273|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Black||28|28273|Bachelors Degree|Single|Medical: Healthcare Worker|28211|0|9|Other|BBBS Board/Staff|Big|General Site|Amachi, mentor2.0 2014, Project Big|Enrollment|0|1|1|0|277|60|598|500000170|500011746|502218304|3|0|2|31|0|2|5|2|-2||4|3||-2|500000294, 500004640, 500014506|-1|0|10|||7671|13|||1|
503833936|502489398|500776719|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|900|Green||2014-09-18|2014-09-28|NaT||||29.6||1|1|1|1|M|Multi-race (Asian & White)||13|No|Mother|28078|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||33|28078|Bachelors Degree|Married|Unemployed|28031|6|2|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503835915|37|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
504139056|503991266|500801765|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|828|Green||2014-12-05|2014-12-09|NaT||||27.2||1|1|1|1|F|Black||13|No|Mother|28217|One Parent: Female|Unknown|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||28|28105|Masters Degree|Married|Business: Mgt, Admin|28211|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|504094626|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|5|||17159|12|||1|
501687330|501733851|500373679|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|374|Yellow|Amachi|2009-07-13|2009-07-17|2010-07-26|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||12.3||1|1|2|2|M|Black||13|Yes|Mother|28262|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|M|Black||50|28078|||Service: Restaurant|28082|0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500010355|501687668|31|0|1|31|0|1|5|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
503063881|503125383|500656877|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|775|Yellow||2012-11-07|2012-11-30|2015-01-14|Volunteer: Moved|Volunteer: Moved||25.5||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||34|28202|Associate Degree|Single|Medical: Healthcare Worker||6|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503065564|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
503594290|503508074|500735488|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1157|Green||2013-12-02|2014-01-14|NaT||||38||1|1|1|1|M|Multi-Race (None of the above)||13|No|Mother|28134|Other Relative|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|Hispanic||26|28205|||Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503596167|7|0|1|3|0|1|10|2|-2||2|1||-2||-2|0|5|||7464|9|||1|
503770823|503850589|500762293|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|985|Green||2014-05-06|2014-05-15|2017-01-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||32.4||1|1|1|1|M|White||13|No|Mother|28211|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||27|28270|Bachelors Degree|Single|Education: Teacher Asst/Aid|28202|0|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503772799|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||46|2|||1|
503689574|503577882|500751079|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|720|Green||2014-02-25|2014-03-20|2016-03-09|Volunteer: Moved|Volunteer: Moved||23.7||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|Unknown|||Y|Yes||Therapist/Counselor|General Community||Enrollment|F|White||33|28210|PHD|Single|Business: Human Resources|28273|0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503691539|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|5|||7464|9|||1|
502884974|503036135|500621875|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|604|Yellow||2012-06-26|2012-07-09|2014-03-05|Volunteer: Time constraint|Volunteer: Time constraint||19.8||1|1|1|1|M|Black||13|Yes|Mother|28217|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||34|28203|Some College|Single|Business: Marketing|28208|1|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502875571|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2||-2|0|10|||7496|10|||1|
503700282|503874948|500771987|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|118|Green||2014-08-12|2014-08-27|2014-12-23|Volunteer: Time constraint|Volunteer: Time constraint||3.9||1|1|1|1|M|Black||13|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|M|Black||42|28214|Some College|Domestic Partner|Service: Restaurant|28208|8|6|Man Up Campaign|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018987|503702247|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|10|||17101|1|||1|
501821947|500353496|500378466|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1182|Red||2009-08-12|2009-08-25|2012-11-19|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||38.8||1|1|4|4|M|Black||13|No|Mother|28105|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||43|28173|Masters Degree|Married|Finance: Banking|28281|7|0|Community Engagement|Special Event|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500011746|501822302|31|0|1|31|0|1|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|10|||18809|8|||1|
501859854|502044100|500469954|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1813|Green|Amachi|2010-09-13|2010-09-29|2015-09-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||59.6||1|1|1|1|F|Black||13|Yes|Mother|28216|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||28|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501860227|31|0|2|31|0|2|10|2|500003586||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
503893808|503976460|500803592|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|312|Red||2014-12-11|2014-12-20|2015-10-28|Volunteer: Moved|Volunteer: Moved||10.3||2|2|1|1|M|Black||13|No|GrandMother|28208|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|Asian||27|28203|Bachelors Degree|Single|Finance: Accountant|28202|1|10|Recruitment Event|BBBS Board/Staff|Big|General Community|mentor2.0 2014|Match Support|0|1|0|1|277|60|598|500000170|500013745|503227914|31|0|1|4|0|1|10|2|-2||4|3||-2|500014506|-2|0|4|||7462|13|||1|
503163476|503119713|500663695|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1567|Green||2012-11-27|2012-11-30|NaT||||51.5||1|1|1|1|M|Black||13|No|Mother|28269|One Parent: Female|$30,000 to $34,999|Yes: Active|No||No||Self|General Community||Match Support|M|Black||32|28217|Masters Degree|Single|Consultant||0|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503165154|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
501582587|501624537|500361275|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|406|Red||2009-05-05|2009-05-13|2010-06-23|Volunteer: Moved|Volunteer: Moved||13.3||1|1|1|1|M|Black||13|Yes|Mother|28215|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|M|White||35|28213|||Finance: Accountant|28117|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501582907|31|0|1|1|0|1|5|2|-2||4|3|500000294|-2||-2|0|10|||7464|9|||1|
502206598|502255565|500465186|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|993|Red|Amachi|2010-08-10|2010-08-20|2013-05-09|Child/Family: Time constraints|Child/Family: Time constraints||32.6||1|1|1|1|M|Black||13|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Service Organization|General Community|Amachi|Match Support|M|Black||34|28208|Bachelors Degree|Single|Finance|28202|9|0|Self|Self|Big|General Site||RTBM|0|1|1|0|277|60|598|500000170|500008321|502207027|31|0|1|31|0|1|10|2|500003586||4|3|500000294|-2||-1|0|11|||7464|9|||1|500000294
502969236|502938930|500612989|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|473|Red||2012-05-02|2012-05-14|2013-08-30|Volunteer: Time constraint|Volunteer: Time constraint||15.5||2|2|1|1|F|Some Other Race||13||Mother|28277|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||34|28277|Bachelors Degree||Medical: Nurse||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502970672|41|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
502969236|503567563|500718760|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|637|Yellow||2013-10-14|2013-10-24|2015-07-23|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||20.9||2|2|1|1|F|Some Other Race||13||Mother|28277|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||30|29730|Bachelors Degree|Single|Finance: Accountant|28273|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|502970672|41|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502728419|502889543|500594026|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|563|Red||2012-01-26|2012-02-06|2013-08-22|Volunteer: Time constraint|Volunteer: Time constraint||18.5||2|2|1|1|M|Black||13|No|Mother|28214|One Parent: Female|$50,000 to $59,999||||No|Big|Neighbor/Friend|General Community|PERL 2014-2016|Match Support|M|White||50|28105|Bachelors Degree|Married|Finance|28217|12|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502729316|31|0|1|1|0|1|10|2|-2||4|3|500014681|-2||-2|6854|8|||7496|10|||1|
502728419|504011804|500802308|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|822|Green|PERL 2014-2016|2014-12-09|2014-12-15|NaT||||27||2|2|1|1|M|Black||13|No|Mother|28214|One Parent: Female|$50,000 to $59,999||||No|Big|Neighbor/Friend|General Community|PERL 2014-2016|Match Support|M|White||25|28202|Bachelors Degree|Single|Tech: Computer/Programmer|28244|2|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|502729316|31|0|1|1|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|6854|8|||17159|12|||1|500014681
502207427|502236275|500464528|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|249|Yellow||2010-08-06|2010-08-15|2011-04-21|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||8.2||1|1|2|2|F|Black||13|No|Mother|28211|One Parent: Female|Unknown||||Yes||Service Organization|General Community||Match Support|F|White||39|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28217|1|7|Radio|Media|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500011639|502207856|31|0|2|1|0|2|10|2|-2||4|2||-2|500000294|-2|0|11|||131|1|||1|
502861545|501631588|500598474|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|242|Red||2012-02-15|2012-03-12|2012-11-09|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||8||1|1|3|3|M|Black||13|No|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Black||31|28203|Juris Doctorate (JD)||Law: Lawyer|28203|1|0|Self|Self|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500011349|502862935|31|0|1|31|0|1|10|2|-2||4|3||-2|500015184|-1|0|4|||7464|9|||1|
502720815|502647072|500566063|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|174|Red||2011-10-17|2011-11-30|2012-05-22|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.7||1|1|1|1|F|Black||13|No|Mother|28205|One Parent: Female|$15,000 to $19,999||||Yes|Big|Neighbor/Friend|General Community||RTBM|F|Black||40|28215|Some College|Single|Medical: Admin||11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502721710|31|0|2|31|0|2|7|2|-2||4|3||-2||-2|6854|8|||7462|13|||1|
502097794|502425119|500510881|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2247|Green||2011-01-13|2011-01-20|NaT||||73.8||1|1|1|1|M|Black||13|No|Mother|28269|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28031|Bachelors Degree|Single|Business: Engineer|28036|0|8|BBBS National Site|Web Link|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020910|502098218|31|0|1|1|0|1|10|2|-2||2|1||-2|500000294, 500004640|-2|34|2|||46|2|||1|
502184849|502513782|500529308|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|525|Green||2011-04-04|2011-04-20|2012-09-26|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||17.2||2|2|1|1|M|Multi-race (Hispanic & White)||13|No|Mother|28211|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||50|28269|Some College|Single|Tech: Engineer|28262|6|2|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011746|502185278|35|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502184849|503145815|500658541|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1549|Green||2012-11-12|2012-12-18|NaT||||50.9||2|2|1|1|M|Multi-race (Hispanic & White)||13|No|Mother|28211|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||28|28210|Bachelors Degree|Single|Business: Marketing|28224|1|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502185278|35|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
502915950|502913149|500602723|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|528|Green||2012-03-07|2012-04-02|2013-09-12|Volunteer: Moved|Volunteer: Moved||17.3||1|1|1|1|F|White||13|No|Mother|28031|One Parent: Female|$15,000 to $19,999|||Y|No||Self|General Community||Match Support|F|White||34|28031|Masters Degree|Single|Education||3|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502917364|1|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7496|10|||1|
503071350|503421602|500705806|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|629|Red||2013-08-05|2013-08-22|2015-05-13|Volunteer: Time constraint|Volunteer: Time constraint||20.7||3|3|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||36|28210|Masters Degree|Divorced|Medical|28209|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503073009|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
503071350|502831401|500625571|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|363|Red|Amachi|2012-07-23|2012-07-27|2013-07-25|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||11.9||3|3|1|1|F|Black||13|Yes|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||27|28226||Single|Student: College||0|0||Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|503073009|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||0|11|||1|500000294
502248033|502841432|500591252|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|535|Red||2012-01-12|2012-02-06|2013-07-25|Volunteer: Moved|Volunteer: Moved||17.6||1|1|1|1|M|Black||13|No|Mother|28273|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||28|28277|Bachelors Degree|Single|Business: Marketing||0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502248464|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||7496|10|||1|
501676480|501599611|500373737|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|276|Green||2009-07-13|2009-07-28|2010-04-30|Volunteer: Moved|Volunteer: Moved||9.1||1|1|1|1|M|Black||13|No|Mother|28214|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|White||31|28202|Bachelors Degree|Single|Finance: Banking||0|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501676818|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502261100|502284382|500512216|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2242|Green||2011-01-20|2011-01-25|NaT||||73.7||1|1|1|1|F|Black||13|No|Mother|28214|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|F|White||35|28209|Bachelors Degree|Single|Retail: Sales||6|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502261532|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|3|||7464|9|||1|
503029036|503070963|500626277|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|552|Green||2012-07-26|2012-08-07|2014-02-10|Volunteer: Moved|Volunteer: Moved||18.1||1|1|1|1|M|Black||13|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Enrollment|M|Asian||33|30097|Bachelors Degree|Single|Business|28255|5|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500002334|503030631|31|0|1|4|0|1|5|2|-2||4|1||-2||-2|0|5|||7464|9|||1|
502252822|502282155|500472826|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1232|Green||2010-09-23|2010-10-11|2014-02-24|Volunteer: Time constraint|Volunteer: Time constraint||40.5||3|3|1|1|F|Black||13|No|GrandMother|28227|Grandparents|Unknown||||No||Self|General Community||Match Support|F|White||34|28270||Single|Personal Trainer/Coach||10|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502253254|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502252822|503769635|500764054|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|203|Green||2014-05-21|2014-06-10|2014-12-30|Volunteer: Moved|Volunteer: Moved||6.7||3|3|1|1|F|Black||13|No|GrandMother|28227|Grandparents|Unknown||||No||Self|General Community||Match Support|F|Asian||26|28209|Bachelors Degree|Single|Business|28203|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502253254|31|0|2|4|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501781969|501902806|500418163|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|841|Yellow||2009-12-03|2009-12-10|2012-03-30|Volunteer: Moved|Volunteer: Moved||27.6||1|1|1|1|M|Black||13|No|Mother|28205|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||36|28205||Married|Law: Lawyer||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501745023|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502083438|502657267|500595491|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1869|Green|Cabarrus County|2012-02-01|2012-02-02|NaT||||61.4||1|1|1|1|F|Black||13|No|Mother|28083|One Parent: Female|Unknown||||Yes||Self|General Community|Cabarrus County|Match Support|F|Black||31|28269|Bachelors Degree|Single|Education: Teacher||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502083853|31|0|2|31|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7496|10|||1|500016374
501853851|502922901|500608304|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1268|Green|Amachi|2012-04-05|2012-04-30|2015-10-20|Child/Family: Moved|Child/Family: Moved||41.7||2|2|1|1|M|Black||13|Yes|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||55|28105|Masters Degree|Married|Law: Lawyer||25|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|501854219|31|0|1|1|0|1|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|500000294
501853851|501874309|500418151|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|627|Yellow|Amachi|2009-12-03|2009-12-14|2011-09-02|Volunteer: Time constraint|Volunteer: Time constraint||20.6||2|2|1|1|M|Black||13|Yes|Mother|28210|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||42|28207||Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|501854219|31|0|1|1|0|1|10|2|500003586||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
502089169|501875977|500452646|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|728|Red||2010-05-13|2010-05-27|2012-05-24|Volunteer: Moved|Volunteer: Moved||23.9||1|1|1|1|F|Black||13|No|Mother|28269|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|White||27|28213||Single|Human Services|28213|1|1|TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502089593|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|10|||130|1|||1|
501814187|500189590|500454641|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|819|Red|Amachi|2010-05-27|2010-06-03|2012-08-30|Volunteer: Time constraint|Volunteer: Time constraint||26.9||1|1|5|5|M|Black||13|Yes|Mother|28226|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|Some Other Race||46|28134|Bachelors Degree|Separated|Unknown||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|501814542|31|0|1|41|0|1|10|2|500003586||4|3|500000294|-2||-2|0|10|||2238|7|||1|500000294
501952951|502166996|500457775|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|432|Green||2010-06-22|2010-06-24|2011-08-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||14.2||1|1|3|3|M|Black||13||Mother|28210|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|Black||56|28277|Bachelors Degree|Married|Business||0|0|Michael Baisden|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501953349|31|0|1|31|0|1|5|2|-2||4|1||-2||-2|0|10|||11272|1|||1|
502619306|502716664|500565374|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1152|Green||2011-10-13|2011-10-22|2014-12-17|Volunteer: Time constraint|Volunteer: Time constraint||37.8||1|1|2|2|F|Hispanic||13|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|White||35|28205|Masters Degree|Married|Education: Teacher|28205|0|1|Recruitment Event|BBBS Board/Staff|Big|General Site|mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500017777|502619917|3|0|2|1|0|2|5|2|-2||4|1||-2|500015184|-1|0|10|||7462|13|||1|
501553422|501564519|500415759|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|235|Green|Amachi|2009-11-25|2009-12-17|2010-08-09|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||7.7||4|4|2|2|F|Black||13|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|F|Black||37|28269|Masters Degree|Single|Human Services: Social Worker|28212|0|6|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500003657|501536657|31|0|2|31|0|2|5|2|500003586||4|1|500000294|-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|500000294
501553422|501491899|500363856|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|110|Green||2009-05-14|2009-07-09|2009-10-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.6||4|4|1|1|F|Black||13|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|F|White||36|28270||Single|Business: Mgt, Admin|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|501536657|31|0|2|1|0|2|5|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|
501553422|502282024|500472224|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|239|Green|Amachi|2010-09-21|2010-09-28|2011-05-25|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||7.9||4|4|1|1|F|Black||13|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|F|White||33|28227|Bachelors Degree|Married|Medical: Nurse||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500003657|501536657|31|0|2|1|0|2|5|2|500003586||4|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|500000294
501553422|502646582|500548206|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1079|Red|Amachi|2011-08-01|2011-08-03|2014-07-17|Volunteer: Time constraint|Volunteer: Time constraint||35.4||4|4|1|1|F|Black||13|No|Mother|28227|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Enrollment|F|Black||31|28212|Masters Degree|Single|Human Services|28211|0|1|Sigma Gamma Rho|Fraternity/Sorority|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|501536657|31|0|2|31|0|2|5|2|500003586||4|3|500000294|-2||-2|0|10|||8700|14|||1|500000294
502882034|502983700|500615277|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1737|Green||2012-05-17|2012-06-13|NaT||||57.1||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Black||27|28208|Bachelors Degree|Single|Business: Mgt, Admin|28213|1|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|501390617|31|0|2|31|0|2|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1|
503584428|503839843|500761714|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1037|Green||2014-04-30|2014-05-14|NaT||||34.1||1|1|1|1|M|Black||13|No|Mother|28213|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|M|Black||27|28216|Some College|Single|Retail: Sales||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503586305|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503575828|503576000|500713280|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|445|Green||2013-09-25|2013-09-28|2014-12-17|Volunteer: Moved|Volunteer: Moved||14.6||3|3|1|1|M|Hispanic||13|No|Mother|28206|One Parent: Female|Unknown||||Yes|Spanish Radio|Media|General Community|PERL 2014-2016|Match Support|M|White||26|28203|Bachelors Degree|Single|Finance: Banking|28202|0|1|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017777|503577713|3|0|1|1|0|1|10|2|-2||4|1|500014681|-2|500000294|-2|7068|1|||7464|9|||1|
503663975|503854225|500762272|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|357|Red||2014-05-06|2014-05-22|2015-05-14|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||11.7||2|2|1|1|M|Black||13|Yes|Mother|28204|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|Black||33|28269|Bachelors Degree|Single|Insurance|28277|5|3|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503665933|31|0|1|31|0|1|10|2|-2||4|3|500000294|-2||-2|0|10|||17159|12|||1|
502634923|501197016|500548227|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1284|Green||2011-08-01|2011-08-16|2015-02-20|Child/Family: Moved|Child/Family: Moved||42.2||1|1|1|1|F|Black||13|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|F|Black||42|28210|Masters Degree|Single|Business: Clerical|28036|3|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502635617|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|3|||46|2|||1|
501573339|501835679|500384135|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|205|Green||2009-09-11|2009-09-30|2010-04-23|Volunteer: Moved|Volunteer: Moved||6.7||2|2|2|2|M|Black||13|No|Mother|28205|One Parent: Female|Unknown||||No||School|General Community||Enrollment|M|White||35|28226|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009242|501524605|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
501573339|501835679|500457932|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|972|Yellow||2010-06-23|2010-06-30|2013-02-26|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.9||2|2|2|2|M|Black||13|No|Mother|28205|One Parent: Female|Unknown||||No||School|General Community||Enrollment|M|White||35|28226|||Business: Sales||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501524605|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|4|||7464|9|||1|
503666549|504106972|500801599|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|826|Green|PERL 2014-2016, Cabarrus County|2014-12-05|2014-12-11|NaT||||27.1||1|1|1|1|M|Black||13|No|Mother|28025|One Parent: Female|$75,000 to $99,999||||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|M|Black||35|28027|Bachelors Degree|Married|Finance|28217|1|9|BBBS National Site|Web Link|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|503668509|31|0|1|31|0|1|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||46|2|||1|500014681, 500016374
503666553|503548907|500727074|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|321|Green||2013-11-04|2013-12-13|2014-10-30|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||10.5||2|2|1|1|F|Black||13|Yes|Mother|28025|One Parent: Female|$75,000 to $99,999||||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|Black||54|28056|PHD|Married|Education: College Professor|28017|4|0|Newspaper|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|503668509|31|0|2|31|0|2|10|2|-2||4|1|500014681, 500016374|-2||-2|0|10|||129|1|||1|
503666553|500991324|500801722|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|826|Green|PERL 2014-2016, Cabarrus County|2014-12-05|2014-12-11|NaT||||27.1||2|2|2|2|F|Black||13|Yes|Mother|28025|One Parent: Female|$75,000 to $99,999||||No||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||29|28027|Associate Degree|Single|Education||5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|503668509|31|0|2|1|0|2|10|2|500016307||2|1|500014681, 500016374|-2|500014681, 500016374|-2|0|10|||2238|7|||1|500014681, 500016374
503034769|503650997|500744436|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1140|Green||2014-01-23|2014-01-31|NaT||||37.5||1|1|1|1|M|Black||13|No|Mother|28226|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|Black||39|28210|Some College|Single|Arts, Entertainment, Sports|28202|7|2|Recruitment Event|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503036365|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7458|9|||1|
502242482|502214770|500466222|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|835|Yellow||2010-08-18|2010-09-10|2012-12-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27.4||1|1|1|1|F|Multi-race (Black & Hispanic)||13|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|White||55|28216|Some College|Divorced|Customer Service||16|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502242913|38|0|2|1|0|2|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503469072|503478672|500700143|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|596|Red||2013-06-10|2013-06-24|2015-02-10|Volunteer: Time constraint|Volunteer: Time constraint||19.6||2|2|1|1|M|White||13||GrandMother|28210|One Parent: Female|Unknown|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|White||35|28217||Married|Finance||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503470938|1|0|1|1|0|1|10|2|-2||4|3|500014681|-2||-2|0|10|||7464|9|||1|
502290605|500908500|500533937|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1130|Red|Amachi|2011-04-29|2011-05-09|2014-06-12|Volunteer: Moved|Volunteer: Moved||37.1||1|1|2|2|M|Black||13|Yes|Mother|28216|One Parent: Female|Unknown||||Yes|Radio|Media|General Community|Amachi|Enrollment|M|Black||48|28269||Divorced|Tech: Engineer||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502291037|31|0|1|31|0|1|5|2|-2||4|3|500000294|-2||-2|55|1|||7496|10|||1|500000294
502637766|503016558|500619500|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1657|Green||2012-06-15|2012-07-12|2017-01-24|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||54.4||1|1|1|1|M|Black||13|No|Mother|28262|One Parent: Female|$50,000 to $59,999||||Yes||School|General Community||Match Support|M|Black||34|28269|Juris Doctorate (JD)|Single|Law: Lawyer|28202|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|502638462|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|4|||7462|13|||1|
502582366|503858870|500766366|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|990|Green||2014-06-12|2014-06-30|NaT||||32.5||1|1|1|1|M|Black||13|No|Mother|28215|One Parent: Female|$45,000 to $49,999||||Yes||Self|General Community||Match Support|M|Black||31|28215|Some College|Single|Transport: Driver|28269|2|4|Local Radio|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502582874|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7437|1|||1|
503465438|503422939|500702504|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|458|Red||2013-07-01|2013-07-30|2014-10-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||15||1|1|1|1|F|Black||13|No|Mother|28215|One Parent: Female|$35,000 to $39,999||||Yes|BBBS National Site|Web Link|General Community||Enrollment|F|Some Other Race||31|28262|Masters Degree|Single|Finance: Accountant|28262|2|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503467304|31|0|2|41|0|2|5|2|-2||4|3||-2||-2|34|2|||7496|10|||1|
503710095|503872736|500766579|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1001|Green||2014-06-13|2014-06-19|NaT||||32.9||1|1|1|1|M|Black||13|No|Mother|28202|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||27|28202|Bachelors Degree|Single|Finance: Accountant|28226|0|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503712061|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1|
503496815|503673962|500739342|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|522|Red||2013-12-17|2014-01-13|2015-06-19|Volunteer: Time constraint|Volunteer: Time constraint||17.1||1|1|1|1|M|Black||13|No|Mother|28034|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||26|28217|Bachelors Degree|Single|Tech: Engineer|28217|0|3|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|503773736|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
503024102|502961739|500617100|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|264|Red||2012-05-30|2012-06-08|2013-02-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.7||2|2|1|1|F|Black||13|No|Mother|28227|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|Black||46|28270|Masters Degree|Single|Tech: Support, Writing|28204|10|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|501001116|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503024102|503465770|500700716|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|466|Red||2013-06-14|2013-06-21|2014-09-30|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||15.3||2|2|1|1|F|Black||13|No|Mother|28227|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||28|28212|Bachelors Degree|Single|Finance|28217|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|501001116|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502747706|502618438|500566066|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1422|Red||2011-10-17|2011-11-17|2015-10-09|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||46.7||1|1|1|1|F|Multi-Race (None of the above)||13|No|Mother|28229|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Enrollment|F|Black||34|28226|Bachelors Degree|Single|Business: Clerical|28208|0|6|Self|Self|Big|General Community|Project Big|Enrollment|0|1|0|1|277|60|598|500000170|500017777|502748616|7|0|2|31|0|2|5|2|-2||4|3||-2|500004640|-2|0|10|||7464|9|||1|
502275237|502264824|500470332|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|458|Yellow|Amachi|2010-09-14|2010-09-28|2011-12-30|Volunteer: Time constraint|Volunteer: Time constraint||15||1|1|1|1|M|Black||13|Yes|Mother|28262|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|M|Multi-Race (None of the above)||50|28027|Bachelors Degree|Married|Human Services: Non-Profit|28205|0|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500012459|502275669|31|0|1|7|0|1|5|2|-2||4|2|500000294|-2|500000294|-2|0|10|||7462|13|||1|500000294
501732944|501784291|500370063|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|998|Green||2009-06-18|2009-07-07|2012-03-31|Child/Family: Moved|Child/Family: Moved||32.8||1|1|1|1|F|Black||13|No|Mother|28262|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|American Indian or Alaska Native||34|28209|Masters Degree|Married|Human Services: Social Worker||0|10|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501733284|31|0|2|6|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
501858025|501664714|500449971|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|952|Red|Amachi, Project Big|2010-04-27|2010-05-14|2012-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||31.3||1|1|2|2|M|Black||13|Yes|Mother|28216|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, Project Big|Match Support|M|Black||44|28273|||Finance: Accountant||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|501858397|31|0|1|31|0|1|10|2|-2||4|3|500000294, 500004640|-2|500000294|-2|0|4|||7464|9|||1|500000294, 500004640
502873189|502882530|500600322|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1625|Yellow||2012-02-24|2012-03-21|2016-09-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||53.4||1|1|1|1|F|Black||13|No|Mother|28206|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Black||40|28216|Masters Degree|Single|Finance||6|0|Charlotte Cares|Service Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502874592|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|4|||11246|6|||1|
502207223|503251424|500703587|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1332|Green||2013-07-15|2013-07-23|NaT||||43.8||2|2|1|1|F|Black||13|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||38|28273|Bachelors Degree|Separated|Customer Service|28134|1|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502207652|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|6854|8|||7464|9|||1|
502207223|502226588|500461272|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|781|Yellow||2010-07-16|2010-07-26|2012-09-14|Volunteer: Time constraint|Volunteer: Time constraint||25.7||2|2|1|1|F|Black||13|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||31|28207|Bachelors Degree|Living w/ Significant Other|Unemployed|28205|3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502207652|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1|
503869451|503940385|500783066|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|64|Green||2014-10-13|2014-10-27|2014-12-30|Volunteer: Moved|Volunteer: Moved||2.1||2|2|1|1|F|White||13|No|Mother|28212|Two Parent|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Enrollment|F|White||30|28205|Masters Degree|Single|Business|28201|2|3|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503871445|1|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|5|||46|2|||1|
503552498|503538554|500744965|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1141|Green||2014-01-27|2014-01-30|NaT||||37.5||1|1|1|1|F|Black||13|No|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||29|28210|Bachelors Degree|Single|Business: Marketing|28277|1|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503554371|31|0|2|1|0|2|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1|
503774057|503665969|500762915|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1028|Green||2014-05-12|2014-05-23|NaT||||33.8||1|1|1|1|F|Multi-race (Black & Hispanic)||13|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|White||61|28211|Bachelors Degree|Divorced|Tech: Management|28202|2|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503776034|38|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503532014|503694720|500753716|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|474|Yellow||2014-03-10|2014-03-21|2015-07-08|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||15.6||2|2|2|2|M|White||12|No|Mother|28025|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community|Amachi, Cabarrus County|Match Support|M|White||58|28075|Masters Degree|Married|Business|32824|0|6|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500012459|503533889|1|0|1|1|0|1|10|2|-2||4|2|500000294, 500016374|-2|500007920, 500011315, 500011316, 500014681, 500016374|-2|0|10|||7464|9|||1|
502630684|502703214|500564807|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|320|Red|Amachi, Project Big AND Amachi|2011-10-13|2011-10-26|2012-09-10|Child: Severity of challenges|Child: Severity of challenges||10.5||1|1|1|1|M|Black||12|Yes|Mother|28214|One Parent: Female|$10,000 to $14,999|||Y|Yes||Therapist/Counselor|General Community||Enrollment|M|Black||31|28214|Bachelors Degree|Single|Finance: Banking|28208|0|4|Radio|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502631339|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|0|5|||131|1|||1|500000294, 500004901
503207102|503688236|500757797|BBBS of Greater Charlotte|Main Office|N|C|Inactive|Match Support|1070|Green||2014-04-01|2014-04-11|NaT||||35.2||1|1|1|1|M|Multi-race (Black & Hispanic)||12|No|Mother|28270|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|M|White||54|28110|Some College|Married|Self-Employed, Entrepreneur|28110|11|6|Relative|Relative|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|0|1|0|1|277|60|598|500000170|500017777|503208876|38|0|1|1|0|1|10|2|-2||3|1||-2|500011312|-2|0|10|||17161|11|||1|
501806165|501706064|500375643|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2779|Green|Amachi|2009-07-27|2009-08-06|NaT||||91.3||1|1|1|1|M|Black||12|Yes|GrandMother|28273|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|M|Black||40|28273|No High School|Single|Business: Human Resources||2|0|Recruitment Event|Workplace Partner|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501806520|31|0|1|31|0|1|10|2|-2||2|1|500000294|-2||-2|0|10|||7446|3|||1|500000294
502787404|503485414|500701279|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1359|Yellow||2013-06-19|2013-06-26|NaT||||44.6||1|1|1|1|M|Black||12|No|Mother|28227|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||32|28262|Some College|Single|Business||0|5|United Way|Service Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502788587|31|0|1|31|0|1|10|2|-2||2|2||-2||-2|0|10|||16263|6|||1|
502740493|502875462|500605781|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|475|Yellow||2012-03-22|2012-04-12|2013-07-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||15.6||1|1|1|1|M|Black||12|No|Mother|28214|One Parent: Female|$60,000 to $74,999||||Yes||Relative|General Community||Match Support|M|Black||45|28217|High School Graduate|Separated|Transport: Driver||0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|502741396|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|3|||7464|9|||1|
502431551|502367677|500515625|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|205|Yellow|Amachi|2011-02-04|2011-02-09|2011-09-02|Child/Family: Unrealistic expectations|Child/Family: Unrealistic expectations||6.7||1|1|2|2|F|Black||12|Yes|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Enrollment|F|Black||36|28208|Some College|Single|Education: Teacher|28226|1|0|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011184|502431994|31|0|2|31|0|2|5|2|500003586||4|2|500000294|-2|500000294, 500004640|-2|0|10|||7464|9|||1|500000294
501832800|502528373|500533462|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|566|Red||2011-04-26|2011-05-03|2012-11-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.6||2|2|1|1|M|Black||12|No|Mother|28213|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|Black||50|28213|Bachelors Degree|Married|Finance||0|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|501833168|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501832800|501895777|500407077|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|254|Red||2009-11-05|2009-11-08|2010-07-20|Volunteer: Moved|Volunteer: Moved||8.3||2|2|1|1|M|Black||12|No|Mother|28213|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|M|White||34|28210|Bachelors Degree|Single|Finance||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009007|501833168|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503995803|503963125|500790223|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|311|Red|PERL 2014-2016|2014-10-30|2014-11-24|2015-10-01|Volunteer: Time constraint|Volunteer: Time constraint||10.2||1|1|1|1|F|Black||12|No|Mother|28206|Two Parent|$10,000 to $14,999|||Y|Yes||Relative|General Community|PERL 2014-2016|Match Support|F|Black||44|28269||Single|Unemployed||0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|503997818|31|0|2|31|0|2|10|2|-2||4|3|500014681|-2|500014681|-2|0|3|||17159|12|||1|500014681
503547661|503731665|500742652|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|560|Green||2014-01-14|2014-01-23|2015-08-06|Child/Family: Moved|Child/Family: Moved||18.4||1|1|1|1|M|Black||12|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||41|28277|Bachelors Degree|Divorced|Business|28273|4|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503549536|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
502904444|502883475|500683493|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|595|Yellow||2013-02-21|2013-03-06|2014-10-22|Child: Family structure changed|Child: Family structure changed||19.5||1|1|1|1|M|Black||12|Yes|Mother|28278|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||36|29715|Bachelors Degree|Single|Tech: Research/Design|28226|0|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502905855|31|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502552445|502545537|500539524|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2104|Green|Project Big|2011-06-02|2011-06-12|NaT||||69.1||1|1|1|1|F|Black||12|No|GrandMother|28208|One Parent: Female|$15,000 to $19,999|||Y|Yes||School|General Community|Project Big|Match Support|F|White||28|28209|Bachelors Degree|Single|Business: Sales|28277|0|9|Self|Self|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020910|502552891|31|0|2|1|0|2|10|2|500004641||2|1|500004640|-2|500000294, 500004640|-2|0|4|||7464|9|||1|500004640
502278991|502263116|500494784|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2295|Green||2010-11-15|2010-12-03|NaT||||75.4||1|1|1|1|F|Black||12|No|Mother|28213|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|Black||40|28269|Bachelors Degree|Married|Tech: Management|28255|1|9|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|502279417|31|0|2|31|0|2|10|2|-2||2|1||-2|500000294|-2|6854|8|||6247|12|||1|
502979757|503161988|500682191|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1461|Red||2013-02-14|2013-02-28|2017-02-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||48||1|1|1|1|M|Black||12|No|Mother|28211|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||31|28210|Bachelors Degree|Single|Business: Engineer||5|0|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502981210|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||17161|11|||1|
502234905|502799047|500583119|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1359|Green|Amachi|2011-11-30|2011-12-05|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||44.6||3|3|1|1|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28083|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|M|White||36|28097|Masters Degree|Divorced|Finance|28026|7|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|502777258|38|0|1|1|0|1|10|2|-2||4|1|500000294, 500014681, 500016374|-2||-2|0|10|||7671|13|||1|500000294
502234905|502570625|500545380|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|133|Yellow|Amachi|2011-07-13|2011-07-20|2011-11-30|Volunteer: Time constraint|Volunteer: Time constraint||4.4||3|3|1|1|M|Multi-race (Black & Hispanic)||12|Yes|Mother|28083|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi, Cabarrus County, PERL 2014-2016|Match Support|M|White||32|28027|||Retail: Sales||0|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502777258|38|0|1|1|0|1|10|2|500003586||4|2|500000294, 500014681, 500016374|-2||-2|0|10|||7464|9|||1|500000294
502280287|502290873|500483592|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|785|Yellow|Project Big|2010-10-20|2010-10-28|2012-12-21|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25.8||1|1|1|1|M|Black||12|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|M|White||50|28105||Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500008321|502280719|31|0|1|1|0|1|10|2|-2||4|2|500004640|-2|500004640|-2|0|10|||7464|9|||1|500004640
502879621|502295287|500603216|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|912|Red||2012-03-09|2012-05-15|2014-11-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||30||1|1|2|2|F|Black||12|No|Mother|28269|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|F|White||47|28078|Juris Doctorate (JD)|Single|Law: Lawyer|28203|8|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502881024|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
503978153|504039547|500798168|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|822|Green|PERL 2014-2016|2014-11-21|2014-12-15|NaT||||27||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Black||37|28227|Associate Degree|Single|Student: College|28223|1|0|Web in a Box, v1|Web Link|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503980164|31|0|2|31|0|2|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||15467|2|||1|500014681
501955885|501863882|500420833|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|790|Green||2009-12-11|2009-12-30|2012-02-28|Child/Family: Moved|Child/Family: Moved||26||1|1|1|1|F|Black||12||Mother|28208|One Parent: Female|Unknown||||Yes||Relative|General Community||Match Support|F|Black||55|28216|||Customer Service||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501873510|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|3|||7464|9|||1|
502933371|503080292|500623322|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1707|Green||2012-07-09|2012-07-13|NaT||||56.1||2|2|1|1|M|Black||12|No|Mother|28206|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Site||Match Support|M|White||37|28209|Bachelors Degree|Married|Unemployed|22202|9|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502934793|31|0|1|1|0|1|10|2|-2||2|1||-1||-2|0|10|||7496|10|||1|
502173768|503831898|500784859|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|862|Red|PERL 2014-2016|2014-10-17|2014-10-20|2017-02-28|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||28.3||3|3|1|1|F|Black||12|Yes|Mother|28211|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|F|Black||58|28269|Bachelors Degree|Married|Self-Employed, Entrepreneur|28269|26|0|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503800801|31|0|2|31|0|2|10|2|-2||4|3|500000294, 500014681|-2|500014681|-2|0|4|||7464|9|||1|500014681
502173768|501454688|500453997|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|452|Yellow|Amachi|2010-05-24|2010-05-28|2011-08-23|Volunteer: Moved|Volunteer: Moved||14.9||3|3|2|2|F|Black||12|Yes|Mother|28211|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|F|White||35|28277|||Education: Teacher|28025|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|503800801|31|0|2|1|0|2|10|2|500003586||4|2|500000294, 500014681|-2||-2|0|4|||7464|9|||1|500000294
502173768|502653258|500557879|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|321|Green|Amachi|2011-09-26|2011-10-20|2012-09-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.5||3|3|1|1|F|Black||12|Yes|Mother|28211|One Parent: Female|Unknown||||Yes||School|General Community|Amachi, PERL 2014-2016|Match Support|F|Black||27|28277||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|503800801|31|0|2|31|0|2|10|2|-2||4|1|500000294, 500014681|-2||-2|0|4|||7464|9|||1|500000294
503636487|503899296|500778337|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|871|Green|PERL 2014-2016|2014-09-25|2014-10-27|NaT||||28.6||1|1|1|1|M|Black||12|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|White||27|28205|Bachelors Degree|Single|Finance: Accountant|28202|1|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500013781|503665377|31|0|1|1|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681
503590328|503874645|500771736|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|763|Red||2014-08-07|2014-08-27|2016-09-28|Volunteer: Time constraint|Volunteer: Time constraint||25.1||1|1|1|1|M|Hispanic||12|No|Mother|28277|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|M|Some Other Race||31|28270|Bachelors Degree|Married|Real Estate: Realtor|28110|0|5|Man Up Campaign|Media|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|0|1|0|1|277|60|598|500000170|500008321|503592205|3|0|1|41|0|1|10|2|-2||4|3||-2|500011312|-2|0|10|||17101|1|||1|
502249038|502254632|500466270|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|822|Red|Amachi|2010-08-19|2010-08-31|2012-11-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||27||1|1|1|1|F|Multi-race (Black & White)||12|Yes|GrandMother|28278|Grandparents|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|White||34|28217|Bachelors Degree|Single|Retail: Sales||2|6|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|502249469|36|0|2|1|0|2|10|2|-2||4|3|500000294|-2|500000294|-2|0|10|||7496|10|||1|500000294
502898016|502951132|500614703|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|505|Yellow||2012-05-14|2012-05-29|2013-10-16|Volunteer: Moved|Volunteer: Moved||16.6||1|1|1|1|F|Black||12|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|Black||25|28205||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502899424|31|0|2|31|0|2|5|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502223076|502226529|500461246|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|370|Green||2010-07-16|2010-07-23|2011-07-28|Volunteer: Time constraint|Volunteer: Time constraint||12.2||2|2|1|1|F|Black||12|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|Black||33|28212|Juris Doctorate (JD)|Single|Law: Lawyer|28212|1|2|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011184|502223507|31|0|2|31|0|2|10|2|-2||4|1|500004640|-2|500000294|-2|0|10|||7464|9|||1|
502223076|502694717|500560829|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1973|Green||2011-10-04|2011-10-21|NaT||||64.8||2|2|1|1|F|Black||12|No|Mother|28216|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|White||30|28205|Bachelors Degree|Single|Business: Mgt, Admin|28204|0|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502223507|31|0|2|1|0|2|10|2|-2||2|1|500004640|-2||-2|0|10|||7464|9|||1|
503895740|503765053|500768490|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|383|Yellow||2014-07-02|2014-08-28|2015-09-15|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12.6||2|2|1|1|F|Black||12|No|Mother|28273|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||34|28214|Some College|Single|Transport: Driver|28273|9|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|503897736|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
501731844|501599513|500374438|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|334|Green|Amachi|2009-07-17|2009-08-07|2010-07-07|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||11||2|2|1|1|F|Black||12|Yes|Father|28210|One Parent: Male|Unknown||||Yes||Self|General Community||Enrollment|F|Black||42|28277|||Law: Police Officer|28202|0|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500003657|501732181|31|0|2|31|0|2|5|2|500003586||4|1||-2||-2|0|10|||7464|9|||1|500000294
501731844|501945149|500478465|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|620|Yellow|Amachi|2010-10-08|2010-10-19|2012-06-30|Volunteer: Moved|Volunteer: Moved||20.4||2|2|1|1|F|Black||12|Yes|Father|28210|One Parent: Male|Unknown||||Yes||Self|General Community||Enrollment|F|Black||36|28273|Associate Degree|Single|Business: Mgt, Admin|28255|0|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500013709|501732181|31|0|2|31|0|2|5|2|-2||4|2||-2|500000294|-2|0|10|||46|2|||1|500000294
502761742|503041890|500699565|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1357|Green|Cabarrus County|2013-06-05|2013-06-28|NaT||||44.6||1|1|2|2|M|Black||12|No|Mother|28083|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||60|28027|Bachelors Degree|Separated|Insurance|28262|24|0|Local Radio|Media|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502762654|31|0|1|1|0|1|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7437|1|||1|500016374
503047019|503070946|500655762|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|468|Red||2012-11-05|2012-11-16|2014-02-27|Volunteer: Time constraint|Volunteer: Time constraint||15.4||1|1|1|1|F|Hispanic||12|No|Mother|28211|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Hispanic||31|28210|Masters Degree|Single|Business||1|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|503048667|3|0|2|3|0|2|10|2|-2||4|3||-2||-2|0|10|||7496|10|||1|
503512877|503893014|500766726|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|853|Green||2014-06-16|2014-07-11|2016-11-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28||1|1|1|1|M|Black||12|No|Mother|28211|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|M|White||27|28226|Bachelors Degree|Single|Tech: Research/Design|28269|0|8|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|503514748|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||17101|1|||1|
502614388|502617891|500547414|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|363|Yellow|Amachi|2011-07-25|2011-09-13|2012-09-10|Volunteer: Moved|Volunteer: Moved||11.9||1|1|1|1|F|Black||12|Yes|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|White||30|28209||Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|502615000|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|5|||7496|10|||1|500000294
504038458|503971368|500800323|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|821|Green||2014-12-02|2014-12-16|NaT||||27||1|1|1|1|F|Black||12|No|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||25|28209|Bachelors Degree|Single|Finance|28202|1|3|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020752|504040320|31|0|2|1|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||17159|12|||1|
501314348|502205797|500460633|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1801|Red||2010-07-12|2010-08-25|2015-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||59.2||1|1|1|1|M|Black||12|No|Mother|28210|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||45|28211|Masters Degree|Married|Finance: Banking||11|0|Friendship Missionar|Faith Organization|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|501314626|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||2230|7|||1|
503565123|503673127|500739078|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|39|Green||2013-12-16|2014-01-23|2014-03-03|Volunteer: Moved|Volunteer: Moved||1.3||1|1|1|1|M|Black||12|No|Mother|28213|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|White||30|28262|Masters Degree|Single|Tech: Engineer|28078|2|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503566998|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503701025|503576358|500731543|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|997|Green||2013-11-15|2013-11-25|2016-08-18|Volunteer: Time constraint|Volunteer: Time constraint||32.8||1|1|1|1|F|Black||12|Yes|Mother|28269|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|White||53|28227|Some College|Married|Customer Service|28105|30|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|501153063|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502090492|503088662|500631918|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|378|Red||2012-09-04|2012-09-13|2013-09-26|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||12.4||1|1|1|1|M|Black||12|No|Mother|28215|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||44|28213|Associate Degree|Single|Laborer|28216|4|6|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502090916|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|0|10|||7438|1|||1|
502280689|502592849|500541235|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|212|Red||2011-06-15|2011-06-28|2012-01-26|Child/Family: Moved|Child/Family: Moved||7||1|1|1|1|M|Black||12|No|Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Enrollment|M|Some Other Race||38|28202|Bachelors Degree|Single|Business: Mgt, Admin||0|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502281121|31|0|1|41|0|1|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502789637|502883706|500604101|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|411|Yellow||2012-03-14|2012-03-29|2013-05-14|Volunteer: Time constraint|Volunteer: Time constraint||13.5||4|4|1|1|F|Black||12|No|Mother|28081|One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|White||51|28025|Some College|Divorced|Medical: Admin|28211|28|4|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502790820|31|0|2|1|0|2|10|2|-2||4|2|500016374|-2||-2|0|4|||7496|10|||1|
502789637|503542037|500708902|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|701|Yellow||2013-09-03|2013-09-23|2015-08-25|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||23||4|4|2|2|F|Black||12|No|Mother|28081|One Parent: Female|Less than $10,000||||Yes||School|General Community|Cabarrus County|Match Support|F|Black||30|28027|Masters Degree|Married|Unemployed|28027|2|5|Self|Self|Big|General Community|Cabarrus County, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500012459|502790820|31|0|2|31|0|2|10|2|-2||4|2|500016374|-2|500007920, 500011315, 500011316, 500016374|-2|0|4|||7464|9|||1|
503355095|503373533|500691042|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1102|Green||2013-04-02|2013-04-26|2016-05-02|Volunteer: Time constraint|Volunteer: Time constraint||36.2||1|1|1|1|F|Black||12|Yes|Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||36|28210|Juris Doctorate (JD)|Single|Law: Lawyer|28202|5|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503356940|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2||-2|0|10|||7496|10|||1|
503401214|503758808|500752693|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1086|Yellow||2014-03-04|2014-03-26|NaT||||35.7||1|1|1|1|M|Black||12|No|Mother|28105|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||31|28226|Bachelors Degree|Single|Finance: Accountant|28217|4|11|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503403071|31|0|1|1|0|1|10|2|-2||2|2||-2||-2|0|10|||7496|10|||1|
503011520|502970448|500617581|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|171|Yellow||2012-06-01|2012-07-05|2012-12-23|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||5.6||1|1|1|1|F|Black||12|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||41|28273|Bachelors Degree|Married|Business: Human Resources|28209|9|9|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503013050|31|0|2|1|0|2|10|2|-2||4|2|500000294|-2||-2|0|10|||7464|9|||1|
502234486|500189813|500462432|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|732|Red|Project Big|2010-07-23|2010-07-30|2012-07-31|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||24||2|2|2|2|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||School|General Site|Project Big|Match Support|F|Black||39|28278|Bachelors Degree|Single|Finance: Accountant|28217|0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|502234907|31|0|2|31|0|2|10|2|500004641||4|3|500004640|-1|500000294|-2|0|4|||2238|7|||1|500004640
502245343|502526001|500532810|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2142|Green|Amachi|2011-04-21|2011-05-05|NaT||||70.4||1|1|1|1|M|Black||12|Yes|Mother|28216|One Parent: Female|Unknown||||No||Self|General Community|Amachi|Match Support|M|White||32|28104|Bachelors Degree|Single|Business|28216|5|3|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502245774|31|0|1|1|0|1|10|2|500003586||2|1|500000294|-2||-2|0|10|||17161|11|||1|500000294
503782875|503732680|500763995|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|160|Green||2014-05-21|2014-05-30|2014-11-06|Agency: Challenges with program/partnership|Agency: Challenges with program/partnership||5.3||1|1|1|1|F|Black||12|No|Mother|28227|Two Parent|$40,000 to $44,999||||No|BBBS National Site|Web Link|General Community||Match Support|F|White||22|28206|Some College|Single|Child/Day Care Worker||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|503784852|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
503472232|503444888|500700046|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1148|Red||2013-06-10|2013-06-17|2016-08-08|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||37.7||1|1|1|1|M|Black||12||Mother|28217|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||48|28273|Some College|Divorced|Transport: Driver|29730|3|0|TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503474098|31|0|1|31|0|1|10|2|-2||4|3||-2||-2|34|2|||130|1|||1|
502347820|502419409|500588112|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1511|Yellow|Amachi|2011-12-20|2011-12-20|2016-02-08|Volunteer: Moved|Volunteer: Moved||49.6||3|3|2|2|F|Black||12|Yes|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Some Other Race||75|28213|Some College|Widowed|Human Services||20|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020990|502348258|31|0|2|41|0|2|10|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
502347820|502419409|500520174|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|14|Green||2011-02-25|2011-03-16|2011-03-30|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||0.5||3|3|2|2|F|Black||12|Yes|Mother|28227|One Parent: Female|Unknown||||Yes||Self|General Community|Amachi|Match Support|F|Some Other Race||75|28213|Some College|Widowed|Human Services||20|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011184|502348258|31|0|2|41|0|2|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|
503689205|503689218|500739856|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|650|Red||2013-12-18|2014-01-08|2015-10-20|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||21.4||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|F|Black||46|28227|Masters Degree|Married|Finance|28202|8|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503691170|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502451190|502532871|500531332|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|877|Red||2011-04-14|2011-06-07|2013-10-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.8||1|1|1|1|M|Black||12|No|Mother|28273|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|M|White||29|28203|Bachelors Degree|Single|Tech: Computer/Programmer|28205|1|3|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502451637|31|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|10|||7462|13|||1|
502391396|503228398|500690843|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1401|Green|Cabarrus County|2013-04-01|2013-05-15|NaT||||46||2|2|1|1|F|Black||12|Yes|Mother|28052|One Parent: Female|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|White||40|28052|Bachelors Degree|Single|Transport: Pilot||1|1|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502391834|31|0|2|1|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
502391396|502202414|500540407|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|623|Red|Amachi, Project Big, Project Big AND Amachi|2011-06-08|2011-06-15|2013-02-27|Volunteer: Time constraint|Volunteer: Time constraint||20.5||2|2|1|1|F|Black||12|Yes|Mother|28052|One Parent: Female|Unknown||||No||Self|General Community|Cabarrus County|Match Support|F|Black||27|28273|Some College|Single|Finance||0|4|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500011746|502391834|31|0|2|31|0|2|10|2|500004772||4|3|500016374|-2|500000294|-2|0|10|||46|2|||1|500000294, 500004640, 500004901
503492220|503521240|500711792|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|726|Yellow||2013-09-18|2013-10-24|2015-10-20|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||23.9||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||27|28205|Bachelors Degree|Single|Business: Clerical|28277|0|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503494082|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
502526979|502616354|500541332|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|916|Green||2011-06-15|2011-06-17|2013-12-19|Child/Family: Moved|Child/Family: Moved||30.1||1|1|1|1|M|Hispanic||12|No|Mother|28209|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community|Project Big|Match Support|M|White||41|28202|Bachelors Degree|Divorced|Finance: Banking|28255|16|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502527432|3|0|1|1|0|1|10|2|-2||4|1|500004640|-2||-2|0|10|||7496|10|||1|
503530345|502460114|500704946|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|1182|Red|Cabarrus County|2013-07-26|2013-08-13|2016-11-07|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||38.8||1|1|2|2|F|Black||12|No|Mother|28025|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|RTBM|F|Black||43|28027|Masters Degree||Education: Teacher|28027|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|501204816|31|0|2|31|0|2|7|2|500016307||4|3|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
503703048|503354824|500753007|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1100|Green||2014-03-05|2014-03-12|NaT||||36.1||1|1|1|1|M|White||12|No|Mother|28226|One Parent: Female|$200,000 or more||||No||Self|General Community||Match Support|M|White||59|28104|Bachelors Degree|Married|Finance||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503705013|1|0|1|1|0|1|10|2|500009594||2|1||-2||-2|0|10|1562|2|7671|13|1561|2|1|
502875668|503114677|500649397|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1003|Red||2012-10-23|2012-10-31|2015-07-31|Volunteer: Time constraint|Volunteer: Time constraint||33||1|1|1|1|M|Black||12|No|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|M|Asian||39|28262|PHD|Married|Business: Mgt, Admin|28202|4|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502877071|31|0|1|4|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502527188|502591019|500544305|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|582|Green||2011-06-30|2011-08-15|2013-03-19|Volunteer: Time constraint|Volunteer: Time constraint||19.1||1|1|1|1|F|Hispanic||12|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes|Come Out and Play|Special Event|General Community||Enrollment|F|Hispanic||35|28207|Some College|Single|Human Services|28277|2|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502527641|3|0|2|3|0|2|5|2|-2||4|1||-2||-2|2203|12|||7462|13|||1|
502004276|502371255|500532829|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|660|Red||2011-04-21|2011-05-10|2013-02-28|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||21.7||1|1|1|1|M|Black||12|No|Mother|28215|One Parent: Female|Unknown||||Yes|AARTF|Neighbor/Friend|General Community||Match Support|M|White||46|28202|Bachelors Degree|Married|Unknown|28207|11|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502004675|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|6855|8|||7496|10|||1|
502697982|502832228|500609452|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|380|Red||2012-04-11|2012-05-16|2013-05-31|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||12.5||1|1|1|1|M|Black||12|No|Mother|28213|One Parent: Female|$60,000 to $74,999|||Y|No||Therapist/Counselor|General Community||Enrollment|M|Black||50|28269|Bachelors Degree|Married|Consultant|28262|8|0|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502698827|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|0|5|||9229|13|||1|
503885975|503885544|500769090|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|444|Red||2014-07-10|2014-08-01|2015-10-19|Volunteer: Moved|Volunteer: Moved||14.6||2|2|1|1|M|Black||12|No|Mother|28216|One Parent: Female|$45,000 to $49,999||||No||Relative|General Community||Match Support|M|White||28|28262|Associate Degree|Single|Finance: Banking|28081|1|1|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503887971|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|3|||17101|1|||1|
503021157|503089640|500658743|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|289|Yellow||2012-11-12|2013-01-23|2013-11-08|Volunteer: Time constraint|Volunteer: Time constraint||9.5||1|1|1|1|M|Black||12|No|Mother|28208|One Parent: Female|Unknown||||Yes||Relative|General Community||Enrollment|M|White||29|28203|Bachelors Degree|Single|Finance: Banking|28255|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500004169|503022696|31|0|1|1|0|1|5|2|-2||4|2||-2||-2|0|3|||7496|10|||1|
502969243|503083846|500628209|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|426|Yellow||2012-08-13|2012-09-04|2013-11-04|Volunteer: Time constraint|Volunteer: Time constraint||14||2|2|1|1|M|Some Other Race||12||Mother|28277|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|Asian||31|28273|Bachelors Degree|Single|Business: Engineer|29745|4|0||Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502970672|41|0|1|4|0|1|10|2|-2||4|2||-2||-2|0|10|||0|11|||1|
502969243|503837125|500759182|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|454|Yellow||2014-04-10|2014-04-25|2015-07-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||14.9||2|2|1|1|M|Some Other Race||12||Mother|28277|One Parent: Female|$20,000 to $24,999||||Yes||Self|General Community||Match Support|M|White||29|28209|Bachelors Degree|Single|Business|28281|0|1|Bowl For Kids Sake|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|502970672|41|0|1|1|0|1|10|2|-2||4|2||-2||-2|0|10|||132|8|||1|
503739899|503802084|500767689|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|987|Green||2014-06-25|2014-07-03|NaT||||32.4||1|1|1|1|F|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Insurance|28277|0|10|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503702247|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502605225|502538030|500540011|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|763|Red|Amachi, Project Big, Project Big AND Amachi|2011-06-06|2011-06-30|2013-08-01|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||25.1||1|1|1|1|F|Black||12|Yes|GrandFather|28216|Grandparents|Unknown||||Yes||School|General Community|Project Big, Project Big AND Amachi|Match Support|F|Black||32|28273|Bachelors Degree|Single|Finance||3|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502605742|31|0|2|31|0|2|10|2|500004772||4|3|500004640, 500004901|-2||-2|0|4|||7464|9|||1|500000294, 500004640, 500004901
503565188|503814392|500758306|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|401|Yellow||2014-04-04|2014-04-22|2015-05-28|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||13.2||2|2|1|1|M|Black||12|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||48|28269|Masters Degree|Married|Finance: Banking|28262|9|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503567063|31|0|1|31|0|1|10|2|-2||4|2||-2||-2|0|10|||46|2|||1|
502629201|502632871|500546227|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|12|Green||2011-07-14|2011-07-21|2011-08-02|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||0.4||2|2|2|2|M|White||12|No|Mother|28277|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|White||36|28226|Some College|Single|Business: Marketing||2|4|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500003657|502629856|1|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502629201|502893231|500603253|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1820|Green||2012-03-09|2012-03-22|NaT||||59.8||2|2|1|1|M|White||12|No|Mother|28277|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|White||32|28210|Bachelors Degree|Single|Business: Mgt, Admin|28226|1|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502629856|1|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503424337|503446943|500703604|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1042|Green||2013-07-15|2013-07-19|2016-05-26|Child/Family: Moved|Child/Family: Moved||34.2||1|1|1|1|F|Black||12||Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|Black||30|28173|Masters Degree|Single|Education|28262|0|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503426202|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|5|||7464|9|||1|
503930457|503544824|500773041|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|115|Green||2014-08-21|2014-08-30|2014-12-23|Child/Family: Moved|Child/Family: Moved||3.8||1|1|1|1|F|Black||12|No|Mother|28217|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||46|28226|Masters Degree|Married|Self-Employed, Entrepreneur|28277|16|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503932464|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||46|2|||1|
502869631|502962077|500618239|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|371|Red||2012-06-06|2012-06-21|2013-06-27|Volunteer: Time constraint|Volunteer: Time constraint||12.2||1|1|1|1|F|Black||12|No|Mother|28206|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Enrollment|F|White||45|28117|Bachelors Degree|Divorced|Business: Human Resources||8|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502871029|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
502290468|502873884|500596681|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1314|Red||2012-02-07|2012-02-10|2015-09-16|Child/Family: Moved|Child/Family: Moved||43.2||1|1|1|1|M|Black||12|No|Mother|28227|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Multi-race (Hispanic & White)||33|28204|PHD||Medical: Doctor, Provider||0|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502290900|31|0|1|35|0|1|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
502222548|502214317|500465659|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2396|Green||2010-08-13|2010-08-24|NaT||||78.7||1|1|1|1|M|Black||12|No|Mother|28216|One Parent: Female|Unknown||||No||School|General Community||Match Support|M|White||40|28211|Bachelors Degree|Married|Finance||2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020753|502222979|31|0|1|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|4|||7496|10|||1|
502367953|502658210|500548740|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1622|Yellow|Amachi|2011-08-04|2011-08-18|2016-01-26|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||53.3||1|1|1|1|M|Black||12|Yes|Mother|28208|One Parent: Female|Unknown|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|Black||43|28212|Masters Degree|Married|Retail: Mgt||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502368391|31|0|1|31|0|1|10|2|500003586||4|2|500000294|-2||-2|6854|8|||46|2|||1|500000294
503524260|503520196|500711429|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|372|Red||2013-09-17|2013-09-25|2014-10-02|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||12.2||1|1|1|1|M|Black||12|No|Mother|28217|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|Amachi|Enrollment|M|Black||30|28278|Associate Degree|Single|Tech: Research/Design|28217|10|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|503526133|31|0|1|31|0|1|5|2|-2||4|3|500000294|-2||-2|0|10|||7464|9|||1|
502068488|503953186|500771917|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|933|Green|Cabarrus County|2014-08-11|2014-08-26|NaT||||30.7||1|1|1|1|M|White||12|No|Mother|28269|One Parent: Female|$60,000 to $74,999||||No|Big|Neighbor/Friend|General Community|Cabarrus County|Match Support|M|White||35|28075|Masters Degree|Single|Finance: Accountant|28202|1|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502068912|1|0|1|1|0|1|10|2|500016307||2|1|500016374|-2|500016374|-2|6854|8|||7464|9|||1|500016374
503486227|503555261|500725969|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1232|Green||2013-10-31|2013-10-31|NaT||||40.5||1|1|1|1|M|Black||12|No|Mother|28270|One Parent: Female|$30,000 to $34,999||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|Black||32|28210|Bachelors Degree|Single|Tech: Research/Design|28273|0|9|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|503186577|31|0|1|31|0|1|10|2|-2||2|1||-2|500000294|-2|34|2|||46|2|||1|
503810996|503799211|500769226|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|959|Green||2014-07-11|2014-07-31|NaT||||31.5||1|1|1|1|M|Black||12|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||63|28078|Bachelors Degree|Married|Retired||0|0|Other|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017732|503812973|31|0|1|31|0|1|10|2|-2||2|1||-2|500007920, 500011315, 500011316|-2|0|10|||7671|13|||1|
502543116|502524371|500531887|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|246|Green|2010-2012 OJJDP JJI|2011-04-19|2011-05-04|2012-01-05|Child/Family: Moved|Child/Family: Moved||8.1||2|2|2|2|M|White||12|No|Mother|28027|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||62|28025||Married|Retired||0|0|Big Champions|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500002335|502543569|1|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|0|10|||7461|12|||1|500005291
502543116|502524371|500607345|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|40|Green||2012-03-30|2012-03-30|2012-05-09|Child: Severity of challenges|Child: Severity of challenges||1.3||2|2|2|2|M|White||12|No|Mother|28027|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|2010-2012 OJJDP JJI|Match Support|M|White||62|28025||Married|Retired||0|0|Big Champions|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500002335|502543569|1|0|1|1|0|1|10|2|-2||4|1|500005291|-2||-2|0|10|||7461|12|||1|
503866348|503862591|500767276|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|990|Green||2014-06-20|2014-06-30|NaT||||32.5||1|1|1|1|M|Black||12|No|GrandMother|28216|Grandparents|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|M|White||45|28269|Bachelors Degree|Married|Finance: Banking|28273|1|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503838583|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1|
502162237|502213773|500460265|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1208|Green|Amachi|2010-07-08|2010-07-12|2013-11-01|Volunteer: Moved|Volunteer: Moved||39.7||2|2|1|1|M|Black||12|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||29|28209|Bachelors Degree|Single|Business: Sales|28146|1|0|AA Task Force|Other Big|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500008321|503458866|31|0|1|1|0|1|10|2|-2||4|1|500000294|-2|500000294|-2|6854|8|||6247|12|||1|500000294
502162237|503151333|500756070|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1085|Red||2014-03-21|2014-03-27|NaT||||35.6||2|2|1|1|M|Black||12|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|Yes|Big|Neighbor/Friend|General Community|Amachi|Match Support|M|White||27|28202|Bachelors Degree|Single|Business|28217|0|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503458866|31|0|1|1|0|1|10|2|-2||2|3|500000294|-2||-2|6854|8|||7464|9|||1|
503941222|503889588|500772492|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|930|Yellow||2014-08-15|2014-08-29|NaT||||30.6||1|1|1|1|F|Black||12|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||28|28205|Masters Degree|Single|Business: Mgt, Admin|28262|2|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503931754|31|0|2|1|0|2|10|2|-2||2|2||-2||-2|0|4|||17159|12|||1|
503929747|503910740|500772491|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|700|Red||2014-08-15|2014-08-29|2016-07-29|Volunteer: Time constraint|Volunteer: Time constraint||23||1|1|1|1|F|Black||12|Yes|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Multi-race (Asian & White)||28|28203|Bachelors Degree|Single|Finance|28211|0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503931754|31|0|2|37|0|2|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
503638969|503503174|500736646|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1182|Green||2013-12-05|2013-12-20|NaT||||38.8||1|1|1|1|F|Black||12|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||23|28227||Single|Student: College|28202|2|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503640929|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
502431040|502609637|500550314|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1822|Green||2011-08-16|2011-08-31|2016-08-26|Child/Family: Moved|Child/Family: Moved||59.9||1|1|1|1|M|Black||12|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||35|28207|Masters Degree|Married|Law: Lawyer|28202|8|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020910|502431483|31|0|1|1|0|1|10|2|-2||4|1||-2|500004640|-2|0|10|||7496|10|||1|
503565637|503604089|500752839|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1097|Green||2014-03-05|2014-03-15|NaT||||36||1|1|1|1|M|Black||12|Yes|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||49|28204|Bachelors Degree|Married|Finance: Accountant|28255|8|0|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|503567522|31|0|1|1|0|1|10|2|-2||2|1|500000294|-2|500000294, 500014681|-2|34|2|||7464|9|||1|
503433257|503384599|500695071|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|485|Green||2013-04-30|2013-05-07|2014-09-04|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||15.9||1|1|1|1|F|Black||12|No|Father|28213|One Parent: Male|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Black||55|28269|Associate Degree|Single|Business||28|0|Self|Self|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500017777|503435122|31|0|2|31|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502527969|503169378|500662254|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|990|Red||2012-11-20|2012-12-01|2015-08-18|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||32.5||1|1|1|1|M|Black||11|No|Mother|28278|One Parent: Female|$35,000 to $39,999||||No||Self|General Community||Match Support|M|White||34|29708|High School Graduate|Single|Business: Mgt, Admin|29730|11|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502528422|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503259350|503370160|500687348|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1462|Green||2013-03-12|2013-03-15|NaT||||48||1|1|1|1|F|Black||11|No|Mother|28212|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Finance|28202|0|4|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503261158|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|34|2|||17161|11|||1|
503001802|502944301|500610527|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|279|Red||2012-04-18|2012-04-27|2013-01-31|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||9.2||1|1|2|2|F|Black||11|No|Mother|28206|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||58|28277|High School Graduate|Divorced|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503003296|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503425375|503546166|500704589|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|289|Red||2013-07-24|2013-07-30|2014-05-15|Child/Family: Moved|Child/Family: Moved||9.5||1|1|2|2|M|Black||11|No|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||49|28031|Associate Degree||Customer Service||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503427238|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503686272|503817633|500766948|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|658|Green||2014-06-18|2014-06-30|2016-04-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.6||1|1|1|1|M|Black||11|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Enrollment|M|White||32|28210|Masters Degree|Single|Finance|28211|8|1|Recruitment Event|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503688237|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7460|12|||1|
503691322|503763297|500752718|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1086|Green||2014-03-04|2014-03-26|NaT||||35.7||1|1|1|1|F|Black||11|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|F|Black||42|28273|Bachelors Degree|Single|Customer Service|28273|4|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503688237|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|5|||7464|9|||1|
503143377|503109316|500649731|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1581|Green||2012-10-23|2012-11-16|NaT||||51.9||1|1|1|1|F|Black||11|No|Mother|28210|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|F|White||28|28226|Bachelors Degree|Single|Education: Teacher|28173|2|6|TV|Media|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|503145049|31|0|2|1|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||130|1|||1|
502934728|503516330|500705674|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1310|Green||2013-08-02|2013-08-14|NaT||||43||1|1|1|1|M|Black||11|No|Mother|28215|One Parent: Female|$35,000 to $39,999||||Yes|Big|Neighbor/Friend|General Community||Match Support|M|Black||41|28211|Bachelors Degree|Single|Finance: Banking|28209|5|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|502936151|31|0|1|31|0|1|10|2|-2||2|1||-2|500000294|-2|6854|8|||7464|9|||1|
503609425|503572418|500730536|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|118|Green||2013-11-13|2013-12-20|2014-04-17|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.9||2|2|1|1|M|Black||11|No|GrandMother|28210|Grandparents|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||35|28210|Some College|Single|Finance: Accountant|28210|8|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500002334|503611302|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7464|9|||1|
503609425|503837417|500762429|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1028|Green||2014-05-07|2014-05-23|NaT||||33.8||2|2|1|1|M|Black||11|No|GrandMother|28210|Grandparents|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||34|28210|Masters Degree|Married|Finance: Banking|28202|8|8|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503611302|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
503723888|503858682|500779634|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|415|Red||2014-10-01|2014-10-13|2015-12-02|Volunteer: Time constraint|Volunteer: Time constraint||13.6||1|1|1|1|M|Black||11|Yes|Mother|28215|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Enrollment|M|Black||26|28227|Bachelors Degree|Single|Customer Service||1|3|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503725860|31|0|1|31|0|1|5|2|-2||4|3||-2||-2|0|10|||17101|1|||1|
502602926|503808719|500769460|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|954|Green||2014-07-14|2014-08-05|NaT||||31.3||1|1|1|1|F|Black||11|No|Mother|28216|One Parent: Female|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|Some Other Race||30|28214|Bachelors Degree|Married|Business|28214|1|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502603443|31|0|2|41|0|2|10|2|-2||2|1||-2||-2|6854|8|||7462|13|||1|
502299232|503510609|500703319|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|748|Yellow||2013-07-11|2013-07-30|2015-08-17|Child: Family structure changed|Child: Family structure changed||24.6||1|1|1|1|M|Black||11|Yes|GrandMother|28273|Foster Home|$25,000 to $29,999|||Y|Yes||Self|General Community|Amachi|Enrollment|M|White||32|28209|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|5|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500015820|501806520|31|0|1|1|0|1|5|2|-2||4|2|500000294|-2|500000294|-2|0|10|||7464|9|||1|
502653228|502192090|500552244|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2013|Green||2011-08-29|2011-09-11|NaT||||66.1||1|1|2|2|F|Black||11|No|Mother|28205|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|White||32|28134|Bachelors Degree|Single|Finance: Banking|28288|0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502653964|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502324604|502242614|500509702|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|946|Yellow||2011-01-07|2011-01-26|2013-08-29|Volunteer: Moved|Volunteer: Moved||31.1||3|3|1|1|F|Black||11|No|Mother|28216|One Parent: Female|Unknown||||Yes|TV|Media|General Community||Match Support|F|White||35|28210||Married|Law: Lawyer|28210|0|0||Relative|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500012459|502325039|31|0|2|1|0|2|10|2|-2||4|2||-2|500004640|-2|56|1|||0|11|||1|
502324604|503589790|500720750|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|372|Yellow||2013-10-18|2013-10-30|2014-11-06|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||12.2||3|3|1|1|F|Black||11|No|Mother|28216|One Parent: Female|Unknown||||Yes|TV|Media|General Community||Match Support|F|White||26|28262||Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|502325039|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|56|1|||7464|9|||1|
502211032|502276859|500508474|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1936|Yellow||2010-12-29|2011-01-14|2016-05-03|Volunteer: Time constraint|Volunteer: Time constraint||63.6||1|1|1|1|M|Black||11|No|Mother|28227|One Parent: Female|Unknown||||No|Big|Neighbor/Friend|General Community||Match Support|M|Some Other Race||38|28209|Bachelors Degree|Single|Business: Mgt, Admin|28205|5|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502211462|31|0|1|41|0|1|10|2|-2||4|2||-2||-2|6854|8|||7464|9|||1|
503492511|503852376|500764721|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|237|Red||2014-05-28|2014-06-13|2015-02-05|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||7.8||1|1|1|1|M|Black||11|No|Mother|28216|One Parent: Female|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||62|28210|Bachelors Degree|Divorced|Business: Engineer|28202|35|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503494379|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
502212246|502730900|500605715|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|243|Red||2012-03-22|2012-04-01|2012-11-30|Volunteer: Time constraint|Volunteer: Time constraint||8||2|2|1|1|F|Black||11|No|Mother|28134|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Enrollment|F|Black||46|28217|Some College|Single|Medical: Healthcare Worker|28210|9|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|501712386|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502212246|502238964|500461303|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|537|Green|Amachi|2010-07-16|2010-07-22|2012-01-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||17.6||2|2|1|1|F|Black||11|No|Mother|28134|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Enrollment|F|White||33|28210|Bachelors Degree|Single|Business: Human Resources|28202|4|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008629|501712386|31|0|2|1|0|2|5|2|500003586||4|1||-2||-2|0|10|||7464|9|||1|500000294
502274606|502441954|500518627|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2208|Green||2011-02-18|2011-02-28|NaT||||72.5||1|1|1|1|F|Black||11|No|Mother|28216|One Parent: Female|Unknown||||Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||29|28207|Bachelors Degree|Single|Human Services: Non-Profit|28212|1|4|Newspaper|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|502275038|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|6854|8|||129|1|||1|
503650948|504063702|500802395|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|149|Green|PERL 2014-2016|2014-12-09|2014-12-16|2015-05-14|Child/Family: Time constraints|Child/Family: Time constraints||4.9||2|2|2|2|M|Black||11|No|GrandMother|28270|Grandparents|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|M|White||57|28105|Bachelors Degree|Married|Business: Sales|28203|11|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018987|503652908|31|0|1|1|0|1|5|2|-2||4|1|500014681|-2|500000294|-2|0|10|||17159|12|||1|500014681
503650948|503605170|500742330|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|40|Green||2014-01-10|2014-02-26|2014-04-07|Volunteer: Time constraint|Volunteer: Time constraint||1.3||2|2|1|1|M|Black||11|No|GrandMother|28270|Grandparents|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|M|White||51|28110|Some College|Married|Arts, Entertainment, Sports||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503652908|31|0|1|1|0|1|5|2|-2||4|1|500014681|-2||-2|0|10|||46|2|||1|
502501346|502540731|500530910|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|429|Yellow|Amachi|2011-04-13|2011-04-26|2012-06-28|Volunteer: Moved|Volunteer: Moved||14.1||1|1|1|1|M|Hispanic||11|Yes|Mother|28213|One Parent: Female|$45,000 to $49,999||||Yes||Therapist/Counselor|General Community|Amachi|Enrollment|M|Hispanic||36|28269|Bachelors Degree|Single|Finance|28202|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|502501795|3|0|1|3|0|1|5|2|500003586||4|2|500000294|-2||-2|0|5|||7496|10|||1|500000294
503470937|500188541|500700189|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1371|Green||2013-06-11|2013-06-14|NaT||||45||1|1|3|3|F|Hispanic||11|No|Mother|28269|Two Parent|Unknown|||Y|Yes||Relative|General Community||Match Support|F|Hispanic||37|28203|Some College|Single|Education: Teacher|28217|5|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020753|502831178|3|0|2|3|0|2|10|2|-2||2|1||-2|500000294|-2|0|3|||2238|7|||1|
502972302|502842406|500603634|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|446|Green||2012-03-13|2012-03-17|2013-06-06|Child/Family: Moved|Child/Family: Moved||14.7||1|1|1|1|M|Black||11|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|Black||61|28027|Associate Degree|Married|Tech: Support, Writing||10|6|AA Task Force|BBBS Board/Staff|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500012459|502083880|31|0|1|31|0|1|10|2|-2||4|1||-2||-2|0|10|||9229|13|||1|
503281015|503585313|500731009|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|388|Green||2013-11-14|2013-11-25|2014-12-18|Child: Family structure changed|Child: Family structure changed||12.7||1|1|1|1|M|Black||11|No|Mother|28105|One Parent: Female|$30,000 to $34,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||45|28173|Bachelors Degree|Married|Finance|28277|13|5|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018987|503282834|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
504083467|504003996|500805363|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|815|Green|PERL 2014-2016|2014-12-19|2014-12-22|NaT||||26.8||1|1|1|1|M|Black||11|No|Mother|28226|One Parent: Female|$30,000 to $34,999||||No||School|General Community|PERL 2014-2016|Match Support|M|White||34|28214|Bachelors Degree||Transport: Flight Attendant|21804|7|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500018851|504085496|31|0|1|1|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681
503503497|503775803|500759857|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1051|Green||2014-04-16|2014-04-30|NaT||||34.5||1|1|1|1|M|Black||11|No|Mother|28216|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||29|28202|Bachelors Degree|Single|Finance|28202|1|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020910|503505371|31|0|1|1|0|1|10|2|-2||2|1|500000294|-2|500000294|-2|0|10|||7464|9|||1|
503580069|503556406|500713513|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|322|Red||2013-09-26|2013-09-30|2014-08-18|Child/Family: Moved|Child/Family: Moved||10.6||1|1|1|1|M|Multi-race (Black & Hispanic)||11|No|Mother|28270|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||27|28203|Bachelors Degree|Single|Finance: Banking|28210|2|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503581946|38|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
503489540|503488404|500707276|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|334|Yellow||2013-08-20|2013-08-31|2014-07-31|Volunteer: Moved|Volunteer: Moved||11||1|1|1|1|F|Black||11||Mother|28210|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Enrollment|F|White||27|28203|Masters Degree|Single|Finance: Accountant|28203|0|7|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|503491406|31|0|2|1|0|2|5|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
502464508|502901720|500609874|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|973|Red|Amachi|2012-04-13|2012-05-23|2015-01-21|Volunteer: Moved|Volunteer: Moved||32|Y|1|1|1|1|M|Black||11|Yes|Mother|28278|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community|Amachi|Match Support|F|White||34|29710|Bachelors Degree|Married|Education: Teacher||0|6|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502211737|31|0|1|1|0|2|10|2|500003586||4|3|500000294|-2||-2|0|10|||17161|11|||1|500000294
503569115|503619714|500735248|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|455|Green||2013-11-27|2013-12-19|2015-03-19|Child/Family: Moved|Child/Family: Moved||14.9||1|1|1|1|F|Black||11|No|Mother|2649|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||33|28203|Bachelors Degree|Single|Education: Teacher|28012|3|0|Self|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500015820|503570990|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502859181|502638002|500597079|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1828|Yellow||2012-02-08|2012-03-14|NaT||||60.1||1|1|1|1|F|Black||11|No|GrandMother|28205|Grandparents|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||40|28227|Masters Degree|Married|Tech: Support, Writing|28262|11|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|500187987|31|0|2|1|0|2|10|2|-2||2|2||-2||-2|0|10|||7462|13|||1|
503795417|503762193|500769015|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|386|Green||2014-07-09|2014-07-23|2015-08-13|Volunteer: Time constraint|Volunteer: Time constraint||12.7||1|1|1|1|F|Black||11|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Therapist/Counselor|General Community||RTBM|F|White||28|28211|Bachelors Degree|Single|Child/Day Care Worker||0|8|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503797394|31|0|2|1|0|2|7|2|-2||4|1||-2||-2|0|5|||17159|12|||1|
503741920|503696505|500754344|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|572|Green||2014-03-12|2014-03-26|2015-10-19|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||18.8||2|2|1|1|M|Black||11|No|Mother|28025|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||73|28226|PHD|Married|Retired||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503743892|31|0|1|1|0|1|10|2|-2||4|1|500016374|-2||-2|0|10|||7464|9|||1|
502675335|502643361|500555080|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|538|Yellow||2011-09-15|2011-09-22|2013-03-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.7||1|1|1|1|M|White||11|No|Mother|28105|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community||Match Support|M|White||51|28210|Bachelors Degree|Married|Self-Employed, Entrepreneur|28210|0|0|Self|Self|Big|General Site|mentor2.0, mentor2.0 2014|RTBM|0|1|1|0|277|60|598|500000170|500011746|502676163|1|0|1|1|0|1|10|2|-2||4|2||-2|500014505, 500014506|-1|0|10|||7464|9|||1|
502298007|501202092|500605225|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1795|Green||2012-03-20|2012-04-16|NaT||||59||2|2|2|2|F|Black||11|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|Black||41|28209|Bachelors Degree|Single|Finance: Banking|28255|0|6|TV|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502234907|31|0|2|31|0|2|10|2|-2||2|1|500004640|-2||-2|0|10|||130|1|||1|
502298007|502177426|500493839|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|320|Yellow|Project Big|2010-11-11|2010-12-09|2011-10-25|Volunteer: Moved|Volunteer: Moved||10.5||2|2|1|1|F|Black||11|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community|Project Big|Match Support|F|Black||27|28209|Some College|Single|Retail: Sales|28211|1|6|Self|Self|Big|General Community|Project Big|Enrollment|0|1|1|0|277|60|598|500000170|500011184|502234907|31|0|2|31|0|2|10|2|500004641||4|2|500004640|-2|500004640|-2|0|10|||7464|9|||1|500004640
502842247|503305101|500687640|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1451|Green||2013-03-13|2013-03-26|NaT||||47.7||1|1|1|1|M|White||11|No|Mother|28269|Other/Unknown|$15,000 to $19,999||||Yes||School|General Community||Match Support|M|White||47|28278|Bachelors Degree|Married|Finance: Banking|28210|0|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|502843540|1|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|
503904008|503820652|500768869|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|976|Green|VOL - Mentoring Hispanic Youth|2014-07-08|2014-07-14|NaT||||32.1||1|1|1|1|F|Hispanic||11|Yes|GrandMother|28216|One Parent: Female|Unknown||||Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||30|28203|Masters Degree|Single|Medical: Pharmacist|28213|0|6|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503906008|3|0|2|1|0|2|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1|500011312
502444611|501519220|500531694|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|178|Red||2011-04-18|2011-05-09|2011-11-03|Child/Family: Moved|Child/Family: Moved||5.8||1|1|2|2|F|Multi-race (Black & Hispanic)||11|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes|Michael Baisden|Media|General Community||Match Support|F|Black||54|28216|PHD|Married|Business: Mgt, Admin|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502445058|38|0|2|31|0|2|10|2|-2||4|3||-2||-2|6749|1|||7464|9|||1|
502619308|502709003|500565252|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|148|Red||2011-10-13|2011-10-31|2012-03-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.9||2|2|1|1|F|Hispanic||11|No|Mother|28212|Two Parent|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Hispanic||41|28215|Some College|Single|Business: Mgt, Admin|28202|6|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502619917|3|0|2|3|0|2|10|2|-2||4|3||-2||-2|0|10|||7462|13|||1|
502619308|503710698|500759246|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|791|Red||2014-04-10|2014-04-29|2016-06-28|Volunteer: Moved|Volunteer: Moved||26||2|2|1|1|F|Hispanic||11|No|Mother|28212|Two Parent|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||29|28206|Masters Degree|Single|Finance: Accountant|28210|3|0|United Way|Service Organization|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017777|502619917|3|0|2|1|0|2|10|2|-2||4|3||-2|500000294|-2|0|10|||16263|6|||1|
503545940|503804018|500760430|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1051|Green||2014-04-21|2014-04-30|NaT||||34.5||1|1|1|1|M|Black||11|No|Mother|28215|One Parent: Female|$45,000 to $49,999||||No||Self|General Community||Match Support|M|White||37|28205|Bachelors Degree|Married|Finance|28205|0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503547815|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1|
503367147|503500228|500704997|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|111|Red||2013-07-26|2013-08-21|2013-12-10|Volunteer: Moved|Volunteer: Moved||3.6||1|1|1|1|M|White||11||Mother|28270|One Parent: Female|$45,000 to $49,999||||No||Self|General Community||RTBM|M|Hispanic||42|28173||Married|Finance|28202|1|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503368992|1|0|1|3|0|1|7|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502664508|503029998|500639359|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|545|Red||2012-09-27|2012-09-28|2014-03-27|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17.9||1|1|1|1|M|Black||11||Aunt|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||36|28025|Some College|Married|Business|28288|7|0|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500013781|502665335|31|0|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
502982459|503565143|500713173|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|758|Green||2013-09-25|2013-09-30|2015-10-28|Volunteer: Time constraint|Volunteer: Time constraint||24.9||2|2|1|1|M|Black||11||Mother|28208|One Parent: Female|Less than $10,000|||Y|No||Self|General Community|PERL 2014-2016|Match Support|M|Black||30|28027|Bachelors Degree|Married|Business: Clerical|28282|3|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020990|502983913|31|0|1|31|0|1|10|2|-2||4|1|500014681|-2||-2|0|10|||7464|9|||1|
503634724|503529603|500753169|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|240|Green||2014-03-06|2014-03-18|2014-11-13|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.9||2|2|3|3|F|White||11|No|Father|28081|One Parent: Male|Unknown||||Yes||Self|General Community|Cabarrus County, PERL 2014-2016|Match Support|F|White||40|28078|Bachelors Degree|Single|Human Services: Social Worker|28277|0|9|Relative|Relative|Big|General Site|mentor2.0, mentor2.0 2015|Match Support|0|1|1|0|277|60|598|500000170|500013781|503636659|1|0|2|1|0|2|10|2|-2||4|1|500014681, 500016374|-2|500014505, 500015184|-1|0|10|||17161|11|||1|
503543014|503546166|500765902|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|994|Green||2014-06-09|2014-06-26|NaT||||32.7||1|1|2|2|M|Black||11|No|Mother|28269|One Parent: Female|$50,000 to $59,999||||No||Self|General Community||Match Support|M|White||49|28031|Associate Degree||Customer Service||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503544889|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502425281|502529075|500530096|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1964|Green||2011-04-08|2011-04-14|2016-08-29|Child/Family: Moved|Child/Family: Moved||64.5||1|1|1|1|F|Black||11|No|Mother|28273|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||61|28211|Bachelors Degree|Widowed|Real Estate: Realtor|28207|16|0|Other|BBBS Board/Staff|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500017777|502425720|31|0|2|1|0|2|10|2|-2||4|1||-2|500000294, 500004640|-2|0|10|||7671|13|||1|
502458411|502479222|500520070|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2200|Green||2011-02-24|2011-03-08|NaT||||72.3||1|1|1|1|F|Multi-race (Hispanic & White)||11|No|GrandMother|28210|Grandparents|$25,000 to $29,999|||Y|Yes|Big|Neighbor/Friend|General Community||Match Support|F|White||31|28211|Bachelors Degree|Single|Finance: Banking|28255|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi, Project Big|Match Support|0|1|0|1|277|60|598|500000170|500020753|502458858|35|0|2|1|0|2|10|2|-2||2|1||-2|500000294, 500004640|-2|6854|8|||7496|10|||1|
502948870|502984009|500616576|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1439|Green|Amachi|2012-05-25|2012-06-11|2016-05-20|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||47.3||1|1|1|1|F|Black||11|Yes|Mother|28216|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||Enrollment|F|White||28|28202|Bachelors Degree|Single|Finance: Banking||0|9|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503287812|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|10|||7496|10|||1|500000294
503381519|503803833|500758686|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1044|Green||2014-04-07|2014-05-07|NaT||||34.3||1|1|1|1|M|Black||11|No|Mother|28206|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||31|28204|Bachelors Degree|Single|Business|28262|1|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503383388|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503067218|503526377|500730492|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|994|Green||2013-11-13|2013-12-09|2016-08-29|Child: Lost interest|Child: Lost interest||32.7||1|1|1|1|M|Black||11|No|Mother|28227|One Parent: Female|$30,000 to $34,999|||Y|Yes||School|General Community||Match Support|M|White||38|28203||Single|Finance|28202|16|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503068877|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
503737886|503844296|500763770|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1015|Green||2014-05-19|2014-06-05|NaT||||33.3||1|1|1|1|M|Black||11|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||49|28205|Masters Degree|Domestic Partner|Business: Mgt, Admin|28277|3|9|Agency Sponsored|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503739858|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||16426|8|||1|
503764144|503784339|500773966|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|929|Green||2014-08-30|2014-08-30|NaT||||30.5||1|1|1|1|F|Black||11|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||37|28105|Masters Degree|Single|Education: Teacher||2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020910|503739858|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502840028|502782718|500589985|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|83|Red||2012-01-05|2012-02-07|2012-04-30|Volunteer: Time constraint|Volunteer: Time constraint||2.7||2|2|1|1|F|Black||11|No|Mother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|F|Black||32|28227||Married|Medical|28262|1|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502841320|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||46|2|||1|
502840028|502849360|500626309|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|92|Red||2012-07-26|2012-07-31|2012-10-31|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3||2|2|2|2|F|Black||11|No|Mother|28215|One Parent: Female|$30,000 to $34,999|||Y|Yes||Self|General Community||Match Support|F|White||28|28213|Bachelors Degree|Single|Medical: Nurse||0|4|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500008321|502841320|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503694415|503723380|500762190|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1016|Green|Cabarrus County|2014-05-05|2014-06-04|NaT||||33.4||1|1|1|1|M|Black||11|No|Mother|28083|One Parent: Female|$45,000 to $49,999|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|M|Black||50|28075|Masters Degree|Married|Law|28212|25|1|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|503696380|31|0|1|31|0|1|10|2|500016307||2|1|500016374|-2|500016374|-2|34|2|||7464|9|||1|500016374
503956230|504026743|500795032|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|846|Green||2014-11-12|2014-11-21|NaT||||27.8||1|1|1|1|M|Black||11|Yes|Mother|28227|One Parent: Female|$30,000 to $34,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Black||29|28210|Bachelors Degree|Single|Tech: Sales, Mktg|28262|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503958239|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1|
503446279|503842555|500759862|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1053|Green||2014-04-16|2014-04-28|NaT||||34.6||1|1|1|1|M|Black||11|No|Mother|28273|One Parent: Female|$40,000 to $44,999||||No||Self|General Community||Match Support|M|White||30|28101|Bachelors Degree|Single|Landscaper/Groundskeeper|28269|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503448145|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502861555|502866782|500595690|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|280|Red||2012-02-02|2012-02-10|2012-11-16|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||9.2||1|1|1|1|F|Black||11|No|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|White||30|28204|Bachelors Degree|Single|Business: Marketing|28226|0|5|BBBS National Site|Web Link|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500011349|502862935|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|4|||46|2|||1|
503585510|503580220|500731042|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|94|Green||2013-11-14|2013-11-22|2014-02-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||3.1||3|3|1|1|M|Black||11|No|Mother|28262|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Black||52|28269|Bachelors Degree|Married|Medical|28269|24|2|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017732|503587387|31|0|1|31|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||46|2|||1|
502656083|503108132|500678455|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1496|Green|Cabarrus County|2013-01-30|2013-02-09|NaT||||49.1||1|1|1|1|M|White||11|No|Mother|28083|One Parent: Female|Unknown||||Yes||Self|General Community|Cabarrus County|Match Support|M|White||59|28025|Some College|Married|Business: Sales|28025|8|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502656820|1|0|1|1|0|1|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
502920379|503497697|500708164|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1294|Green||2013-08-27|2013-08-30|NaT||||42.5||1|1|1|1|M|Black||11|Yes|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||28|28209|Bachelors Degree||Finance|28202|2|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|502921794|31|0|1|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
503867922|503834583|500766160|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|961|Green||2014-06-10|2014-07-29|NaT||||31.6||1|1|1|1|F|Black||11|No|Mother|28226|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||46|28207|Bachelors Degree|Married|Arts, Entertainment, Sports|28209|1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503126373|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
504004518|504055712|500800042|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|647|Green||2014-12-02|2014-12-22|2016-09-29|Volunteer: Time constraint|Volunteer: Time constraint||21.3||1|1|1|1|F|Some Other Race||11|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||Enrollment|F|White||24|28209|Bachelors Degree|Single|Business|28207|0|2|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500021785|504006533|41|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|4|||46|2|||1|
502782687|502760157|500595472|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1206|Red||2012-02-01|2012-03-06|2015-06-25|Volunteer: Moved|Volunteer: Moved||39.6||1|1|1|1|F|Black||11|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||26|28269|Some College||Medical|28216|0|3|Recruitment Event|BBBS Board/Staff|Big|General Community|Project Big|Match Support|0|1|0|1|277|60|598|500000170|500008321|502783868|31|0|2|31|0|2|10|2|-2||4|3||-2|500004640|-2|0|10|||7462|13|1207|5|1|
503296668|503922155|500777025|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|269|Yellow|PERL 2014-2016|2014-09-19|2014-09-29|2015-06-25|Child/Family: Moved|Child/Family: Moved||8.8||1|1|1|1|F|Black||11|No|Mother|28234|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|F|Multi-race (Black & White)||41|28270|Associate Degree|Divorced|Law: Security Officer|28262|1|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503298492|31|0|2|36|0|2|10|2|-2||4|2|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681
503388408|503761210|500769224|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|561|Red||2014-07-11|2014-07-29|2016-02-10|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||18.4||2|2|1|1|F|Black||11|No|Mother|28277|One Parent: Female|$30,000 to $34,999|||Y|No||School|General Community||Enrollment|F|Black||31|28270|Bachelors Degree|Single|Business: Sales||0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503390265|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
503388408|503432435|500696590|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|335|Red||2013-05-13|2013-06-21|2014-05-22|Volunteer: Time constraint|Volunteer: Time constraint||11||2|2|1|1|F|Black||11|No|Mother|28277|One Parent: Female|$30,000 to $34,999|||Y|No||School|General Community||Enrollment|F|Black||31|28270|High School Graduate|Single|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500013781|503390265|31|0|2|31|0|2|5|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
502882555|503438025|500695316|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|670|Green||2013-05-01|2013-05-16|2015-03-17|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||22||1|1|1|1|M|Black||11|No|Mother|28215|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|White||29|28208|Bachelors Degree|Single|Law: Police Officer|28216|3|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500011349|501090456|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
503411965|503792970|500754286|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1087|Green||2014-03-12|2014-03-25|NaT||||35.7||1|1|1|1|M|Black||11|No|Mother|28227|One Parent: Female|$45,000 to $49,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|White||26|28202|Bachelors Degree|Single|Consultant|28244|2|5|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503413822|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|34|2|||46|2|||1|
503383959|503572248|500713580|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1258|Green||2013-09-26|2013-10-05|NaT||||41.3||1|1|1|1|M|Black||11|Yes|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|M|White||27|28203|Bachelors Degree|Single|Real Estate: Realtor|28202|4|0|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|503554371|31|0|1|1|0|1|10|2|-2||2|1|500000294|-2|500000294|-2|0|10|||46|2|||1|
502869627|502932955|500608271|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1794|Green|Amachi|2012-04-05|2012-04-17|NaT||||58.9||1|1|1|1|F|Black||10|No|Mother|28206|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|F|White||28|28208|Bachelors Degree|Single|Business: Marketing|28269|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502871029|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|500000294
503297711|503353908|500681652|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1079|Yellow||2013-02-13|2013-02-26|2016-02-10|Child: Lost interest|Child: Lost interest||35.4||1|1|1|1|F|White||10|No|Mother|28226|One Parent: Female|$25,000 to $29,999||||No||School|General Community||Match Support|F|White||27|28207|Bachelors Degree|Single|Arts, Entertainment, Sports|28207|0|0|Billboard|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503299535|1|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|4|||125|1|||1|
504058316|503984749|500800274|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|820|Green||2014-12-02|2014-12-17|NaT||||26.9||1|1|1|1|M|Black||10|No|Mother|28208|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||29|28203|Masters Degree|Married|Business|28202|0|2|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|504060340|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|34|2|||7462|13|||1|
504030099|503994598|500793822|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|850|Green||2014-11-10|2014-11-17|NaT||||27.9||1|1|1|1|M|Black||10|No|Mother|28105|One Parent: Female|Unknown|||Y|Yes||School|General Community||Match Support|M|White||44|28211|Bachelors Degree|Married|Business: Human Resources|28255|9|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504032117|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|4|||7671|13|||1|
502776079|503573272|500711993|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1254|Green|Cabarrus County|2013-09-19|2013-10-09|NaT||||41.2||1|1|1|1|M|Black||10|Yes|Mother|28083|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Cabarrus County|Match Support|M|White||33|28269|Bachelors Degree|Single|Retail: Sales|28027|0|6|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|502777258|31|0|1|1|0|1|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
502643841|503991357|500783837|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|102|Green||2014-10-15|2014-10-20|2015-01-30|Volunteer: Time constraint|Volunteer: Time constraint||3.4||3|3|1|1|F|Black||10|Yes|Aunt|28227|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||53|28215||Married|Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500011349|502255582|31|0|2|31|0|2|10|2|-2||4|1|500000294|-2||-2|0|10|||7464|9|||1|
502643841|502638170|500548648|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1069|Yellow|Amachi|2011-08-04|2011-09-16|2014-08-20|Volunteer: Time constraint|Volunteer: Time constraint||35.1||3|3|1|1|F|Black||10|Yes|Aunt|28227|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||44|28269||Single|Business||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|502255582|31|0|2|31|0|2|10|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
502610111|501041084|500701839|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|943|Green||2013-06-25|2013-07-03|2016-02-01|Volunteer: Moved|Volunteer: Moved||31||1|1|1|1|F|Black||10|No|Mother|28211|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Enrollment|F|Black||46|28256|Associate Degree|Single|Finance: Banking||7|6|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|501288299|31|0|2|31|0|2|5|2|-2||4|1||-2||-2|0|10|||46|2|||1|
503076808|503688665|500758530|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|645|Green||2014-04-07|2014-05-20|2016-02-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||21.2||2|2|1|1|F|Multi-race (Black & White)||10|No|Mother|28115|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|White||46|28211|Bachelors Degree|Married|Finance|28105|11|4|BBBS National Site|Web Link|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500018851|503078467|36|0|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||46|2|||1|
503076808|503029978|500622847|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|469|Green|Amachi|2012-07-05|2012-07-23|2013-11-04|Volunteer: Moved|Volunteer: Moved||15.4||2|2|1|1|F|Multi-race (Black & White)||10|No|Mother|28115|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|White||30|28203|Bachelors Degree|Single|Finance: Accountant|28202|0|1|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|503078467|36|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|500000294
503389942|503191064|500695067|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1416|Green||2013-04-30|2013-04-30|NaT||||46.5||1|1|1|1|F|Black||10|No|Mother|28278|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||29|28205|Masters Degree|Single|Finance|28203|0|6|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020752|503239061|31|0|2|1|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
503047027|503087288|500639223|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|455|Red||2012-09-27|2012-11-29|2014-02-27|Volunteer: Time constraint|Volunteer: Time constraint||14.9||1|1|1|1|F|Hispanic||10|No|Mother|28211|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community||Match Support|F|Hispanic||36|28226|Bachelors Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|503045507|3|0|2|3|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502873192|502855289|500597685|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|480|Red||2012-02-10|2012-03-21|2013-07-14|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||15.8||1|1|1|1|F|Black||10|No|Mother|28206|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|F|White||25|28262|High School Graduate|Single|Customer Service|28269|0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502874592|31|0|2|1|0|2|5|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
503355399|503428702|500703056|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1336|Green||2013-07-09|2013-07-19|NaT||||43.9||1|1|1|1|F|Hispanic||10|No|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|M|White||35|28273|Masters Degree|Single|Finance: Accountant|28201|9|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020753|503348836|3|0|2|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
503585540|503485941|500709459|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|211|Yellow||2013-09-06|2013-09-24|2014-04-23|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||6.9||3|3|1|1|F|Black||10|No|GrandMother|28083|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|Black||45|28027|Masters Degree||Tech: Management|28262|13|0|Coworker|Workplace Partner|Big|General Community||RTBM|0|1|1|0|277|60|598|500000170|500012459|503587420|31|0|2|31|0|2|10|2|-2||4|2|500014681|-2||-2|34|2|||7447|3|||1|
503585540|503798839|500767384|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|372|Green||2014-06-23|2014-07-16|2015-07-23|Volunteer: Health|Volunteer: Health||12.2||3|3|1|1|F|Black||10|No|GrandMother|28083|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||37|28027|Some College|Married|Business: Mgt, Admin|28255|2|6|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|503587420|31|0|2|1|0|2|10|2|-2||4|1|500014681|-2||-2|34|2|||7439|1|||1|
503931637|504068281|500789322|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|867|Green||2014-10-29|2014-10-31|NaT||||28.5||1|1|1|1|M|Black||10|No|Mother|28208|One Parent: Female|$25,000 to $29,999|||Y|Yes||School|General Community||Match Support|M|White||40|28204|Bachelors Degree|Single|Business|28027|8|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503933644|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|4|||46|2|||1|
503246892|503350295|500691065|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1430|Green||2013-04-02|2013-04-16|NaT||||47||1|1|1|1|F|Black||10|Yes|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||29|28202|Bachelors Degree|Single|Business|28226|1|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503248691|31|0|2|1|0|2|10|2|-2||2|1|500000294|-2||-2|0|10|||7464|9|||1|
502688939|503023856|500619498|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1301|Yellow||2012-06-15|2012-06-21|2016-01-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||42.7||2|2|1|1|F|Black||10|No|Mother|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||37|28270|Bachelors Degree|Single|Finance: Banking||0|0|Recruitment Event|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500013781|501750989|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7458|9|||1|
502688939|502668908|500556512|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|156|Yellow||2011-09-21|2011-10-25|2012-03-29|Volunteer: Moved|Volunteer: Moved||5.1||2|2|1|1|F|Black||10|No|Mother|28215|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|Some Other Race||36|28078|Masters Degree|Separated|Finance: Accountant|28273|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501750989|31|0|2|41|0|2|10|2|-2||4|2||-2||-2|0|10|||7496|10|||1|
502543702|503346987|500702244|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1226|Green||2013-06-27|2013-07-10|2016-11-17|Volunteer: Time constraint|Volunteer: Time constraint||40.3|Y|2|2|1|1|M|Black||10|No|Mother|28269|One Parent: Female|$40,000 to $44,999||||No||School|General Community||Match Support|M|White||34|28078|Bachelors Degree|Married|Business: Mgt, Admin|28262|2|10|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017732|502544155|31|0|1|1|0|1|10|2|-2||4|1||-2|500000294|-2|0|4|||7464|9|||1|
502544010|502641777|500549950|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|2022|Green||2011-08-12|2011-08-31|2017-03-14|Volunteer: Time constraint|Volunteer: Time constraint||66.4||1|1|1|1|F|Black||10|No|Mother|28269|One Parent: Female|$40,000 to $44,999||||No||School|General Community||Enrollment|F|White||29|28202|Bachelors Degree|Single|Service: Hotel||0|3|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|502544463|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502950100|502466985|500691514|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|175|Red|Amachi|2013-04-04|2013-04-24|2013-10-16|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.7||1|1|1|1|M|Black||10|Yes|GrandMother|28215|Grandparents|Unknown||||Yes||Self|General Community||RTBM|M|Black||25|28208|High School Graduate|Single|Business: Mgt, Admin|28227|1|2|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500011746|502951526|31|0|1|31|0|1|7|2|-2||4|3||-2||-2|0|10|||7464|9|||1|500000294
502661304|502640462|500548919|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1071|Yellow|Amachi|2011-08-07|2011-08-25|2014-07-31|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||35.2||1|1|1|1|F|Black||10|Yes|GrandMother|28208|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|Amachi|Enrollment|F|Black||28|28215|Bachelors Degree|Single|Tech: Management|28217|0|4|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|502662054|31|0|2|31|0|2|5|2|500003586||4|2|500000294|-2||-2|0|10|||7464|9|||1|500000294
503569406|503534366|500706542|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1295|Green||2013-08-13|2013-08-29|NaT||||42.5||1|1|1|1|F|Multi-race (Black & Hispanic)||10|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||28|28207|PHD|Married|Medical: Healthcare Worker|28025|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503567063|38|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502931159|503802032|500759587|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1051|Green||2014-04-14|2014-04-30|NaT||||34.5||1|1|1|1|M|Black||10|No|Mother|28214|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||45|28214|Masters Degree|Married|Business|28207|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502932575|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503402178|503468005|500700142|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1338|Green||2013-06-10|2013-07-17|NaT||||44||1|1|1|1|M|Black||10|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|M|White||31|28203|Bachelors Degree|Single|Finance|28202|5|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503404035|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|3|||7496|10|||1|
503586001|503568168|500711704|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|720|Red||2013-09-18|2013-09-26|2015-09-16|Child: Lost interest|Child: Lost interest||23.7||1|1|1|1|F|Black||10|No|Mother|28212|One Parent: Female|$35,000 to $39,999|||Y|Yes||Self|General Community||Match Support|F|Black||38|28262|Masters Degree|Divorced|Finance|28202|3|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503587878|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
503586069|503541572|500711744|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|720|Red||2013-09-18|2013-09-26|2015-09-16|Child: Lost interest|Child: Lost interest||23.7||1|1|1|1|F|Black||10|No|Mother|28212|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|F|Black||47|28269|Bachelors Degree|Married|Medical: Nurse|28078|8|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503587878|31|0|2|31|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502934732|503537424|500722866|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1234|Green||2013-10-24|2013-10-29|NaT||||40.5||1|1|1|1|M|Black||10|No|Mother|28215|One Parent: Female|$35,000 to $39,999||||Yes||Self|General Community||Match Support|M|White||29|28211|Bachelors Degree|Single|Business: Marketing|28262|3|0|Recruitment Event|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|502936151|31|0|1|1|0|1|10|2|-2||2|1||-2|500000294|-2|0|10|||7458|9|||1|
502843866|502951469|500609886|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|881|Red||2012-04-13|2012-04-26|2014-09-24|Child/Family: Moved|Child/Family: Moved||28.9||1|1|1|1|F|Black||10|No|Mother|28212|One Parent: Female|$20,000 to $24,999|Yes: Active|No||Yes||Relative|General Community||Match Support|F|White||31|28203|Bachelors Degree|Single|Business|27401|0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|502845159|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|0|3|||7496|10|||1|
503471046|503489178|500703315|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1115|Green||2013-07-11|2013-07-30|2016-08-18|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||36.6||1|1|1|1|M|White||10|No|Mother|28210|One Parent: Female|$60,000 to $74,999||||No||Self|General Community||Match Support|M|Asian||29|28134|Masters Degree|Single|Finance: Accountant|28202|1|8|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500021785|503472912|1|0|1|4|0|1|10|2|-2||4|1||-2|500000294|-2|0|10|||7496|10|||1|
502778215|503291713|500682140|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1484|Green||2013-02-14|2013-02-21|NaT||||48.8||1|1|1|1|M|Black||10|No|Mother|28217|One Parent: Female|Less than $10,000|||Y|Yes||Relative|General Community||Match Support|M|White||28|28209|Masters Degree|Single|Finance: Accountant||0|6|Relative|Relative|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502610737|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|3|||17161|11|||1|
503259551|503371077|500700569|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|603|Red||2013-06-13|2013-06-26|2015-02-19|Volunteer: Time constraint|Volunteer: Time constraint||19.8||2|2|1|1|F|Black||10||Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||55|28209|Some College|Divorced|Business: Clerical|28273|20|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503261359|31|0|2|1|0|2|10|2|-2||4|3||-2||-2|34|2|||7464|9|||1|
503834826|503675532|500767892|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|168|Red||2014-06-26|2014-07-16|2014-12-31|Volunteer: Time constraint|Volunteer: Time constraint||5.5||2|2|2|2|F|Black||10|No|Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Enrollment|F|White||39|28134|Masters Degree|Separated|Business: Human Resources|28202|1|0|Self|Self|Big|General Site||Enrollment|0|1|1|0|277|60|598|500000170|500008321|503836805|31|0|2|1|0|2|5|2|-2||4|3||-2||-1|0|10|||7464|9|||1|
503873009|503953864|500789610|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|374|Red||2014-10-29|2014-11-21|2015-11-30|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||12.3||1|1|1|1|M|White||10|No|Mother|28270|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Enrollment|M|White||28|28270|Bachelors Degree|Living w/ Significant Other|Law: Police Officer|28211|0|9|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503875005|1|0|1|1|0|1|5|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
502946633|502893902|500605537|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1787|Green||2012-03-21|2012-04-24|NaT||||58.7||1|1|1|1|F|Black||10|No|GrandMother|28208|Grandparents|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||31|28209|Masters Degree|Single|Medical: Healthcare Worker|28079|0|4|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|502948059|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|4|||7464|9|||1|
503582752|503771996|500766377|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|997|Green||2014-06-12|2014-06-23|NaT||||32.8||1|1|1|1|F|Black||10|No|Mother|28212|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|Black||35|28104|Some College|Single|Medical: Healthcare Worker|28105|2|7|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500020910|502908938|31|0|2|31|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
503634722|503597445|500743535|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1150|Green|Cabarrus County|2014-01-17|2014-01-21|NaT||||37.8||1|1|1|1|F|White||10|No|Father|28081|One Parent: Male|Unknown|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|White||50|28226|Bachelors Degree||Human Services: Non-Profit|28208|0|6|Self|Self|Big|General Community|Cabarrus County|Enrollment|0|1|0|1|277|60|598|500000170|500013781|503636659|1|0|2|1|0|2|10|2|-2||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
503671417|504022116|500799802|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|822|Green||2014-12-01|2014-12-15|NaT||||27||1|1|1|1|M|Black||10|No|Mother|28206|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|M|White||28|28203|Masters Degree|Single|Business|28277|0|1|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503673378|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|34|2|||17159|12|||1|
503230851|503317475|500693795|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|661|Yellow||2013-04-19|2013-04-22|2015-02-12|Child/Family: Moved|Child/Family: Moved||21.7||1|1|1|1|F|Black||10|No|Mother|28216|One Parent: Female|$10,000 to $14,999|||Y|Yes|Big|Neighbor/Friend|General Community||Enrollment|F|White||28|28205|Bachelors Degree|Single|Business|28255|0|3|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500015820|503232639|31|0|2|1|0|2|5|2|-2||4|2||-2|500000294|-2|6854|8|||7464|9|||1|
503144476|503453981|500700084|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|1197|Red||2013-06-10|2013-06-18|2016-09-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||39.3||1|1|1|1|M|Black||10|Yes|GrandMother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes|AARTF|BBBS Board/Staff|General Community|Amachi|Enrollment|M|White||29|28269|Masters Degree|Living w/ Significant Other|Business: Mgt, Admin|28203|0|7|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|503146148|31|0|1|1|0|1|5|2|-2||4|3|500000294|-2|500000294|-2|7294|13|||7464|9|||1|
503836529|503876514|500775633|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|911|Green||2014-09-12|2014-09-17|NaT||||29.9||1|1|1|1|M|Multi-race (Black & Hispanic)||10|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||27|28211|Bachelors Degree|Single|Finance|29715|1|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503838508|38|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1|
503662361|503740772|500758213|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|573|Green||2014-04-03|2014-04-25|2015-11-19|Volunteer: Time constraint|Volunteer: Time constraint||18.8||1|1|1|1|M|Black||10|Yes|Mother|28216|One Parent: Female|$45,000 to $49,999|||Y|Yes||Self|General Community||Match Support|M|White||33|28031|Bachelors Degree|Single|Tech: Engineer|28081|6|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503664337|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503835875|503926804|500772936|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|917|Green||2014-08-20|2014-09-11|NaT||||30.1||1|1|1|1|M|Black||10|No|Mother|28217|One Parent: Female|$25,000 to $29,999|||Y|Yes||Relative|General Community||Match Support|M|White||47|28278|Bachelors Degree|Married|Business: Mgt, Admin|29732|4|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503837854|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|3|||17159|12|||1|
503804106|503988181|500777910|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|380|Green||2014-09-24|2014-09-29|2015-10-14|Volunteer: Moved|Volunteer: Moved||12.5||2|2|1|1|M|Black||10|No|Mother|28202|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||RTBM|M|White||25|28209|Bachelors Degree|Single|Tech: Computer/Programmer|28202|0|1|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503712061|31|0|1|1|0|1|7|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
504051221|503972520|500786442|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|288|Yellow||2014-10-22|2014-11-10|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||9.5||1|1|1|1|F|Black||10|No|Mother|28203|One Parent: Female|Less than $10,000|||Y|Yes||School|General Community||RTBM|F|White||34|28203|Masters Degree|Single|Business||0|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|504053245|31|0|2|1|0|2|7|2|-2||4|2||-2||-2|0|4|||17159|12|||1|
503224812|503385277|500692915|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1430|Green||2013-04-15|2013-04-16|NaT||||47||1|1|1|1|F|Black||10|No|Mother|28215|One Parent: Female|$15,000 to $19,999||||Yes||Self|General Community||Match Support|F|White||33|28210|Bachelors Degree|Single|Tech: Support, Writing|28217|0|6|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503226552|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1|
503589761|503582412|500718535|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|718|Yellow||2013-10-11|2013-10-28|2015-10-16|Volunteer: Health|Volunteer: Health||23.6||2|2|1|1|F|Black||10|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||27|28203|Bachelors Degree|Single|Child/Day Care Worker|28214|10|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|503591638|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503001538|503380945|500686972|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|876|Green||2013-03-11|2013-03-27|2015-08-20|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||28.8||1|1|1|1|M|Black||10|No|Mother|28205|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||34|28203|Masters Degree|Single|Real Estate: Realtor||5|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018987|503003032|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
503321228|503412979|500691563|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1401|Green||2013-04-04|2013-05-15|NaT||||46||1|1|1|1|M|Multi-race (Black & White)||10||Mother|28226|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Multi-race (Asian & White)||35|28209|Bachelors Degree|Single|Business: Mgt, Admin||1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503323062|36|0|1|37|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503650774|503526078|500746685|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1108|Green||2014-02-03|2014-03-04|NaT||||36.4||1|1|1|1|M|Black||10|No|Mother|28226|One Parent: Female|$20,000 to $24,999||||No|BBBS National Site|Web Link|General Community||Match Support|M|Some Other Race||38|28277|Masters Degree|Married|Finance: Banking|28228|7|0|Big For A Day|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503652734|31|0|1|41|0|1|10|2|-2||2|1||-2||-2|34|2|||16422|8|||1|
503995241|503924249|500783860|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|572|Green|PERL 2014-2016|2014-10-15|2014-10-22|2016-05-16|Volunteer: Time constraint|Volunteer: Time constraint||18.8||1|1|1|1|F|Black||10|No|Mother|28213|One Parent: Female|$30,000 to $34,999|||Y|Yes|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|F|White||32|28270|Associate Degree|Married|Arts, Entertainment, Sports|28203|3|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500018851|503997256|31|0|2|1|0|2|10|2|-2||4|1|500014681|-2|500014681|-2|34|2|||17159|12|||1|500014681
503468785|503856524|500765157|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1015|Green||2014-06-02|2014-06-05|NaT||||33.3||1|1|1|1|M|Black||10|No|Mother|28262|One Parent: Female|$50,000 to $59,999|Yes: Active|No||No||Self|General Community||Match Support|M|Black||46|28078||Married|Unemployed||0|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503470651|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||7671|13|||1|
503565647|503577080|500758415|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|329|Yellow||2014-04-04|2014-04-10|2015-03-05|Volunteer: Time constraint|Volunteer: Time constraint||10.8||2|2|1|1|M|Black||10|Yes|Mother|28216|One Parent: Female|Less than $10,000||||Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|White||43|28269|Bachelors Degree|Married|Business: Marketing|28262|2|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|503567522|31|0|1|1|0|1|10|2|-2||4|2|500000294|-2||-2|34|2|||7464|9|1360|3|1|
503461190|503672434|500753717|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|519|Yellow||2014-03-10|2014-03-24|2015-08-25|Volunteer: Time constraint|Volunteer: Time constraint||17.1||1|1|1|1|M|Multi-race (Black & White)||10|No|Mother|28081|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|White||51|28027|Some College|Married|Business: Marketing|28027|1|5|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|503463056|36|0|1|1|0|1|10|2|||4|2||-2||-2|0|10|||7464|9|||1|
503681425|503786945|500773494|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|747|Red|PERL 2014-2016|2014-08-26|2014-09-18|2016-10-04|Child: Family structure changed|Child: Family structure changed||24.5||1|1|2|2|M|Multi-race (Black & White)||10|Yes|Mother|28025|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County, PERL 2014-2016, VOL - Incarcerated Parents|Match Support|M|Asian||27|28075|Bachelors Degree|Single|Finance: Banking|28202|3|0|Local Print|Media|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|503683390|36|0|1|4|0|1|10|2|-2||4|3|500007918, 500014681, 500016374|-2|500014681, 500016374|-2|34|2|||7439|1|||1|500014681
503602769|503919845|500787263|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|413|Green||2014-10-23|2014-11-10|2015-12-28|Volunteer: Moved|Volunteer: Moved||13.6||2|2|1|1|F|Black||10|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|F|Black||25|28213|Bachelors Degree|Single|Finance: Banking|28216|0|10|Billboard|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020990|503604646|31|0|2|31|0|2|10|2|-2||4|1|500007920, 500011315, 500011316, 500014681|-2||-2|0|10|||125|1|||1|
503226693|503035671|500682567|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1486|Green||2013-02-18|2013-02-19|NaT||||48.8||1|1|1|1|F|Black||10|No|Father|28213|One Parent: Male|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|Black||56|28269|Bachelors Degree|Single|Business: Mgt, Admin|28262|25|0|Other|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503228481|31|0|2|31|0|2|10|2|500014421||2|1||-2||-2|0|4|||7671|13|||1|
503883171|502138981|500769877|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|936|Green||2014-07-17|2014-08-23|NaT||||30.8||1|1|3|3|F|Black||9|No|Mother|28213|One Parent: Female|$30,000 to $34,999||||Yes||Self|General Community||Match Support|F|Black||29|28262|Bachelors Degree|Single|Student: College||1|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503885167|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||7496|10|||1|
503587467|503886373|500768974|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|966|Green||2014-07-09|2014-07-24|NaT||||31.7||1|1|1|1|M|Black||9|Yes|Mother|28262|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|M|White||31|28117|Bachelors Degree|Single|Finance: Accountant|28677|0|5|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503587387|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1|
503778456|503787440|500763996|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|797|Green||2014-05-21|2014-05-31|2016-08-05|Volunteer: Moved|Volunteer: Moved||26.2||1|1|1|1|M|Black||9|No|Mother|28208|One Parent: Female|$10,000 to $14,999|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|M|White||31|28277|Bachelors Degree|Single|Finance: Economist|28277|1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503780433|31|0|1|1|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
503589735|503488419|500720851|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|601|Green||2013-10-18|2013-10-25|2015-06-18|Volunteer: Moved|Volunteer: Moved||19.7||1|1|1|1|F|Black||9|No|Mother|28208|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|F|White||26|28209|Bachelors Degree|Single|Retail: Sales|28209|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503591612|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
503062537|503455629|500695323|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1400|Green||2013-05-01|2013-05-16|NaT||||46||2|2|1|1|F|Black||9|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|White||54|28211|Bachelors Degree|Separated|Retired||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501090456|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7462|13|||1|
503062537|502911343|500623747|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|217|Yellow||2012-07-11|2012-08-14|2013-03-19|Volunteer: Time constraint|Volunteer: Time constraint||7.1||2|2|1|1|F|Black||9|No|Mother|28215|One Parent: Female|Unknown||||Yes||Self|General Community||Match Support|F|Black||28|28215|Bachelors Degree|Single|Business||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011349|501090456|31|0|2|31|0|2|10|2|-2||4|2||-2||-2|0|10|||7464|9|||1|
503774068|503866555|500767047|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|996|Green||2014-06-18|2014-06-24|NaT||||32.7||1|1|1|1|M|Multi-race (Black & Hispanic)||9|No|Mother|28215|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|M|Hispanic||37|28202|Bachelors Degree|Single|Consultant|27607|1|0|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503776034|38|0|1|3|0|1|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1|
503866363|503946948|500771529|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|945|Green||2014-08-06|2014-08-14|NaT||||31||1|1|1|1|F|Black||9|No|GrandMother|28216|Grandparents|$25,000 to $29,999|||Y|Yes||Self|General Community||Match Support|F|White||48|28269|Some College|Married|Finance: Banking|28262|0|0|Current/Previous Big|Relative|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500008321|503838583|31|0|2|1|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||17160|11|||1|
503862843|503926694|500788150|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|800|Green|PERL 2014-2016|2014-10-27|2014-11-04|2017-01-12|Volunteer: Time constraint|Volunteer: Time constraint||26.3||1|1|1|1|F|Black||9|No|Aunt|28208|Other Relative|Less than $10,000|||Y|Yes||Self|General Community|PERL 2014-2016|Enrollment|F|White||54|28078|Associate Degree|Single|Medical|28025|10|7|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020910|502431630|31|0|2|1|0|2|5|2|-2||4|1|500014681|-2|500000294, 500014681|-2|0|10|||7464|9|||1|500014681
503476611|503495634|500704993|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|678|Red||2013-07-26|2013-08-15|2015-06-24|Volunteer: Moved|Volunteer: Moved||22.3||1|1|1|1|M|Multi-race (Black & Asian)||9||Mother|28226|One Parent: Female|$20,000 to $24,999|||Y|Yes||School|General Community||Match Support|M|White||29|28208|Bachelors Degree|Single|Unknown|28202|0|2|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503478477|39|0|1|1|0|1|10|2|-2||4|3||-2||-2|0|4|||7464|9|||1|
504106075|503995246|500799241|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|822|Green|PERL 2014-2016|2014-11-25|2014-11-28|2017-02-27|Volunteer: Time constraint|Volunteer: Time constraint||27||1|1|1|1|F|Black||9|No|Mother|28208|One Parent: Female|$25,000 to $29,999||||No||School|General Community|PERL 2014-2016|Enrollment|F|Black||22|28208|Bachelors Degree|Single|Medical: Nurse|28278|0|7|Self|Self|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500018851|503933644|31|0|2|31|0|2|5|2|-2||4|1|500014681|-2|500014681|-2|0|4|||7464|9|||1|500014681
503454717|503349725|500691603|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|419|Red||2013-04-05|2013-04-26|2014-06-19|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||13.8||2|2|1|1|F|Black||9|No|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||50|28214|Associate Degree|Single|Medical|28210|2|5|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500013781|504995618|31|0|2|31|0|2|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|10|||7464|9|||1|
503225825|502916764|500679932|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|586|Green||2013-02-05|2013-02-21|2014-09-30|Volunteer: Time constraint|Volunteer: Time constraint||19.3||3|3|1|1|F|White||9|No|Mother|28027|Two Parent|Unknown||||Yes||School|General Community|Cabarrus County|Match Support|F|White||47|28075|Masters Degree|Divorced|Business: Marketing|28282|5|6|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500015820|503227613|1|0|2|1|0|2|10|2|-2||4|1|500016374|-2||-2|0|4|||7464|9|||1|
503225825|503551624|500794940|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|720|Red||2014-11-12|2014-11-19|2016-11-08|Volunteer: Time constraint|Volunteer: Time constraint||23.7||3|3|1|1|F|White||9|No|Mother|28027|Two Parent|Unknown||||Yes||School|General Community|Cabarrus County|Match Support|F|White||29|28138|Bachelors Degree|Single|Customer Service|28269|2|5|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500020753|503227613|1|0|2|1|0|2|10|2|-2||4|3|500016374|-2|500016374|-2|0|4|||7464|9|||1|
503585543|500189320|500709465|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1150|Red|Cabarrus County|2013-09-06|2013-09-25|2016-11-18|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||37.8||1|1|3|3|F|Black||9|No|GrandMother|28083|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community|Cabarrus County|Match Support|F|Black||46|28025|Some College|Single|Finance: Banking|28204|0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|503587420|31|0|2|31|0|2|10|2|500016307||4|3|500016374|-2|500016374|-2|34|2|||7464|9|||1|500016374
503953662|503952799|500772194|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|795|Green|Amachi|2014-08-13|2014-08-29|2016-11-01|Volunteer: Time constraint|Volunteer: Time constraint||26.1||1|1|1|1|F|Black||9|Yes|Mother|28208|One Parent: Female|Less than $10,000||||Yes||Therapist/Counselor|General Community||Enrollment|F|White||26|28209|Masters Degree|Single|Education: Teacher|28212|2|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|503955662|31|0|2|1|0|2|5|2|-2||4|1||-2||-2|0|5|||7496|10|||1|500000294
503798419|502994003|500761356|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|519|Yellow|Amachi|2014-04-28|2014-04-30|2015-10-01|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||17.1||1|1|1|1|F|Black||9|Yes|Mother|28269|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community|Amachi|Match Support|F|Black||26|28212|Some College||Medical: Nurse||2|0|Recruitment Event|BBBS Board/Staff|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500012459|503800396|31|0|2|31|0|2|10|2|-2||4|2|500000294|-2|500000294|-2|34|2|||7462|13|||1|500000294
503286862|503386901|500701858|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1359|Green||2013-06-25|2013-06-26|NaT||||44.6||1|1|1|1|F|Black||9||Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||29|28269|Bachelors Degree|Single|Medical: Nurse||1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503261359|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503663973|503865770|500763734|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|287|Red||2014-05-19|2014-05-22|2015-03-05|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||9.4||2|2|2|2|M|Black||9|Yes|Mother|28204|One Parent: Female|$25,000 to $29,999||||Yes||Self|General Community||Match Support|M|White||42|28205|Bachelors Degree|Married|Arts, Entertainment, Sports|28205|14|0|Current/Previous Big|Other Big|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017777|503665933|31|0|1|1|0|1|10|2|-2||4|3||-2|500000294|-2|0|10|||17159|12|||1|
503739912|503929189|500772941|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|932|Green||2014-08-20|2014-08-27|NaT||||30.6||1|1|1|1|M|Black||9|No|Mother|28208|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|Black||35|28217|Some College|Married|Law: Police Officer|28229|0|8|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503702247|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|0|10|||17101|1|||1|
503663417|504057497|500800835|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|818|Green||2014-12-03|2014-12-19|NaT||||26.9||1|1|1|1|M|Black||9|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|M|White||34|28269|Bachelors Degree|Living w/ Significant Other|Tech: Sales, Mktg|28117|2|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503665377|31|0|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503530548|503635342|500756727|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1086|Green||2014-03-26|2014-03-26|NaT||||35.7||1|1|1|1|F|Black||9|Yes|GrandMother|28208|One Parent: Female|$15,000 to $19,999|||Y|Yes||Self|General Community|Amachi|Match Support|F|Black||31|28269||Single|Unemployed||0|0|Recruitment Event|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503146148|31|0|2|31|0|2|10|2|500003586||2|1|500000294|-2||-2|0|10|||7458|9|||1|
503833932|503698988|500761753|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|687|Green||2014-04-30|2014-05-12|2016-03-29|Child/Family: Time constraints|Child/Family: Time constraints||22.6||1|1|2|2|F|Black||9|No|Mother|28208|Two Parent|$15,000 to $19,999|||Y|Yes|BBBS National Site|Web Link|General Community||Enrollment|F|White||48|28031|Bachelors Degree|Separated|Business: Marketing|28601|16|0|BBBS National Site|Web Link|Big|General Community|Amachi, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500018851|503835911|31|0|2|1|0|2|5|2|-2||4|1||-2|500000294, 500007920, 500011315, 500011316|-2|34|2|||46|2|||1|
503834833|503968276|500783899|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|869|Green|PERL 2014-2016|2014-10-15|2014-10-29|NaT||||28.6||1|1|1|1|M|Black||9|No|Mother|28206|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community|PERL 2014-2016|Match Support|M|Hispanic||30|28227|Bachelors Degree|Single|Retail: Sales|28105|8|0|Current/Previous Big|Relative|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500008321|503836805|31|0|1|3|0|1|10|2|-2||2|1|500014681|-2|500014681|-2|0|10|||17160|11|||1|500014681
503955220|503874105|500772805|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|925|Green||2014-08-19|2014-09-03|NaT||||30.4||1|1|1|1|F|Multi-race (Black & Hispanic)||9|No|Mother|28212|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||28|28203|Bachelors Degree|Single|Education: Teacher|28078|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|503838508|38|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
503366783|503493458|500709610|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1273|Green||2013-09-09|2013-09-20|NaT||||41.8||1|1|1|1|M|Black||9|No|Mother|28216|One Parent: Female|$45,000 to $49,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|Black||35|28216|Some College|Married|Tech: Engineer|28120|0|7|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503368628|31|0|1|31|0|1|10|2|-2||2|1||-2||-2|34|2|||7464|9|||1|
503496397|503797696|500772113|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|932|Green||2014-08-12|2014-08-27|NaT||||30.6||1|1|1|1|F|Hispanic||9|No|Mother|28212|One Parent: Female|Unknown|||Y|Yes||Relative|General Community||Match Support|F|Hispanic||25|28210|Bachelors Degree|Single|Business: Sales|28277|2|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503498265|3|0|2|3|0|2|10|2|-2||2|1||-2||-2|0|3|||7464|9|||1|
503558194|503527934|500705245|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1312|Green||2013-07-30|2013-08-12|NaT||||43.1||1|1|1|1|F|Black||9|Yes|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|Black||47|28269|Associate Degree|Single|Tech: Computer/Programmer|28269|21|0|Big For A Day|Special Event|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|503560069|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||16422|8|||1|
503575837|503825634|500766748|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|993|Green|VOL - Mentoring Hispanic Youth|2014-06-16|2014-06-27|NaT||||32.6||1|1|1|1|F|Hispanic||9|No|Mother|28206|One Parent: Female|Unknown||||Yes|Spanish Radio|Media|General Community||Match Support|F|Hispanic||37|28206|Masters Degree|Single|Unknown|28223|1|0|Local Radio|Media|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|503577713|3|0|2|3|0|2|10|2|-2||2|1||-2|500014681|-2|7068|1|||7437|1|||1|500011312
503579909|503552956|500707000|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1296|Green||2013-08-16|2013-08-28|NaT||||42.6||1|1|1|1|F|Black||8|No|Mother|28203|One Parent: Female|$10,000 to $14,999|||Y|Yes||Self|General Community||Match Support|F|White||40|28204|Masters Degree|Single|Finance: Banking|28212|5|7|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500018851|502958068|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
503798824|503895001|500783536|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|881|Green||2014-10-14|2014-10-17|NaT||||28.9||1|1|1|1|F|Black||8|Yes|Mother|28211|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community|Amachi|Match Support|F|White||26|28277|Bachelors Degree|Single|Business|28273|1|9|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503800801|31|0|2|1|0|2|10|2|-2||2|1|500000294|-2||-2|0|10|||7439|1|||1|
503554921|503556149|500742082|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|553|Green||2014-01-09|2014-01-30|2015-08-06|Child/Family: Moved|Child/Family: Moved||18.2||1|1|1|1|F|Black||8|No|Mother|28203|One Parent: Female|Less than $10,000|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||33|28277|Bachelors Degree|Single|Insurance|28277|3|0|Self|Self|Big|General Community||Enrollment|0|1|0|1|277|60|598|500000170|500015820|503556796|31|0|2|1|0|2|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
503654738|503853843|500772115|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|931|Green||2014-08-12|2014-08-28|NaT||||30.6||2|2|1|1|F|Black||8|No|Mother|28216|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|Asian||31|28202|Bachelors Degree|Single|Business: Sales|28217|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|500740560|31|0|2|4|0|2|10|2|-2||2|1||-2||-2|34|2|||7496|10|||1|
503654738|503646353|500737114|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|162|Yellow||2013-12-06|2013-12-31|2014-06-11|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.3||2|2|1|1|F|Black||8|No|Mother|28216|One Parent: Female|$25,000 to $29,999|||Y|Yes|BBBS National Site|Web Link|General Community||Match Support|F|White||24|28031||Single|Student: College||0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500012459|500740560|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|34|2|||46|2|||1|
503717075|503842851|500762275|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|419|Yellow||2014-05-06|2014-05-16|2015-07-09|Volunteer: Moved|Volunteer: Moved||13.8||2|2|1|1|F|Black||8|Yes|Mother|28216|One Parent: Female|Less than $10,000|||Y|Yes||Self|General Community||Match Support|F|White||33|28202|Masters Degree|Single|Consultant|28202|0|1|Man Up Campaign|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500015820|503719040|31|0|2|1|0|2|10|2|-2||4|2||-2||-2|0|10|||17101|1|||1|
503572810|503785317|500764166|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|516|Green||2014-05-22|2014-05-31|2015-10-29|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||17||1|1|1|1|M|Multi-race (Black & White)||8|No|Mother|28115|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|White||45|28031|Bachelors Degree|Married|Real Estate: Realtor|28031|20|0|Local Print|Media|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500012459|503078467|36|0|1|1|0|1|5|2|-2||4|1||-2||-2|0|10|||7439|1|||1|
503993975|503947272|500797389|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|829|Green||2014-11-19|2014-12-08|NaT||||27.2||1|1|1|1|F|Black||8|Yes|Mother|28262|One Parent: Female|$25,000 to $29,999||||No||Self|General Community||Match Support|F|White||40|28205|Bachelors Degree|Divorced|Law|28204|2|6|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503969639|31|0|2|1|0|2|10|2|-2||2|1||-2||-2|0|10|||17159|12|||1|
504069856|502591360|500786507|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|841|Green|Cabarrus County|2014-10-22|2014-11-26|NaT||||27.6||1|1|2|2|F|Black||8|No|Mother|28083|One Parent: Female|$25,000 to $29,999|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||69|28027||Married|Business: Mgt, Admin||0|0|Self|Self|Big|General Community|Cabarrus County|Match Support|0|1|0|1|277|60|598|500000170|500022817|504071884|31|0|2|31|0|2|10|2|500016307||2|1|500016374|-2|500016374|-2|0|10|||7464|9|||1|500016374
504096330|503992956|500794009|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|731|Red|Cabarrus County|2014-11-10|2014-11-21|2016-11-21|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||24||1|1|1|1|F|Black||8|Yes|GrandMother|28083|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Amachi, Cabarrus County|Match Support|F|White||25|28081||Single|Medical: Admin||0|0|BBBS National Site|Web Link|Big|General Community|Cabarrus County|Enrollment|0|1|0|1|277|60|598|500000170|500022817|503587420|31|0|2|1|0|2|10|2|500016307||4|3|500000294, 500016374|-2|500016374|-2|0|10|||46|2|||1|500016374
504096289|503776419|500790461|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|731|Red|Cabarrus County|2014-10-30|2014-11-21|2016-11-21|Child/Family: Infraction of match rules/agency policies|Child/Family: Infraction of match rules/agency policies||24||1|1|1|1|F|Black||8|Yes|GrandMother|28083|One Parent: Female|Unknown|||Y|Yes||Self|General Community|Cabarrus County|Match Support|F|Black||28|28027|Masters Degree|Single|Human Services: Social Worker|28202|1|1|Self|Self|Big|General Community|Cabarrus County, PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500022817|503587420|31|0|2|31|0|2|10|2|500016307||4|3|500016374|-2|500014681, 500016374|-2|0|10|||7464|9|||1|500016374
504044312|503862152|500783874|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|875|Green||2014-10-15|2014-10-23|NaT||||28.7||1|1|1|1|F|Black||8|No|Mother|28213|One Parent: Female|$20,000 to $24,999|||Y|Yes||Self|General Community||Match Support|F|Black||27|28269|Some College|Single|Business|28269|4|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|504046330|31|0|2|31|0|2|10|2|-2||2|1||-2||-2|0|10|||46|2|||1|
503774486|503792812|500766439|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|875|Green||2014-06-12|2014-06-27|2016-11-18|Volunteer: Moved|Volunteer: Moved||28.7||1|1|1|1|F|Black||8|No|Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|Yes|BBBS National Site|Web Link|General Community||RTBM|F|Black||63|28213||Single|Retired||0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017732|503776463|31|0|2|31|0|2|7|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
502242649|502576783|500536543|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|348|Red|2010-2012 OJJDP JJI|2011-05-17|2011-05-27|2012-05-09|Volunteer: Moved|Volunteer: Moved||11.4||1|1|1|1|M|Hispanic|Dominican|17|No|Mother|28212|One Parent: Female|Unknown|||Y|No|Big|Neighbor/Friend|General Community|2010-2012 OJJDP JJI|Enrollment|M|Hispanic||44|28211|Masters Degree|Married|Finance: Banking|28277|2|10|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502243080|3|13|1|3|0|1|5|2|-2||4|3|500005291|-2||-2|6854|8|||7462|13|||1|500005291
501023404|501510589|500359415|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|375|Green||2009-04-24|2009-05-01|2010-05-11|Volunteer: Moved|Volunteer: Moved||12.3||2|2|1|1|F|Hispanic|Mexican|22|No|Mother|28273|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|F|White||33|28202|Juris Doctorate (JD)|Single|Law: Lawyer|28202|0|3|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500009242|501023677|3|10|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502627461|502615885|500550750|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|398|Red|2010-2012 OJJDP JJI|2011-08-18|2011-08-26|2012-09-27|Volunteer: Time constraint|Volunteer: Time constraint||13.1||1|1|1|1|F|Hispanic|Mexican|20|Yes|Mother|28269|One Parent: Female|Unknown|||Y|Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|F|White||52|28205|Some College|Single|Self-Employed, Entrepreneur||16|0|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500011746|502628116|3|10|2|1|0|2|10|2|-2||4|3|500005291|-2|500005291|-2|0|4|||7464|9|||1|500005291
502527168|501646021|500618440|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1532|Red||2012-06-07|2012-06-19|2016-08-29|Child: Graduated|Child: Graduated||50.3||1|1|2|2|M|Hispanic|Mexican|19|No|Mother|28215|One Parent: Female|Less than $10,000|||Y|Yes|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|M|Hispanic||30|28227|||Business: Engineer|28202|0|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502527621|3|10|1|3|0|1|10|2|-2||4|3|500005291|-2||-2|2203|12|||7464|9|||1|
502528773|502552143|500539575|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|349|Red|2010-2012 OJJDP JJI|2011-06-03|2011-06-16|2012-05-30|Volunteer: Moved|Volunteer: Moved||11.5||1|1|1|1|F|Hispanic|Mexican|18|No|Mother|28215|One Parent: Female|Unknown||||No|Come Out and Play|Special Event|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||36|28262|Masters Degree|Single|Finance|28273|3|10|BBBS National Site|Web Link|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500011746|502529226|3|10|2|3|0|2|10|2|-2||4|3|500005291|-2|500005291|-2|2203|12|||46|2|||1|500005291
502627468|503419352|500696276|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|367|Green||2013-05-09|2013-05-17|2014-05-19|Child: Lost interest|Child: Lost interest||12.1||1|1|1|1|M|Hispanic|Mexican|18|No|Mother|28269|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|White||30|28036|Some College|Single|Business|28078|0|1|Neighbor/Friend|Neighbor/Friend|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500017777|502628116|3|10|1|1|0|1|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1|
502627466|502800101|500591158|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|848|Green||2012-01-11|2012-01-18|2014-05-15|Volunteer: Moved|Volunteer: Moved||27.9||1|1|1|1|M|Hispanic|Mexican|18|No|Mother|28269|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Multi-race (Hispanic & White)||28|28202|Bachelors Degree|Single|Finance||0|3|Local TV|Media|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502628116|3|10|1|35|0|1|10|2|-2||4|1||-2||-2|0|4|||7438|1|||1|
502853025|503009880|500621608|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|321|Green||2012-06-25|2012-07-11|2013-05-28|Child: Lost interest|Child: Lost interest||10.5||1|1|1|1|F|Hispanic|Mexican|17|No|Mother|28205|Two Parent|Unknown|||Y|Yes||School|General Community||Match Support|F|Hispanic||40|28277|Some College|Married|Self-Employed, Entrepreneur||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502854420|3|10|2|3|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
500841232|500834757|500166629|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|918|Green||2007-03-13|2007-03-20|2009-09-23|Volunteer: Time constraint|Volunteer: Time constraint||30.2||1|1|1|1|M|Hispanic|Mexican|16|No|Mother|28269|One Parent: Female|Unknown||||No||Self|General Community||Enrollment|M|Hispanic|Mexican|48|28269|Bachelors Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500009242|500829324|3|10|1|3|10|1|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
502374716|502014837|500491463|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|686|Green|Project Big|2010-11-05|2010-11-11|2012-09-27|Volunteer: Moved|Volunteer: Moved||22.5||2|2|1|1|M|Hispanic|Mexican|16|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Hispanic||38|28204||Single|Finance: Banking||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community|Project Big|Match Support|0|1|1|0|277|60|598|500000170|500011746|502375154|3|10|1|3|0|1|10|2|500004641||4|1||-2|500004640|-2|0|4|||7496|10|||1|500004640
502374716|503560077|500723012|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1234|Green||2013-10-24|2013-10-29|NaT||||40.5||2|2|1|1|M|Hispanic|Mexican|16|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|M|Hispanic||29|28214|Bachelors Degree|Single|Self-Employed, Entrepreneur|28214|0|0|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|502375154|3|10|1|3|0|1|10|2|-2||2|1||-2||-2|0|4|||46|2|||1|
502627470|502672424|500552887|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|980|Green||2011-09-01|2011-09-12|2014-05-19|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||32.2||1|1|1|1|M|Hispanic|Mexican|16|No|Mother|28269|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|Asian||26|28105|Some College|Single|Student: College||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502628116|3|10|1|4|0|1|5|2|-2||4|1||-2||-2|0|4|||7496|10|||1|
503490571|503645850|500738556|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|510|Red|VOL - Mentoring Hispanic Youth|2013-12-12|2013-12-20|2015-05-14|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||16.8||1|1|1|1|F|Hispanic|Mexican|16|No|Mother|28208|Two Parent|Unknown|||Y|Yes|Spanish Radio|Media|General Community||Match Support|F|White||35|28214|Bachelors Degree|Single|Transport: Flight Attendant|85034|0|3|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500017777|503492439|3|10|2|1|0|2|10|2|-2||4|3||-2|500000294|-2|7068|1|||7464|9|||1|500011312
502859440|503046471|500623399|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|628|Green||2012-07-10|2012-08-01|2014-04-21|Volunteer: Time constraint|Volunteer: Time constraint||20.6||1|1|1|1|F|Hispanic|Mexican|15|No|Mother|28215|Two Parent|Unknown||||Yes||School|General Community||Match Support|F|Multi-race (Hispanic & White)||30|28202|Bachelors Degree|Married|Finance: Banking|28255|4|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502860839|3|10|2|35|0|2|10|2|-2||4|1||-2||-2|0|4|||7496|10|||1|
502874566|502894480|500607372|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1240|Green||2012-03-30|2012-05-24|2015-10-16|Volunteer: Moved|Volunteer: Moved||40.7||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28205|One Parent: Female|$10,000 to $14,999|||Y|Yes||School|General Community||Match Support|F|White||28|27235|Bachelors Degree||Business: Engineer||1|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502875969|3|10|2|1|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502339704|502539104|500552221|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|393|Red|2010-2012 OJJDP JJI|2011-08-29|2011-08-31|2012-09-27|Child/Family: Moved|Child/Family: Moved||12.9||2|2|1|1|F|Hispanic|Mexican|14|No|Mother|28212|One Parent: Female|Unknown||||No||Relative|General Community|2010-2012 OJJDP JJI|Match Support|F|Black||39|28211|Masters Degree|Single|Business|28211|0|6|Self|Self|Big|General Community|2010-2012 OJJDP JJI|Match Support|0|1|1|0|277|60|598|500000170|500011746|502340140|3|10|2|31|0|2|10|2|-2||4|3|500005291|-2|500005291|-2|0|3|||7464|9|||1|500005291
502339704|502275098|500499962|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|218|Green||2010-11-29|2010-12-06|2011-07-12|Volunteer: Moved|Volunteer: Moved||7.2||2|2|1|1|F|Hispanic|Mexican|14|No|Mother|28212|One Parent: Female|Unknown||||No||Relative|General Community|2010-2012 OJJDP JJI|Match Support|F|Hispanic||34|28262||Single|Education: Teacher||0|0|Neighbor/Friend|Neighbor/Friend|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500010765|502340140|3|10|2|3|0|2|10|2|-2||4|1|500005291|-2||-2|0|3|||7496|10|||1|
503895506|504026849|500784082|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|877|Green|VOL - Mentoring Hispanic Youth, PERL 2014-2016|2014-10-15|2014-10-21|NaT||||28.8||1|1|1|1|F|Hispanic|Mexican|14|No|Mother|28212|Two Parent|Unknown|||Y|Yes||School|General Community|PERL 2014-2016|Match Support|F|Hispanic||30|28226||Single|Unemployed||0|0|Relative|Relative|Big|General Community|PERL 2014-2016|Match Support|0|1|0|1|277|60|598|500000170|500020753|503897502|3|10|2|3|0|2|10|2|-2||2|1|500014681|-2|500014681|-2|0|4|||17161|11|||1|500011312, 500014681
503706992|503709061|500761338|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1051|Green|VOL - Mentoring Hispanic Youth|2014-04-28|2014-04-30|NaT||||34.5||1|1|1|1|F|Hispanic|Mexican|13|No|Mother|28205|One Parent: Female|Unknown|||Y|Yes|BBBS National Site|Web Link|General Community|VOL - Mentoring Hispanic Youth|Match Support|F|White||44|28213|Bachelors Degree|Married|Medical|28216|2|6|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020753|503708958|3|10|2|1|0|2|10|2|-2||2|1|500011312|-2||-2|34|2|||7464|9|||1|500011312
503398288|503473834|500707156|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|479|Yellow||2013-08-19|2013-08-31|2014-12-23|Volunteer: Moved|Volunteer: Moved||15.7||1|1|1|1|M|Hispanic|Mexican|12|No|Mother|28206|One Parent: Female|$15,000 to $19,999|||Y|Yes||Therapist/Counselor|General Community||Match Support|M|White||28|28202|Masters Degree|Single|Consultant||0|11|Neighbor/Friend|Neighbor/Friend|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017777|503400145|3|10|1|1|0|1|10|2|-2||4|2||-2|500000294|-2|0|5|||7496|10|||1|
500970181|500969057|500203109|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1764|Red||2007-10-11|2007-10-31|2012-08-29|Child: Severity of challenges|Child: Severity of challenges||58||1|1|1|1|M|Black|Other African|20|No|Mother|28208|One Parent: Female|$15,000 to $19,999|||Y|No|BBBS National Site|Web Link|General Community||Match Support|M|White||37|28210|Bachelors Degree|Single|Finance: Accountant||1|0|BBBS National Site|Web Link|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500001281|500970452|31|31|1|1|0|1|10|2|-2||4|3||-2||-2|34|2|||46|2|||1|
501872144|502063676|500460156|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2421|Green||2010-07-07|2010-07-30|NaT||||79.5||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown|||Y|Yes||Relative|General Community||Match Support|M|White||35|28205|Masters Degree|Married|Tech: Engineer|28115|1|1|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500020752|501872517|31|31|1|1|0|1|10|2|-2||2|1||-2||-2|0|3|||46|2|||1|
501860404|501893096|500425993|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|922|Green||2010-01-11|2010-01-21|2012-07-31|Volunteer: Moved|Volunteer: Moved||30.3||1|1|1|1|M|Black|Other African|17|No|Mother|28269|One Parent: Female|Unknown||||No|BBBS National Site|Web Link|General Community||Enrollment|M|White||30|28202||Single|Finance||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|501860777|31|31|1|1|0|1|5|2|-2||4|1||-2||-2|34|2|||7464|9|||1|
502632678|503007956|500616542|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|98|Yellow||2012-05-25|2012-06-08|2012-09-14|Child: Family structure changed|Child: Family structure changed||3.2||1|1|1|1|M|Black|Other African|17|No|Mother|28212|One Parent: Female|$20,000 to $24,999|||Y|Yes||Relative|General Community||Match Support|M|Black||54|28269|Masters Degree|Single|Tech: Computer/Programmer|28212|5|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500001281|502633334|31|31|1|31|0|1|10|2|-2||4|2||-2||-2|0|3|||7462|13|||1|
502455004|502680045|500553363|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|2004|Green|2010-2012 OJJDP JJI|2011-09-06|2011-09-20|NaT||||65.8||1|1|1|1|M|Black|Other African|15|No|Mother|29732|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI|Match Support|M|White||31|29720|Bachelors Degree|Married|Business: Sales|28134|4|0|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500013781|502074089|31|31|1|1|0|1|10|2|-2||2|1|500005291|-2||-2|0|4|||7464|9|||1|500005291
502859604|502863229|500604130|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|997|Green||2012-03-14|2012-03-26|2014-12-18|Volunteer: Time constraint|Volunteer: Time constraint||32.8||1|1|1|1|F|Hispanic|Other Central American|19|No|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community||Match Support|F|Hispanic||40|28214|Some College|Single|Student: College||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502860998|3|14|2|3|0|2|10|2|-2||4|1||-2||-2|0|4|||7464|9|||1|
502421671|502272620|500524198|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|43|Red|Project Big, 2010-2012 OJJDP JJI|2011-03-09|2011-03-31|2011-05-13|Child/Family: Lost contact with volunteer/agency|Child/Family: Lost contact with volunteer/agency||1.4||1|1|1|1|F|Hispanic|Other Central American|16|No|Mother|28213|One Parent: Female|Unknown||||Yes||School|General Community|2010-2012 OJJDP JJI, Project Big|Match Support|F|White||31|28202|Some College|Single|Business: Marketing||3|0|Self|Self|Big|General Community|Project Big|Enrollment|0|1|1|0|277|60|598|500000170|500010765|502422110|3|14|2|1|0|2|10|2|500004641||4|3|500004640, 500005291|-2|500004640|-2|0|4|||7464|9|||1|500004640, 500005291
502838495|502707985|500605723|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|42|Green||2012-03-22|2012-04-24|2012-06-05|Volunteer: Unrealistic expectations|Volunteer: Unrealistic expectations||1.4||1|1|1|1|F|Hispanic|Other Central American|16|No|Mother|28213|Grandparents|Unknown|||Y|Yes||School|General Community||Match Support|F|Hispanic||38|28202||Single|Unknown||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502839787|3|14|2|3|0|2|10|2|-2||4|1||-2||-2|0|4|||7462|13|||1|
502859599|502864237|500610310|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|735|Green||2012-04-17|2012-04-30|2014-05-05|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||24.1||1|1|1|1|M|Hispanic|Other Central American|14|No|Mother|28205|One Parent: Female|Unknown||||Yes||School|General Community||Enrollment|M|Hispanic|Other South American|35|28209|High School Graduate|Married|Business||0|1|Relative|Relative|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502860998|3|14|1|3|15|1|5|2|-2||4|1||-2||-2|0|4|||17161|11|||1|
504059280|503998203|500796014|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|622|Red|VOL - Mentoring Hispanic Youth|2014-11-15|2014-12-16|2016-08-29|Child: Family structure changed|Child: Family structure changed||20.4||1|1|1|1|M|Hispanic|Other Central American|13|No|Mother|28214|One Parent: Female|Unknown|||Y|Yes||Therapist/Counselor|General Community|VOL - Mentoring Hispanic Youth|Match Support|M|Hispanic||37|28078|Associate Degree|Single|Finance|28217|0|3|Coworker|Workplace Partner|Big|General Community|VOL - Mentoring Hispanic Youth|Match Support|0|1|0|1|277|60|598|500000170|500017777|504061304|3|14|1|3|0|1|10|2|-2||4|3|500011312|-2|500011312|-2|0|5|||7447|3|||1|500011312
502859609|502863010|500601876|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|790|Green||2012-03-02|2012-03-20|2014-05-19|Volunteer: Moved|Volunteer: Moved||26||1|1|1|1|F|Hispanic|Other Central American|11|No|Mother|28205|Two Parent: Not Married|Unknown||||Yes||School|General Community||Match Support|F|Black||34|28205|Bachelors Degree|Single|Business: Mgt, Admin|95354|2|6|AA Task Force|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|502860998|3|14|2|31|0|2|10|2|-2||4|1||-2||-2|0|4|||9229|13|||1|
503355390|503468187|500703060|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|390|Red||2013-07-09|2013-07-17|2014-08-11|Volunteer: Time constraint|Volunteer: Time constraint||12.8||2|2|1|1|F|Hispanic|Other Central American|10|No|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|RTBM|F|White||42|29708|Bachelors Degree|Single|Tech: Sales, Mktg||0|0|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017777|503348836|3|14|2|1|0|2|7|2|-2||4|3|500011312, 500014681|-2|500000294|-2|0|10|||7464|9|||1|
503355390|503843020|500777040|BBBS of Greater Charlotte|Main Office|N|C|Completed|RTBM|375|Yellow|VOL - Mentoring Hispanic Youth|2014-09-19|2014-09-29|2015-10-09|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||12.3||2|2|2|2|F|Hispanic|Other Central American|10|No|Mother|28217|One Parent: Female|Unknown||||Yes||Self|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|RTBM|F|Hispanic||23|28226|Some College|Single|Student: College|28207|3|0|Self|Self|Big|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|0|1|277|60|598|500000170|500017777|503348836|3|14|2|3|0|2|7|2|-2||4|2|500011312, 500014681|-2|500007920, 500011312, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|500011312
503467766|503543048|500717156|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|1241|Green||2013-10-08|2013-10-22|NaT||||40.8||1|1|1|1|F|Hispanic|Other Central American|9|No|Mother|28262|One Parent: Female|Unknown|||Y|Yes||Self|General Community||Match Support|F|White||30|28214|Bachelors Degree|Single|Law: Paralegal|28214|2|5|Self|Self|Big|General Community|Amachi|Match Support|0|1|0|1|277|60|598|500000170|500013781|502751081|3|14|2|1|0|2|10|2|-2||2|1||-2|500000294|-2|0|10|||7464|9|||1|
500896588|500924445|500183434|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|3253|Green||2007-07-10|2007-07-20|2016-06-15|Child: Graduated|Child: Graduated||106.9||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28273|Two Parent|Less than $10,000|||Y|No||Self|General Community||Match Support|F|White||36|28269|Masters Degree|Married|Education|28205|6|6|Other|BBBS Board/Staff|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020752|500896858|3|15|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7671|13|||1|
502738004|502620216|500579434|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|114|Red||2011-11-17|2011-11-30|2012-03-23|Volunteer: Infraction of match rules/agency policies|Volunteer: Infraction of match rules/agency policies||3.7||1|1|1|1|F|Hispanic|Other South American|18|No|Mother|28262|Two Parent: Not Married|Unknown|||Y|No||Self|General Community||Match Support|F|Hispanic||36|28202||Single|Finance: Banking||1|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502738904|3|15|2|3|0|2|10|2|-2||4|3||-2||-2|0|10|||7464|9|||1|
501023408|501356600|500296545|BBBS of Greater Charlotte|Main Office|N|C|Active|Match Support|3053|Green||2008-10-08|2008-11-05|NaT||||100.3||1|1|1|1|M|Hispanic|Other South American|17|No|Mother|28273|One Parent: Female|Less than $10,000||||Yes||Self|General Community||Match Support|M|White||32|28203|Bachelors Degree|Single|Business: Sales||0|1|Self|Self|Big|General Community||Match Support|1|0|0|1|277|60|598|500000170|500020753|501023677|3|15|1|1|0|1|10|2|-2||2|1||-2||-2|0|10|||7464|9|||1|
502215233|503558339|500709090|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|457|Red||2013-09-04|2013-09-16|2014-12-17|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||15||2|2|1|1|F|Hispanic|Other South American|14|No|Mother|28212|Two Parent|Unknown||||Yes|Big|Neighbor/Friend|General Community|PERL 2014-2016, VOL - Mentoring Hispanic Youth|Match Support|F|White||34|28270||Married|Unknown|28236|1|0|Big For A Day|Special Event|Big|General Community|Amachi|Enrollment|0|1|1|0|277|60|598|500000170|500017777|502215660|3|15|2|1|0|2|10|2|-2||4|3|500011312, 500014681|-2|500000294|-2|6854|8|||16422|8|||1|
502485856|502253272|500537140|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|810|Yellow||2011-05-20|2011-06-02|2013-08-20|Child/Family: Moved|Child/Family: Moved||26.6||2|2|1|1|F|Hispanic|Other South American|13|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Hispanic||63|28227|Bachelors Degree|Married|Education: Teacher||0|0|Recruitment Event|BBBS Board/Staff|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500011746|502486303|3|15|2|3|0|2|5|2|-2||4|2||-2||-2|0|10|||7462|13|||1|
502485856|503544124|500726848|BBBS of Greater Charlotte|Main Office|N|C|Completed|Enrollment|697|Green||2013-11-04|2013-11-15|2015-10-13|Volunteer: Time constraint|Volunteer: Time constraint||22.9||2|2|1|1|F|Hispanic|Other South American|13|No|Mother|28208|One Parent: Female|Unknown||||Yes||Self|General Community||Enrollment|F|Hispanic||39|28278|Associate Degree|Married|Finance||1|8|Self|Self|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500017777|502486303|3|15|2|3|0|2|5|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500553077|500542775|500120499|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1128|Green|Amachi|2006-08-31|2006-09-07|2009-10-09|Child: Family structure changed|Child: Family structure changed||37.1||1|1|1|1|F|Hispanic|Puerto Rican|24||Mother|28269||Unknown||||No||Therapist/Counselor|General Community|Amachi|Match Support|F|White||57|28210||Single|Business: Marketing|28403|2|6|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500003657|500553329|3|11|2|1|0|2|10|2|500003586||4|1|500000294|-2|500000294|-2|0|5|||2238|7|||1|500000294
500905608|500772804|500178425|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1238|Green||2007-05-29|2007-05-31|2010-10-20|Child/Family: Moved|Child/Family: Moved||40.7||1|1|1|1|M|Hispanic|Puerto Rican|22|No|Mother|28025|Two Parent|Unknown||||No||Self|General Community||Match Support|M|White||42|28036|Associate Degree|Divorced|Business: Clerical|28078|9|5|Recruitment Event|Neighbor/Friend|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500905873|3|11|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||7459|10|||1|
500905603|500783324|500185515|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|1188|Green||2007-07-20|2007-07-20|2010-10-20|Child/Family: Moved|Child/Family: Moved||39||2|3|2|2|F|Hispanic|Puerto Rican|20|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||35|28081|Some College|Single|Law: Police Officer||0|0|Bellafonte Presbyter|Faith Organization|Big|General Community|Amachi|Match Support|1|0|1|0|277|60|598|500000170|500002335|500905873|3|11|2|1|0|2|10|2|-2||4|1||-2|500000294|-2|0|10|||2238|7|||1|
500905606|501315871|500283022|BBBS of Greater Charlotte|Main Office|N|C|Completed|Match Support|784|Green||2008-08-21|2008-08-27|2010-10-20|Child/Family: Moved|Child/Family: Moved||25.8||1|1|1|1|F|Hispanic|Puerto Rican|19|No|Mother|28025|One Parent: Female|Unknown||||No||Self|General Community||Match Support|F|White||30|28081|High School Graduate|Married|Finance: Banking||0|0|Self|Self|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500002335|500905873|3|11|2|1|0|2|10|2|-2||4|1||-2||-2|0|10|||7464|9|||1|
500186428|500189441|500037496|BBBS of Greater Charlotte|Main Office|Y|C|Completed|Match Support|3619|Green||2003-11-03|2003-11-03|2013-09-30|Child: Graduated|Child: Graduated||118.9||1|2|2|3|M|Black||21||Mother|28262|One Parent: Female|Unknown||||No||Self|General Community||Match Support|M|White||40|28211|Bachelors Degree|Single|Unknown||0|0|Brochure|Media|Big|General Community||Match Support|1|0|1|0|277|60|598|500000170|500004169|500187986|31|0|1|1|0|1|10|2|-2||4|1||-2||-2|0|10|||127|1|||1|
500186175|500189134|500037134|BBBS of Greater Charlotte|Main Office|Y|C|Completed|Match Support|1820|Green||2004-10-07|2004-10-07|2009-10-01|Child: Graduated|Child: Graduated||59.8||1|2|1|2|M|Black||19||Mother|28273|Other/Unknown|Unknown||||No||Self|General Site||Match Support|F|Multi-Race (None of the above)||46|28277|Bachelors Degree|Single|Business: Sales|28277|7|0|Neighbor/Friend|Neighbor/Friend|Big|General Site||Match Support|1|0|1|0|277|60|598|500000170|500009242|500187759|31|0|1|7|0|2|10|2|-2||4|1||-1||-1|0|10|||7496|10|||1|
500186802|500189243|500037245|BBBS of Greater Charlotte|Main Office|Y|C|Completed|Match Support|1848|Green||2004-09-28|2004-09-28|2009-10-20|Child: Changed school/site|Child: Changed school/site||60.7||1|2|2|3|F|Black||19||Mother|28217|Other/Unknown|Unknown||||No||Self|General Site||Match Support|F|White||51|29732|Some College|Divorced|Business: Clerical|29732|13|0|Recruitment Event|Neighbor/Friend|Big|General Site||Enrollment|1|0|1|0|277|60|598|500000170|500009242|500188104|31|0|2|1|0|2|10|2|-2||4|1||-1||-1|0|10|||7459|10|||1|
503457000|503552518|500710586|BBBS of Greater Charlotte|Main Office|Y|C|Active|Match Support|1265|Green||2013-09-12|2013-09-28|NaT||||41.6||1|3|1|3|F|Black||9|Yes|Mother|28205|One Parent: Female|$20,000 to $24,999|||Y|No||Self|General Community|Amachi|Match Support|F|White||33|28205|Masters Degree|Single|Education: Admin|28027|0|5|Recruitment Event|Other Big|Big|General Community||Match Support|0|1|0|1|277|60|598|500000170|500008321|503458866|31|0|2|1|0|2|10|2|500014421||2|1|500000294|-2||-2|0|10|||7460|12|||1|
