MatchNum|OfficeName|TeamName|Hybrid|MatchType|MatchStatus|MatchName|QueueDescription|TimeInQueue|MatchSupportLevel|MatchReportSources|PendingMatchDate|MatchOpenDate|MatchCloseDate|MatchClosureReasons|MatchClosurePrimaryReason|MatchClosureSecondaryReason|MatchLength|CouplesMatch|MatchCountChild|SegmentMatchCountChild|MatchCountVolunteer|SegmentMatchCountVolunteer|ChildGender|ChildEthnicity|ChildNationality|ChildAge|IncarceratedParent|AdultChildRelationship|ChildZip|ChildGrade|ChildLivingSituation|ChildIncomeLevel|MilitaryParent|ParentDeployed|ChildFamilyAssistance|ChildFreeReducedlunch|CustodialAdultEmployerCity|CustodialAdultEmployerState|CustodialAdultEmployerZipCode|ChildReferralSource|ChildReferralType|ChildAutomaticProgramName|ChildReportSources|ChildActiveQueue|VolGender|VolEthnicity|VolNationality|VolAge|VolZip|VolEducationLevel|VolMaritalStatus|VolOccupation|VolEmployerZipCode|VolEmploymentLengthYears|VolEmploymentLengthMonths|VolReferralSource|VolReferralType|VolunteerType|VolAutomaticProgramName|VolReportSources|VolActiveQueue|Beg|Open|Close|End|AgencyID|AgencyGroupKey|LocationKey|TeamKey|UserKey|ChildPartKey|CustodialAdultKey|ChildEthnicityKey|ChildNationalityKey|ChildGenderKey|VolPartKey|VolEthnicityKey|VolNationalityKey|VolGenderKey|MatchKey|QueueKey|MatchTypeKey|MatchActivityKey|MatchSiteKey|StatusKey|MatchSupportLevelKey|ChildReportSourcesKey|ChildAutomaticProgramKey|VolReportSourcesKey|VolAutomaticProgramKey|ChildReferralSourceKey|ChildReferralSourceTypeKey|ChildPartnerAffiliationKey|ChildPartnerAffiliationTypeKey|VolReferralSourceKey|VolReferralSourceTypeKey|VolPartnerAffiliationKey|VolPartnerAffiliationTypeKey|VolunteerTypeKey|MatchReportSourcesKey|CustodialAdultEmployerHash
CM2|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM2|Enrollment|21|Yellow||2015-12-09|2015-12-18|2016-01-08|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||0.7||1|1|1|1|F|Black||15|No|Mother|28269|8|One Parent: Female|$30,000 to $34,999||||Yes|Charlotte|NC|28269||School|General Community|VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|F|White||26|28078|Masters Degree|Single|Business: Marketing|28269|2|0|Self|Self|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|RTBM|0|1|1|0|277|60|598|500000170|500017777|504458036|504460294|31|0|2|504416792|1|0|2|500866388|5|2|-2||4|2|500011315, 500011316|-2|500007920, 500011315, 500011316|-2|0|4|||7464|9|||1||3086452374500817499
CM6|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM6|Match Support|56|Green||2015-04-23|2015-04-30|2015-06-25|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||1.8||2|2|1|1|F|Black||11|No|Mother|28269|5|One Parent: Female|$50,000 to $59,999|||Y|No|Charlotte|NC|28211||School|General Community||Match Support|F|White||27|28202|Some College|Single|Transport: Flight Attendant||2|1|Local TV|Media|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500017732|504243465|504245581|31|0|2|504173742|1|0|2|500824646|10|2|-2||4|1||-2||-2|0|4|||7438|1|||1||2806833304218536184
CM8|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM8|Match Support|68|Red||2016-12-01|2016-12-22|2017-02-28|Child/Family: Moved|Child/Family: Moved||2.2||1|1|1|1|M|Black||14|No|Mother|28215|9|One Parent: Female|Less than $10,000|||Y|Yes|||||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|M|Black||32|28213|Masters Degree|Married|Finance: Auditor|28202|0|5|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500020753|504851045|504853547|31|0|1|504774982|31|0|1|500932246|10|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316|-2|0|5|||46|2|||1||2141487034287122220
CM9|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM9|Match Support|86|Red|PERL 2014-2016|2015-06-16|2015-06-29|2015-09-23|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||2.8||2|2|1|1|M|American Indian or Alaska Native||12|No|Mother|28269|4|One Parent: Female|$10,000 to $14,999|||Y|Yes|Charlotte|NC|28262||School|General Community|PERL 2014-2016|Match Support|M|White||26|28031||Single|Service: Restaurant|28078|0|2|Self|Self|Big|General Community|Amachi, PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500020752|504150685|504152735|6|0|1|504186384|1|0|1|500830331|10|2|-2||4|3|500014681|-2|500000294, 500014681|-2|0|4|||7464|9|||1|500014681|3402014428779854546
CM10|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM10|Match Support|97|Green|Amachi|2015-09-11|2015-09-23|2015-12-29|Child: Lost interest|Child: Lost interest||3.2||1|1|1|1|F|Black||10|Yes|GrandMother|28217|4|Grandparents|Less than $10,000|||Y|Yes|||||School|General Community|Amachi|Match Support|F|White||32|28277|Masters Degree|Divorced|Tech: Computer/Programmer|28277|0|3|Self|Self|Big|General Community|Amachi|Match Support|0|1|1|0|277|60|598|500000170|500017732|504195472|504197572|31|0|2|504222207|1|0|2|500839514|10|2|-2||4|1|500000294|-2|500000294|-2|0|4|||7464|9|||1|500000294|0
CM13|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM13|Enrollment|111|Red|PERL 2014-2016|2015-08-06|2015-08-11|2015-11-30|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.6||1|1|1|1|F|Multi-race (Black & White)||13|No|Mother|28212|6|One Parent: Female|$10,000 to $14,999|||Y|Yes|Charlotte|NC|28212||Relative|General Community|PERL 2014-2016|Enrollment|F|White||47|28270|Some College|Married|Homemaker|29020|18|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500008321|504280484|504282684|36|0|2|504226821|1|0|2|500835375|5|2|-2||4|3|500014681|-2||-2|0|3|||7464|9|||1|500014681|4694273237201497095
CM14|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM14|Match Support|111|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-01-14|2016-01-30|2016-05-20|Volunteer: Moved|Volunteer: Moved||3.6||2|2|1|1|F|Black||12|No|Mother|28214|5|One Parent: Female|$15,000 to $19,999|||Y|Yes|Charlotte|NC|28262|BBBS National Site|Web Link|General Community||Match Support|F|White||32|28208|Bachelors Degree|Single|Journalist/Media||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017777|503976557|503978568|31|0|2|504365048|1|0|2|500871811|10|2|-2||4|1||-2||-2|34|2|||7464|9|||1|500007920, 500011315, 500011316|3198188609986797983
CM16|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM16|Enrollment|120|Green|PERL 2014-2016|2016-10-24|2016-10-31|2017-02-28|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||3.9||4|4|1|1|F|Black||13|Yes|Mother|28217|8|One Parent: Female|Unknown||||Yes|||||Self|General Community|PERL 2014-2016|Enrollment|F|White||31|28278|Doctor of Medicine (MD)|Living w/ Significant Other|Medical: Pharmacist||0|0|BBBS National Site|Web Link|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500013781|501319029|500948399|31|0|2|504558901|1|0|2|500918750|5|2|-2||4|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||46|2|||1|500014681|0
CM22|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM22|Enrollment|135|Green|PERL 2014-2016|2015-10-01|2015-10-21|2016-03-04|Child/Family: Moved|Child/Family: Moved||4.4||1|1|2|2|M|Black||14|No|Mother|28212|5|One Parent: Female|$10,000 to $14,999|||Y|Yes|||||Therapist/Counselor|General Community|Amachi, PERL 2014-2016|Enrollment|M|White||30|28209|Bachelors Degree|Married|Real Estate: Realtor|28217|0|9|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|503863366|503865360|31|0|1|504322037|1|0|1|500843765|5|2|-2||4|1|500000294, 500014681|-2||-2|0|5|||46|2|||1|500014681|0
CM25|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM25|RTBM|136|Green||2016-05-11|2016-06-20|2016-11-03|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||4.5||1|1|1|1|F|Black||14|No|GrandMother|28105|9|Grandparents|$45,000 to $49,999||||Yes||||BBBS National Site|Web Link|General Community||RTBM|F|Black||39|28105|Bachelors Degree|Single|Unemployed||0|0|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504631841|504634252|31|0|2|504167347|31|0|2|500892753|7|2|-2||4|1||-2||-2|34|2|||7464|9|||1||5605796235524810842
CM30|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM30|Enrollment|157|Green|PERL 2014-2016|2015-11-17|2015-12-14|2016-05-19|Volunteer: Moved|Volunteer: Moved||5.2||1|1|1|1|F|Black||16|No|Mother|28215|8|One Parent: Female|Less than $10,000|||Y|Yes|||||Self|General Community|PERL 2014-2016|Enrollment|F|White||25|28205|Bachelors Degree|Single|Business|28031|0|0|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500017777|503611723|503613600|31|0|2|504295160|1|0|2|500860670|5|2|-2||4|1|500014681|-2|500014681|-2|0|10|||17159|12|||1|500014681|0
CM31|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM31|Match Support|161|Yellow||2015-07-30|2015-07-30|2016-01-07|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||5.3||1|1|1|1|M|Black||14|No|Mother|28217|6|One Parent: Female|$10,000 to $14,999|||Y|Yes|Charlotte|NC|28217|BBBS National Site|Web Link|General Community||Match Support|M|White||31|28209|Bachelors Degree|Single|Human Services|28203|1|8|Current/Previous Big|Other Big|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500018851|503063769|503065429|31|0|1|504299841|1|0|1|500834948|10|2|-2||4|2||-2||-2|34|2|||17159|12|||1||2141487034287122220
CM33|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM33|Match Support|167|Yellow||2015-07-28|2015-07-28|2016-01-11|Child/Family: Feels incompatible with volunteer|Child/Family: Feels incompatible with volunteer||5.5||1|1|1|1|F|Black||13|No|Mother|28217|6|One Parent: Female|$10,000 to $14,999|||Y|Yes|Charlotte|NC|28217||School|General Community||Match Support|F|White||26|28203|Bachelors Degree|Single|Finance: Banking||2|2|Self|Self|Big|General Community||Enrollment|0|1|1|0|277|60|598|500000170|500018851|504230613|503065429|31|0|2|503995309|1|0|2|500834694|10|2|-2||4|2||-2||-2|0|4|||7464|9|||1||2141487034287122220
CM34|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM34|Match Support|169|Red||2015-11-10|2015-12-07|2016-05-24|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||5.6||1|1|1|1|M|Black||14|No|Mother|28027|7|One Parent: Female|$25,000 to $29,999||||Yes|Charlotte|NC|28217||School|General Community||Match Support|M|White||24|28262||Single|Medical: Healthcare Worker|28025|1|0|Current/Previous Big|Other Big|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020753|502129820|502130249|31|0|1|504474407|1|0|1|500858150|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|4|||17159|12|||1||2881622112345502539
CM39|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM39|Pending Match|176|Red|PERL 2014-2016|2015-03-26|2015-04-14|2015-10-07|Volunteer: Moved|Volunteer: Moved||5.8||1|2|1|1|F|Multi-race (Hispanic & White)||13|No|Mother|28205|7|One Parent: Female|$10,000 to $14,999|||Y|Yes|Charlotte|NC|28202||Therapist/Counselor|General Community||Pending Match|F|White||30|28205|Bachelors Degree|Separated|Business|28205|0|7|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500013781|504205508|504207619|35|0|2|504157187|1|0|2|500820606|9|2|-2||4|3||-2|500014681|-2|0|5|||17159|12|||1|500014681|610388910998118020
CM42|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM42|Match Support|194|Green||2015-05-28|2015-06-18|2015-12-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||6.4||1|1|1|1|M|Black||13|Yes|Mother|28214|5|One Parent: Female|$20,000 to $24,999|||Y|Yes|Charlotte|NC|28269|BBBS National Site|Web Link|General Community|Amachi|Match Support|M|Asian|Indian|49|28203|Bachelors Degree|Married|Tech: Engineer|28204|10|0|Current/Previous Big|Other Big|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504217755|504219869|31|0|1|504131744|4|18|1|500828564|10|2|-2||4|1|500000294|-2||-2|34|2|||17159|12|||1||7000602719972091240
CM51|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM51|Match Support|221|Green|PERL 2014-2016|2016-01-11|2016-01-21|2016-08-29|Volunteer: Feels incompatible with child/family|Volunteer: Feels incompatible with child/family||7.3||1|1|1|1|M|Black||15|No|Mother|28269|7|One Parent: Female|$10,000 to $14,999|||Y|Yes|Charlotte|NC|28217||School|General Community|PERL 2014-2016|Match Support|M|Multi-race (Black & White)||27|28115|Bachelors Degree|Single|Business|28115|4|4|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500017777|504268284|504270481|31|0|1|503172653|36|0|1|500871097|10|2|-2||4|1|500014681|-2|500007920, 500011315, 500011316, 500014681|-2|0|4|||7464|9|||1|500014681|2378213070582218846
CM56|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM56|RTBM|228|Green|PERL 2014-2016|2015-11-09|2016-01-14|2016-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.5||1|1|1|1|F|Black||10|No|Mother|28056|4|One Parent: Female|$15,000 to $19,999|||Y|Yes|||||Self|General Community||RTBM|F|White||30|28209|Bachelors Degree|Single|Finance: Banking|28211|3|2|Self|Self|Big|General Community|PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500017777|504407275|504409521|31|0|2|504393547|1|0|2|500857377|7|2|-2||4|1||-2|500007920, 500011315, 500011316, 500014681|-2|0|10|||7464|9|||1|500014681|0
CM60|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM60|Match Support|238|Red||2016-05-04|2016-05-27|2017-01-20|Child: Severity of challenges|Child: Severity of challenges||7.8||1|1|1|1|M|Black||14|No|Mother|28215|7|One Parent: Female|$15,000 to $19,999|||Y|Yes|||||School|General Community||Match Support|M|White||23|28205|Bachelors Degree|Single|Finance|28210|0|11|BBBS National Site|Web Link|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Enrollment|0|1|1|0|277|60|598|500000170|500008321|504318423|504320644|31|0|1|504561410|1|0|1|500891770|10|2|-2||4|3||-2|500007920, 500011315, 500011316|-2|0|4|||46|2|||1||2141487034287122220
CM62|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM62|Match Support|241|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment|2016-05-02|2016-05-31|2017-01-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||7.9||1|1|2|2|M|White||14|No|Mother|28214|7|One Parent: Female|$10,000 to $14,999|||Y|Yes|||||Relative|General Community||Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500013781|504231264|504233379|1|0|1|504230177|1|0|1|500891315|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|0|3|||7462|13|||1|500007920, 500011315, 500011316|0
CM64|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM64|Match Support|241|Red|PERL 2014-2016|2015-06-28|2015-06-28|2016-02-24|Child/Family: Time constraints|Child/Family: Time constraints||7.9||1|1|2|2|M|Black||11|No|Mother|28226|3|One Parent: Female|$30,000 to $34,999|||Y|Yes|||||School|General Community|PERL 2014-2016|Match Support|M|White||26|28012|Some College|Single|Finance|28255|4|4|Recruitment Event|BBBS Board/Staff|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500013781|504198439|504200550|31|0|1|504230177|1|0|1|500831539|10|2|-2||4|3|500014681|-2|500007920, 500011315, 500011316|-2|0|4|||7462|13|||1|500014681|0
CM70|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM70|Match Support|254|Green|PERL 2014-2016|2015-06-23|2015-06-23|2016-03-03|Child/Family: Moved|Child/Family: Moved||8.3||1|1|1|1|F|Black||13|No|Mother|28134|6|One Parent: Female|Less than $10,000|||Y|Yes|||||Therapist/Counselor|General Community|PERL 2014-2016|Match Support|F|White||30|28277|Bachelors Degree|Single|Business: Clerical|28277|1|7|Self|Self|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500018851|502205926|502206355|31|0|2|504225335|1|0|2|500831147|10|2|-2||4|1|500014681|-2||-2|0|5|||7464|9|||1|500014681|6178126991714892144
CM71|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM71|RTBM|256|Green|VOL - PreMatch, VOL - PreMatchILT, VOL - PreMatch Training Final Assessment, PERL 2014-2016|2015-12-07|2015-12-17|2016-08-29|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||8.4||1|1|1|1|M|Black||14|No|Mother|28269|7|One Parent: Female|Less than $10,000|||Y|Yes|||||School|General Community||RTBM|M|Black||40|28269|Bachelors Degree|Married|Tech: Support, Writing|28269|4|0|Local Radio|Media|Big|General Community|Amachi, PERL 2014-2016, VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500017777|504245120|504247236|31|0|1|504396885|31|0|1|500865817|7|2|-2||4|1||-2|500000294, 500007920, 500011315, 500011316, 500014681|-2|0|4|||7437|1|||1|500007920, 500011315, 500011316, 500014681|1546374315672654438
CM74|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM74|Match Support|275|Green||2016-05-10|2016-05-24|2017-02-23|Volunteer: Moved|Volunteer: Moved||9||1|1|1|1|M|Black||15|No|Mother|28208|9|One Parent: Female|$20,000 to $24,999|||Y|Yes||||BBBS National Site|Web Link|General Community||Match Support|M|White||32|28203|PHD|Single|Self-Employed, Entrepreneur|30604|4|0|Local Print|Media|Big|General Community|VOL - PreMatch, VOL - PreMatch Training Final Assessment, VOL - PreMatchILT|Match Support|0|1|1|0|277|60|598|500000170|500020910|504347348|504349572|31|0|1|504566830|1|0|1|500892524|10|2|-2||4|1||-2|500007920, 500011315, 500011316|-2|34|2|||7439|1|||1||7044657180546140448
CM78|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM78|Match Support|288|Yellow|PERL 2014-2016|2015-05-14|2015-05-31|2016-03-14|Child/Family: Moved|Child/Family: Moved||9.5||1|1|1|1|M|Multi-race (Black & White)||13|No|Mother|28134|4|One Parent: Female|$10,000 to $14,999|||Y|Yes|Pineville|NC|28134||School|General Community|PERL 2014-2016|Match Support|M|White||26|28273|Bachelors Degree|Single|Architect|28273|0|11|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500008321|504202968|504205079|36|0|1|504285700|1|0|1|500827095|10|2|-2||4|2|500014681|-2|500014681|-2|0|4|||17159|12|||1|500014681|7165641474360673060
CM87|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM87|Match Support|330|Red|PERL 2014-2016|2015-05-05|2015-06-02|2016-04-27|Volunteer: Lost contact with child/agency|Volunteer: Lost contact with child/agency||10.8||1|1|1|1|M|Black||15|No|Mother|28273|8|One Parent: Female|$35,000 to $39,999||||No|Charlotte|NC|28273|BBBS National Site|Web Link|General Community|PERL 2014-2016|Match Support|M|White||30|28208|Bachelors Degree|Single|Self-Employed, Entrepreneur|28078|2|3|Current/Previous Big|Other Big|Big|General Community|PERL 2014-2016|Match Support|0|1|1|0|277|60|598|500000170|500013781|504159888|504161941|31|0|1|504240720|1|0|1|500825834|10|2|-2||4|3|500014681|-2|500014681|-2|34|2|||17159|12|||1|500014681|8491998754880714879
CM92|BBBS of Greater Charlotte|Main Office|N|C|Completed|CM92|RTBM|332|Green||2015-10-09|2015-10-26|2016-09-22|Volunteer: Moved|Volunteer: Moved||10.9||1|1|1|1|M|Black||9|No|Mother|28211|4|One Parent: Female|$25,000 to $29,999|Yes: Active|No|Y|Yes|Charlotte|NC|28216||Self|General Community||RTBM|M|Multi-race (Black & White)||26|28211|Some College|Single|Finance|28210|0|5|BBBS National Site|Web Link|Big|General Community||Match Support|0|1|1|0|277|60|598|500000170|500017732|504345299|504347523|31|0|1|504397824|36|0|1|500846354|7|2|-2||4|1||-2||-2|0|10|||46|2|||1||1981915209225039472
